// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 28 2022 12:21:15

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__37833;
    wire N__37832;
    wire N__37831;
    wire N__37822;
    wire N__37821;
    wire N__37820;
    wire N__37813;
    wire N__37812;
    wire N__37811;
    wire N__37804;
    wire N__37803;
    wire N__37802;
    wire N__37795;
    wire N__37794;
    wire N__37793;
    wire N__37786;
    wire N__37785;
    wire N__37784;
    wire N__37777;
    wire N__37776;
    wire N__37775;
    wire N__37768;
    wire N__37767;
    wire N__37766;
    wire N__37759;
    wire N__37758;
    wire N__37757;
    wire N__37750;
    wire N__37749;
    wire N__37748;
    wire N__37741;
    wire N__37740;
    wire N__37739;
    wire N__37732;
    wire N__37731;
    wire N__37730;
    wire N__37723;
    wire N__37722;
    wire N__37721;
    wire N__37714;
    wire N__37713;
    wire N__37712;
    wire N__37705;
    wire N__37704;
    wire N__37703;
    wire N__37696;
    wire N__37695;
    wire N__37694;
    wire N__37687;
    wire N__37686;
    wire N__37685;
    wire N__37678;
    wire N__37677;
    wire N__37676;
    wire N__37669;
    wire N__37668;
    wire N__37667;
    wire N__37660;
    wire N__37659;
    wire N__37658;
    wire N__37651;
    wire N__37650;
    wire N__37649;
    wire N__37642;
    wire N__37641;
    wire N__37640;
    wire N__37633;
    wire N__37632;
    wire N__37631;
    wire N__37624;
    wire N__37623;
    wire N__37622;
    wire N__37615;
    wire N__37614;
    wire N__37613;
    wire N__37606;
    wire N__37605;
    wire N__37604;
    wire N__37597;
    wire N__37596;
    wire N__37595;
    wire N__37588;
    wire N__37587;
    wire N__37586;
    wire N__37579;
    wire N__37578;
    wire N__37577;
    wire N__37570;
    wire N__37569;
    wire N__37568;
    wire N__37561;
    wire N__37560;
    wire N__37559;
    wire N__37552;
    wire N__37551;
    wire N__37550;
    wire N__37543;
    wire N__37542;
    wire N__37541;
    wire N__37534;
    wire N__37533;
    wire N__37532;
    wire N__37525;
    wire N__37524;
    wire N__37523;
    wire N__37516;
    wire N__37515;
    wire N__37514;
    wire N__37507;
    wire N__37506;
    wire N__37505;
    wire N__37498;
    wire N__37497;
    wire N__37496;
    wire N__37489;
    wire N__37488;
    wire N__37487;
    wire N__37480;
    wire N__37479;
    wire N__37478;
    wire N__37471;
    wire N__37470;
    wire N__37469;
    wire N__37462;
    wire N__37461;
    wire N__37460;
    wire N__37453;
    wire N__37452;
    wire N__37451;
    wire N__37444;
    wire N__37443;
    wire N__37442;
    wire N__37435;
    wire N__37434;
    wire N__37433;
    wire N__37426;
    wire N__37425;
    wire N__37424;
    wire N__37417;
    wire N__37416;
    wire N__37415;
    wire N__37408;
    wire N__37407;
    wire N__37406;
    wire N__37399;
    wire N__37398;
    wire N__37397;
    wire N__37390;
    wire N__37389;
    wire N__37388;
    wire N__37381;
    wire N__37380;
    wire N__37379;
    wire N__37372;
    wire N__37371;
    wire N__37370;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37343;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37327;
    wire N__37324;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37298;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37253;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37119;
    wire N__37116;
    wire N__37115;
    wire N__37114;
    wire N__37113;
    wire N__37112;
    wire N__37111;
    wire N__37110;
    wire N__37109;
    wire N__37108;
    wire N__37107;
    wire N__37106;
    wire N__37105;
    wire N__37100;
    wire N__37097;
    wire N__37092;
    wire N__37083;
    wire N__37082;
    wire N__37081;
    wire N__37080;
    wire N__37079;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37034;
    wire N__37031;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36981;
    wire N__36978;
    wire N__36977;
    wire N__36976;
    wire N__36975;
    wire N__36974;
    wire N__36973;
    wire N__36972;
    wire N__36971;
    wire N__36970;
    wire N__36969;
    wire N__36968;
    wire N__36967;
    wire N__36966;
    wire N__36965;
    wire N__36964;
    wire N__36963;
    wire N__36962;
    wire N__36961;
    wire N__36960;
    wire N__36959;
    wire N__36958;
    wire N__36957;
    wire N__36956;
    wire N__36955;
    wire N__36954;
    wire N__36953;
    wire N__36952;
    wire N__36951;
    wire N__36950;
    wire N__36949;
    wire N__36948;
    wire N__36947;
    wire N__36946;
    wire N__36945;
    wire N__36944;
    wire N__36943;
    wire N__36942;
    wire N__36941;
    wire N__36940;
    wire N__36939;
    wire N__36938;
    wire N__36937;
    wire N__36936;
    wire N__36935;
    wire N__36934;
    wire N__36933;
    wire N__36932;
    wire N__36931;
    wire N__36930;
    wire N__36929;
    wire N__36928;
    wire N__36927;
    wire N__36926;
    wire N__36925;
    wire N__36924;
    wire N__36923;
    wire N__36922;
    wire N__36921;
    wire N__36920;
    wire N__36919;
    wire N__36918;
    wire N__36917;
    wire N__36916;
    wire N__36915;
    wire N__36914;
    wire N__36913;
    wire N__36912;
    wire N__36911;
    wire N__36910;
    wire N__36909;
    wire N__36908;
    wire N__36907;
    wire N__36906;
    wire N__36905;
    wire N__36904;
    wire N__36903;
    wire N__36902;
    wire N__36901;
    wire N__36900;
    wire N__36899;
    wire N__36898;
    wire N__36897;
    wire N__36896;
    wire N__36895;
    wire N__36894;
    wire N__36893;
    wire N__36892;
    wire N__36891;
    wire N__36890;
    wire N__36889;
    wire N__36888;
    wire N__36887;
    wire N__36886;
    wire N__36885;
    wire N__36884;
    wire N__36883;
    wire N__36882;
    wire N__36881;
    wire N__36880;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36876;
    wire N__36875;
    wire N__36874;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36870;
    wire N__36869;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36864;
    wire N__36863;
    wire N__36862;
    wire N__36861;
    wire N__36860;
    wire N__36859;
    wire N__36858;
    wire N__36857;
    wire N__36856;
    wire N__36855;
    wire N__36854;
    wire N__36853;
    wire N__36852;
    wire N__36851;
    wire N__36850;
    wire N__36849;
    wire N__36848;
    wire N__36847;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36575;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36565;
    wire N__36562;
    wire N__36561;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36540;
    wire N__36535;
    wire N__36532;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36411;
    wire N__36408;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36387;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36356;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36348;
    wire N__36345;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36334;
    wire N__36333;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36325;
    wire N__36324;
    wire N__36323;
    wire N__36318;
    wire N__36315;
    wire N__36314;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36303;
    wire N__36302;
    wire N__36301;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36272;
    wire N__36267;
    wire N__36260;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36252;
    wire N__36249;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36222;
    wire N__36219;
    wire N__36214;
    wire N__36211;
    wire N__36204;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36182;
    wire N__36177;
    wire N__36174;
    wire N__36169;
    wire N__36166;
    wire N__36159;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36147;
    wire N__36144;
    wire N__36143;
    wire N__36142;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36129;
    wire N__36128;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36105;
    wire N__36104;
    wire N__36103;
    wire N__36102;
    wire N__36101;
    wire N__36100;
    wire N__36099;
    wire N__36098;
    wire N__36097;
    wire N__36096;
    wire N__36095;
    wire N__36094;
    wire N__36093;
    wire N__36092;
    wire N__36091;
    wire N__36090;
    wire N__36089;
    wire N__36088;
    wire N__36087;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36035;
    wire N__36030;
    wire N__36029;
    wire N__36028;
    wire N__36027;
    wire N__36026;
    wire N__36025;
    wire N__36024;
    wire N__36023;
    wire N__36022;
    wire N__36021;
    wire N__36020;
    wire N__36019;
    wire N__36018;
    wire N__36017;
    wire N__36016;
    wire N__36015;
    wire N__36014;
    wire N__36013;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36009;
    wire N__36008;
    wire N__36007;
    wire N__36006;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35864;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35849;
    wire N__35848;
    wire N__35847;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35839;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35831;
    wire N__35830;
    wire N__35827;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35802;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35762;
    wire N__35759;
    wire N__35754;
    wire N__35751;
    wire N__35746;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35730;
    wire N__35727;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35709;
    wire N__35708;
    wire N__35707;
    wire N__35706;
    wire N__35705;
    wire N__35704;
    wire N__35703;
    wire N__35702;
    wire N__35701;
    wire N__35700;
    wire N__35699;
    wire N__35698;
    wire N__35697;
    wire N__35696;
    wire N__35695;
    wire N__35694;
    wire N__35693;
    wire N__35692;
    wire N__35691;
    wire N__35690;
    wire N__35689;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35674;
    wire N__35667;
    wire N__35658;
    wire N__35645;
    wire N__35644;
    wire N__35643;
    wire N__35642;
    wire N__35641;
    wire N__35638;
    wire N__35631;
    wire N__35630;
    wire N__35629;
    wire N__35628;
    wire N__35627;
    wire N__35626;
    wire N__35625;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35609;
    wire N__35606;
    wire N__35601;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35584;
    wire N__35577;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35559;
    wire N__35554;
    wire N__35545;
    wire N__35542;
    wire N__35541;
    wire N__35540;
    wire N__35535;
    wire N__35532;
    wire N__35525;
    wire N__35520;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35481;
    wire N__35478;
    wire N__35475;
    wire N__35472;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35385;
    wire N__35382;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35361;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35343;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35310;
    wire N__35307;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35285;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35270;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35234;
    wire N__35233;
    wire N__35230;
    wire N__35229;
    wire N__35228;
    wire N__35225;
    wire N__35224;
    wire N__35221;
    wire N__35220;
    wire N__35219;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35204;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35189;
    wire N__35184;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35172;
    wire N__35169;
    wire N__35168;
    wire N__35165;
    wire N__35164;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35137;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35114;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35080;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35055;
    wire N__35050;
    wire N__35047;
    wire N__35040;
    wire N__35039;
    wire N__35038;
    wire N__35037;
    wire N__35036;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35007;
    wire N__34998;
    wire N__34997;
    wire N__34996;
    wire N__34995;
    wire N__34994;
    wire N__34993;
    wire N__34992;
    wire N__34991;
    wire N__34988;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34956;
    wire N__34955;
    wire N__34954;
    wire N__34953;
    wire N__34948;
    wire N__34943;
    wire N__34938;
    wire N__34931;
    wire N__34928;
    wire N__34921;
    wire N__34914;
    wire N__34913;
    wire N__34912;
    wire N__34911;
    wire N__34910;
    wire N__34907;
    wire N__34906;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34890;
    wire N__34889;
    wire N__34886;
    wire N__34881;
    wire N__34878;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34840;
    wire N__34833;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34829;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34821;
    wire N__34820;
    wire N__34819;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34772;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34754;
    wire N__34749;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34717;
    wire N__34710;
    wire N__34709;
    wire N__34708;
    wire N__34703;
    wire N__34700;
    wire N__34699;
    wire N__34694;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34683;
    wire N__34682;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34676;
    wire N__34675;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34640;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34608;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34577;
    wire N__34574;
    wire N__34573;
    wire N__34570;
    wire N__34569;
    wire N__34566;
    wire N__34561;
    wire N__34558;
    wire N__34553;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34529;
    wire N__34526;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34490;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34445;
    wire N__34444;
    wire N__34443;
    wire N__34442;
    wire N__34441;
    wire N__34440;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34428;
    wire N__34425;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34417;
    wire N__34414;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34359;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34307;
    wire N__34304;
    wire N__34303;
    wire N__34302;
    wire N__34301;
    wire N__34298;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34244;
    wire N__34241;
    wire N__34236;
    wire N__34231;
    wire N__34228;
    wire N__34215;
    wire N__34214;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34190;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34176;
    wire N__34175;
    wire N__34174;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34157;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34137;
    wire N__34136;
    wire N__34135;
    wire N__34132;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34112;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34086;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34062;
    wire N__34059;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34037;
    wire N__34034;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34019;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33982;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33935;
    wire N__33934;
    wire N__33933;
    wire N__33932;
    wire N__33931;
    wire N__33928;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33907;
    wire N__33906;
    wire N__33903;
    wire N__33898;
    wire N__33897;
    wire N__33894;
    wire N__33889;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33864;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33850;
    wire N__33847;
    wire N__33846;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33836;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33792;
    wire N__33791;
    wire N__33790;
    wire N__33787;
    wire N__33786;
    wire N__33785;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33777;
    wire N__33776;
    wire N__33775;
    wire N__33774;
    wire N__33773;
    wire N__33772;
    wire N__33771;
    wire N__33768;
    wire N__33761;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33749;
    wire N__33748;
    wire N__33743;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33725;
    wire N__33720;
    wire N__33717;
    wire N__33714;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33697;
    wire N__33694;
    wire N__33687;
    wire N__33684;
    wire N__33675;
    wire N__33666;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33639;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33613;
    wire N__33612;
    wire N__33605;
    wire N__33602;
    wire N__33601;
    wire N__33600;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33582;
    wire N__33581;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33524;
    wire N__33521;
    wire N__33516;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33493;
    wire N__33490;
    wire N__33483;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33459;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33432;
    wire N__33429;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33411;
    wire N__33408;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33400;
    wire N__33395;
    wire N__33392;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33372;
    wire N__33371;
    wire N__33364;
    wire N__33361;
    wire N__33360;
    wire N__33359;
    wire N__33356;
    wire N__33355;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33334;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33312;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33257;
    wire N__33252;
    wire N__33251;
    wire N__33250;
    wire N__33247;
    wire N__33246;
    wire N__33245;
    wire N__33244;
    wire N__33241;
    wire N__33240;
    wire N__33239;
    wire N__33236;
    wire N__33233;
    wire N__33228;
    wire N__33227;
    wire N__33224;
    wire N__33219;
    wire N__33216;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33183;
    wire N__33174;
    wire N__33171;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33065;
    wire N__33064;
    wire N__33061;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33040;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33032;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33005;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32984;
    wire N__32983;
    wire N__32982;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32964;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32938;
    wire N__32937;
    wire N__32930;
    wire N__32927;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32909;
    wire N__32908;
    wire N__32903;
    wire N__32900;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32882;
    wire N__32879;
    wire N__32878;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32847;
    wire N__32844;
    wire N__32843;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32831;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32799;
    wire N__32798;
    wire N__32795;
    wire N__32794;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32747;
    wire N__32744;
    wire N__32743;
    wire N__32740;
    wire N__32739;
    wire N__32738;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32728;
    wire N__32725;
    wire N__32722;
    wire N__32721;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32706;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32681;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32660;
    wire N__32657;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32621;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32557;
    wire N__32554;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32444;
    wire N__32443;
    wire N__32442;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32430;
    wire N__32427;
    wire N__32426;
    wire N__32421;
    wire N__32418;
    wire N__32417;
    wire N__32414;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32406;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32303;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32268;
    wire N__32267;
    wire N__32266;
    wire N__32263;
    wire N__32258;
    wire N__32255;
    wire N__32250;
    wire N__32249;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32217;
    wire N__32216;
    wire N__32215;
    wire N__32214;
    wire N__32213;
    wire N__32212;
    wire N__32211;
    wire N__32210;
    wire N__32209;
    wire N__32208;
    wire N__32207;
    wire N__32206;
    wire N__32205;
    wire N__32204;
    wire N__32203;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32138;
    wire N__32137;
    wire N__32134;
    wire N__32129;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32103;
    wire N__32100;
    wire N__32099;
    wire N__32098;
    wire N__32097;
    wire N__32094;
    wire N__32089;
    wire N__32086;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32070;
    wire N__32067;
    wire N__32066;
    wire N__32065;
    wire N__32064;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32052;
    wire N__32049;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31831;
    wire N__31830;
    wire N__31825;
    wire N__31820;
    wire N__31815;
    wire N__31812;
    wire N__31811;
    wire N__31810;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31797;
    wire N__31796;
    wire N__31791;
    wire N__31788;
    wire N__31783;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31763;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31739;
    wire N__31738;
    wire N__31737;
    wire N__31734;
    wire N__31727;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31706;
    wire N__31703;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31685;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31661;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31639;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31625;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31598;
    wire N__31595;
    wire N__31590;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31578;
    wire N__31575;
    wire N__31566;
    wire N__31563;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31555;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31539;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31493;
    wire N__31492;
    wire N__31491;
    wire N__31490;
    wire N__31489;
    wire N__31488;
    wire N__31487;
    wire N__31486;
    wire N__31485;
    wire N__31484;
    wire N__31483;
    wire N__31482;
    wire N__31481;
    wire N__31480;
    wire N__31479;
    wire N__31476;
    wire N__31465;
    wire N__31458;
    wire N__31451;
    wire N__31442;
    wire N__31431;
    wire N__31428;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31406;
    wire N__31401;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31393;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31369;
    wire N__31362;
    wire N__31361;
    wire N__31360;
    wire N__31357;
    wire N__31356;
    wire N__31355;
    wire N__31352;
    wire N__31351;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31307;
    wire N__31304;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31292;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31264;
    wire N__31263;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31236;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31215;
    wire N__31214;
    wire N__31213;
    wire N__31210;
    wire N__31209;
    wire N__31206;
    wire N__31205;
    wire N__31202;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31184;
    wire N__31179;
    wire N__31178;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31159;
    wire N__31156;
    wire N__31149;
    wire N__31148;
    wire N__31147;
    wire N__31146;
    wire N__31145;
    wire N__31144;
    wire N__31143;
    wire N__31142;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31127;
    wire N__31126;
    wire N__31125;
    wire N__31124;
    wire N__31123;
    wire N__31122;
    wire N__31121;
    wire N__31120;
    wire N__31119;
    wire N__31118;
    wire N__31117;
    wire N__31116;
    wire N__31115;
    wire N__31112;
    wire N__31111;
    wire N__31108;
    wire N__31107;
    wire N__31106;
    wire N__31105;
    wire N__31104;
    wire N__31103;
    wire N__31102;
    wire N__31101;
    wire N__31098;
    wire N__31097;
    wire N__31090;
    wire N__31085;
    wire N__31084;
    wire N__31083;
    wire N__31082;
    wire N__31077;
    wire N__31076;
    wire N__31073;
    wire N__31068;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31049;
    wire N__31046;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31004;
    wire N__31003;
    wire N__31002;
    wire N__31001;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30987;
    wire N__30982;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30949;
    wire N__30948;
    wire N__30947;
    wire N__30946;
    wire N__30945;
    wire N__30944;
    wire N__30943;
    wire N__30940;
    wire N__30935;
    wire N__30932;
    wire N__30923;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30905;
    wire N__30898;
    wire N__30891;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30854;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30815;
    wire N__30812;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30797;
    wire N__30794;
    wire N__30787;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30771;
    wire N__30770;
    wire N__30765;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30728;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30692;
    wire N__30691;
    wire N__30690;
    wire N__30687;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30669;
    wire N__30668;
    wire N__30667;
    wire N__30666;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30620;
    wire N__30615;
    wire N__30606;
    wire N__30605;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30597;
    wire N__30594;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30572;
    wire N__30569;
    wire N__30558;
    wire N__30557;
    wire N__30556;
    wire N__30553;
    wire N__30552;
    wire N__30549;
    wire N__30548;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30519;
    wire N__30516;
    wire N__30507;
    wire N__30506;
    wire N__30505;
    wire N__30500;
    wire N__30497;
    wire N__30492;
    wire N__30489;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30481;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30443;
    wire N__30442;
    wire N__30439;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30417;
    wire N__30416;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30393;
    wire N__30390;
    wire N__30387;
    wire N__30378;
    wire N__30377;
    wire N__30376;
    wire N__30375;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30347;
    wire N__30344;
    wire N__30339;
    wire N__30332;
    wire N__30327;
    wire N__30324;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30284;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30256;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30230;
    wire N__30229;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30215;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30110;
    wire N__30107;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30067;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30030;
    wire N__30029;
    wire N__30026;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29969;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29945;
    wire N__29942;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29918;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29898;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29820;
    wire N__29819;
    wire N__29816;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29799;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29763;
    wire N__29762;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29751;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29736;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29711;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29700;
    wire N__29699;
    wire N__29698;
    wire N__29697;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29685;
    wire N__29684;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29662;
    wire N__29657;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29633;
    wire N__29630;
    wire N__29619;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29586;
    wire N__29585;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29552;
    wire N__29549;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29519;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29496;
    wire N__29493;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29481;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29417;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29406;
    wire N__29403;
    wire N__29402;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29376;
    wire N__29375;
    wire N__29374;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29349;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29319;
    wire N__29318;
    wire N__29317;
    wire N__29316;
    wire N__29315;
    wire N__29312;
    wire N__29307;
    wire N__29300;
    wire N__29299;
    wire N__29298;
    wire N__29297;
    wire N__29292;
    wire N__29289;
    wire N__29284;
    wire N__29277;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29240;
    wire N__29239;
    wire N__29236;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29214;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29107;
    wire N__29106;
    wire N__29103;
    wire N__29102;
    wire N__29099;
    wire N__29098;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29083;
    wire N__29082;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29069;
    wire N__29068;
    wire N__29067;
    wire N__29066;
    wire N__29065;
    wire N__29064;
    wire N__29063;
    wire N__29062;
    wire N__29061;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29046;
    wire N__29043;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29029;
    wire N__29026;
    wire N__29025;
    wire N__29024;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29016;
    wire N__29015;
    wire N__29012;
    wire N__29011;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__29002;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28990;
    wire N__28989;
    wire N__28986;
    wire N__28985;
    wire N__28982;
    wire N__28981;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28961;
    wire N__28958;
    wire N__28955;
    wire N__28952;
    wire N__28949;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28939;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28892;
    wire N__28887;
    wire N__28878;
    wire N__28875;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28854;
    wire N__28853;
    wire N__28852;
    wire N__28851;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28843;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28826;
    wire N__28813;
    wire N__28810;
    wire N__28809;
    wire N__28808;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28779;
    wire N__28778;
    wire N__28777;
    wire N__28772;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28757;
    wire N__28754;
    wire N__28753;
    wire N__28750;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28738;
    wire N__28737;
    wire N__28736;
    wire N__28733;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28704;
    wire N__28691;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28660;
    wire N__28653;
    wire N__28652;
    wire N__28649;
    wire N__28642;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28603;
    wire N__28600;
    wire N__28595;
    wire N__28590;
    wire N__28587;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28547;
    wire N__28546;
    wire N__28545;
    wire N__28542;
    wire N__28537;
    wire N__28534;
    wire N__28527;
    wire N__28524;
    wire N__28523;
    wire N__28522;
    wire N__28521;
    wire N__28518;
    wire N__28511;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28494;
    wire N__28493;
    wire N__28490;
    wire N__28489;
    wire N__28486;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28462;
    wire N__28461;
    wire N__28460;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28445;
    wire N__28444;
    wire N__28441;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28421;
    wire N__28416;
    wire N__28413;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28265;
    wire N__28264;
    wire N__28263;
    wire N__28262;
    wire N__28261;
    wire N__28260;
    wire N__28259;
    wire N__28246;
    wire N__28241;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28195;
    wire N__28194;
    wire N__28193;
    wire N__28192;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28160;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28109;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28098;
    wire N__28097;
    wire N__28096;
    wire N__28095;
    wire N__28094;
    wire N__28091;
    wire N__28090;
    wire N__28089;
    wire N__28088;
    wire N__28087;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28071;
    wire N__28070;
    wire N__28069;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28053;
    wire N__28050;
    wire N__28043;
    wire N__28036;
    wire N__28033;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28010;
    wire N__28009;
    wire N__28008;
    wire N__28007;
    wire N__28002;
    wire N__27997;
    wire N__27994;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27927;
    wire N__27924;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27869;
    wire N__27868;
    wire N__27865;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27841;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27825;
    wire N__27824;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27816;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27789;
    wire N__27788;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27751;
    wire N__27738;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27720;
    wire N__27717;
    wire N__27716;
    wire N__27715;
    wire N__27714;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27660;
    wire N__27659;
    wire N__27656;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27624;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27606;
    wire N__27605;
    wire N__27604;
    wire N__27603;
    wire N__27602;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27585;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27557;
    wire N__27554;
    wire N__27543;
    wire N__27540;
    wire N__27539;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27503;
    wire N__27498;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27476;
    wire N__27473;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27462;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27447;
    wire N__27442;
    wire N__27435;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27404;
    wire N__27401;
    wire N__27400;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27370;
    wire N__27363;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27319;
    wire N__27318;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27303;
    wire N__27298;
    wire N__27291;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27276;
    wire N__27273;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27250;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27222;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27180;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27169;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27161;
    wire N__27160;
    wire N__27155;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27126;
    wire N__27125;
    wire N__27124;
    wire N__27123;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27107;
    wire N__27102;
    wire N__27097;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27073;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27054;
    wire N__27053;
    wire N__27052;
    wire N__27051;
    wire N__27050;
    wire N__27049;
    wire N__27048;
    wire N__27047;
    wire N__27046;
    wire N__27045;
    wire N__27044;
    wire N__27043;
    wire N__27042;
    wire N__27039;
    wire N__27038;
    wire N__27037;
    wire N__27036;
    wire N__27033;
    wire N__27026;
    wire N__27023;
    wire N__27018;
    wire N__27017;
    wire N__27016;
    wire N__27011;
    wire N__27008;
    wire N__27007;
    wire N__27006;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26989;
    wire N__26986;
    wire N__26985;
    wire N__26980;
    wire N__26975;
    wire N__26970;
    wire N__26965;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26946;
    wire N__26943;
    wire N__26942;
    wire N__26941;
    wire N__26940;
    wire N__26939;
    wire N__26936;
    wire N__26931;
    wire N__26920;
    wire N__26915;
    wire N__26910;
    wire N__26907;
    wire N__26898;
    wire N__26883;
    wire N__26880;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26860;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26853;
    wire N__26850;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26808;
    wire N__26805;
    wire N__26800;
    wire N__26797;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26776;
    wire N__26775;
    wire N__26772;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26754;
    wire N__26753;
    wire N__26750;
    wire N__26749;
    wire N__26748;
    wire N__26747;
    wire N__26746;
    wire N__26745;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26698;
    wire N__26693;
    wire N__26690;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26674;
    wire N__26669;
    wire N__26664;
    wire N__26663;
    wire N__26662;
    wire N__26661;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26653;
    wire N__26652;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26569;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26555;
    wire N__26554;
    wire N__26553;
    wire N__26552;
    wire N__26551;
    wire N__26550;
    wire N__26549;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26538;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26523;
    wire N__26520;
    wire N__26519;
    wire N__26518;
    wire N__26515;
    wire N__26510;
    wire N__26509;
    wire N__26506;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26478;
    wire N__26475;
    wire N__26468;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26439;
    wire N__26438;
    wire N__26437;
    wire N__26436;
    wire N__26435;
    wire N__26434;
    wire N__26433;
    wire N__26432;
    wire N__26431;
    wire N__26430;
    wire N__26429;
    wire N__26426;
    wire N__26425;
    wire N__26424;
    wire N__26423;
    wire N__26422;
    wire N__26421;
    wire N__26420;
    wire N__26419;
    wire N__26418;
    wire N__26417;
    wire N__26416;
    wire N__26415;
    wire N__26414;
    wire N__26413;
    wire N__26412;
    wire N__26405;
    wire N__26404;
    wire N__26403;
    wire N__26398;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26377;
    wire N__26370;
    wire N__26365;
    wire N__26358;
    wire N__26353;
    wire N__26348;
    wire N__26345;
    wire N__26340;
    wire N__26335;
    wire N__26332;
    wire N__26317;
    wire N__26316;
    wire N__26315;
    wire N__26314;
    wire N__26313;
    wire N__26312;
    wire N__26311;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26291;
    wire N__26282;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26218;
    wire N__26217;
    wire N__26216;
    wire N__26215;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26207;
    wire N__26206;
    wire N__26205;
    wire N__26204;
    wire N__26199;
    wire N__26196;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26184;
    wire N__26179;
    wire N__26174;
    wire N__26173;
    wire N__26170;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26151;
    wire N__26148;
    wire N__26143;
    wire N__26130;
    wire N__26129;
    wire N__26126;
    wire N__26125;
    wire N__26124;
    wire N__26123;
    wire N__26120;
    wire N__26115;
    wire N__26112;
    wire N__26107;
    wire N__26106;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26091;
    wire N__26086;
    wire N__26083;
    wire N__26076;
    wire N__26073;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26065;
    wire N__26062;
    wire N__26059;
    wire N__26056;
    wire N__26055;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26043;
    wire N__26042;
    wire N__26041;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26029;
    wire N__26028;
    wire N__26025;
    wire N__26024;
    wire N__26021;
    wire N__26020;
    wire N__26019;
    wire N__26018;
    wire N__26017;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25980;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25953;
    wire N__25952;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25934;
    wire N__25931;
    wire N__25926;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25890;
    wire N__25885;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25875;
    wire N__25868;
    wire N__25861;
    wire N__25854;
    wire N__25851;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25829;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25818;
    wire N__25817;
    wire N__25816;
    wire N__25815;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25803;
    wire N__25798;
    wire N__25795;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25779;
    wire N__25776;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25743;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25726;
    wire N__25723;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25711;
    wire N__25708;
    wire N__25707;
    wire N__25704;
    wire N__25697;
    wire N__25694;
    wire N__25689;
    wire N__25684;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25665;
    wire N__25664;
    wire N__25663;
    wire N__25662;
    wire N__25659;
    wire N__25658;
    wire N__25655;
    wire N__25650;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25629;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25599;
    wire N__25596;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25551;
    wire N__25548;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25505;
    wire N__25504;
    wire N__25503;
    wire N__25502;
    wire N__25501;
    wire N__25500;
    wire N__25499;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25487;
    wire N__25486;
    wire N__25485;
    wire N__25484;
    wire N__25483;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25472;
    wire N__25469;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25459;
    wire N__25456;
    wire N__25451;
    wire N__25448;
    wire N__25443;
    wire N__25436;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25419;
    wire N__25408;
    wire N__25403;
    wire N__25392;
    wire N__25391;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25358;
    wire N__25357;
    wire N__25354;
    wire N__25353;
    wire N__25352;
    wire N__25351;
    wire N__25350;
    wire N__25349;
    wire N__25348;
    wire N__25347;
    wire N__25346;
    wire N__25341;
    wire N__25338;
    wire N__25329;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25307;
    wire N__25304;
    wire N__25299;
    wire N__25296;
    wire N__25295;
    wire N__25294;
    wire N__25293;
    wire N__25292;
    wire N__25291;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25277;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25266;
    wire N__25259;
    wire N__25256;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25231;
    wire N__25230;
    wire N__25229;
    wire N__25224;
    wire N__25219;
    wire N__25214;
    wire N__25209;
    wire N__25206;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25183;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25163;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25155;
    wire N__25154;
    wire N__25153;
    wire N__25150;
    wire N__25145;
    wire N__25142;
    wire N__25137;
    wire N__25128;
    wire N__25127;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25119;
    wire N__25118;
    wire N__25117;
    wire N__25112;
    wire N__25109;
    wire N__25108;
    wire N__25103;
    wire N__25100;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25075;
    wire N__25072;
    wire N__25067;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25055;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25047;
    wire N__25046;
    wire N__25045;
    wire N__25044;
    wire N__25041;
    wire N__25036;
    wire N__25031;
    wire N__25026;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24980;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24951;
    wire N__24948;
    wire N__24943;
    wire N__24940;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24812;
    wire N__24811;
    wire N__24810;
    wire N__24809;
    wire N__24808;
    wire N__24805;
    wire N__24804;
    wire N__24803;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24780;
    wire N__24777;
    wire N__24776;
    wire N__24775;
    wire N__24774;
    wire N__24773;
    wire N__24772;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24711;
    wire N__24708;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24658;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24639;
    wire N__24634;
    wire N__24627;
    wire N__24624;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24616;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24605;
    wire N__24602;
    wire N__24597;
    wire N__24594;
    wire N__24593;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24586;
    wire N__24585;
    wire N__24584;
    wire N__24583;
    wire N__24582;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24493;
    wire N__24492;
    wire N__24489;
    wire N__24484;
    wire N__24469;
    wire N__24460;
    wire N__24459;
    wire N__24456;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24414;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24368;
    wire N__24367;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24359;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24345;
    wire N__24342;
    wire N__24337;
    wire N__24334;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24313;
    wire N__24306;
    wire N__24305;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24281;
    wire N__24280;
    wire N__24279;
    wire N__24276;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24254;
    wire N__24251;
    wire N__24240;
    wire N__24239;
    wire N__24238;
    wire N__24237;
    wire N__24236;
    wire N__24235;
    wire N__24234;
    wire N__24233;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24225;
    wire N__24224;
    wire N__24223;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24206;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24153;
    wire N__24150;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24129;
    wire N__24126;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24110;
    wire N__24109;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24081;
    wire N__24072;
    wire N__24071;
    wire N__24068;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24023;
    wire N__24020;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23969;
    wire N__23968;
    wire N__23965;
    wire N__23964;
    wire N__23963;
    wire N__23962;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23947;
    wire N__23946;
    wire N__23943;
    wire N__23942;
    wire N__23939;
    wire N__23938;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23840;
    wire N__23837;
    wire N__23832;
    wire N__23829;
    wire N__23826;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23791;
    wire N__23784;
    wire N__23783;
    wire N__23782;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23766;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23748;
    wire N__23743;
    wire N__23740;
    wire N__23735;
    wire N__23730;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23706;
    wire N__23705;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23687;
    wire N__23684;
    wire N__23683;
    wire N__23682;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23667;
    wire N__23666;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23637;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23629;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23537;
    wire N__23536;
    wire N__23533;
    wire N__23526;
    wire N__23519;
    wire N__23518;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23510;
    wire N__23507;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23478;
    wire N__23469;
    wire N__23468;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23381;
    wire N__23378;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23355;
    wire N__23354;
    wire N__23353;
    wire N__23352;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23341;
    wire N__23338;
    wire N__23337;
    wire N__23336;
    wire N__23335;
    wire N__23334;
    wire N__23331;
    wire N__23330;
    wire N__23329;
    wire N__23328;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23220;
    wire N__23217;
    wire N__23210;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23186;
    wire N__23185;
    wire N__23184;
    wire N__23183;
    wire N__23182;
    wire N__23181;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23158;
    wire N__23155;
    wire N__23142;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23127;
    wire N__23124;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23112;
    wire N__23111;
    wire N__23110;
    wire N__23109;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23094;
    wire N__23093;
    wire N__23090;
    wire N__23089;
    wire N__23088;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23055;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23011;
    wire N__23008;
    wire N__23001;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22958;
    wire N__22951;
    wire N__22948;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22926;
    wire N__22925;
    wire N__22924;
    wire N__22921;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22887;
    wire N__22884;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22872;
    wire N__22869;
    wire N__22868;
    wire N__22865;
    wire N__22864;
    wire N__22863;
    wire N__22860;
    wire N__22859;
    wire N__22858;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22854;
    wire N__22853;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22801;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22745;
    wire N__22742;
    wire N__22737;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22703;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22691;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22651;
    wire N__22646;
    wire N__22639;
    wire N__22626;
    wire N__22625;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22604;
    wire N__22603;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22592;
    wire N__22591;
    wire N__22588;
    wire N__22587;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22570;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22559;
    wire N__22558;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22554;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22459;
    wire N__22456;
    wire N__22449;
    wire N__22448;
    wire N__22443;
    wire N__22438;
    wire N__22431;
    wire N__22428;
    wire N__22423;
    wire N__22422;
    wire N__22421;
    wire N__22420;
    wire N__22415;
    wire N__22412;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22371;
    wire N__22368;
    wire N__22367;
    wire N__22366;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22358;
    wire N__22357;
    wire N__22356;
    wire N__22353;
    wire N__22352;
    wire N__22349;
    wire N__22348;
    wire N__22347;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22335;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22309;
    wire N__22306;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22231;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22212;
    wire N__22205;
    wire N__22204;
    wire N__22203;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22170;
    wire N__22165;
    wire N__22160;
    wire N__22153;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22128;
    wire N__22127;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22099;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22088;
    wire N__22085;
    wire N__22084;
    wire N__22083;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22071;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22060;
    wire N__22059;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22047;
    wire N__22046;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21956;
    wire N__21951;
    wire N__21948;
    wire N__21947;
    wire N__21944;
    wire N__21937;
    wire N__21936;
    wire N__21935;
    wire N__21928;
    wire N__21925;
    wire N__21920;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21894;
    wire N__21885;
    wire N__21884;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21767;
    wire N__21766;
    wire N__21765;
    wire N__21764;
    wire N__21763;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21753;
    wire N__21750;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21734;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21662;
    wire N__21661;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21520;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21495;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21474;
    wire N__21471;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21447;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21393;
    wire N__21384;
    wire N__21383;
    wire N__21378;
    wire N__21375;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21336;
    wire N__21335;
    wire N__21334;
    wire N__21331;
    wire N__21326;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21258;
    wire N__21257;
    wire N__21256;
    wire N__21249;
    wire N__21246;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21202;
    wire N__21199;
    wire N__21194;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21174;
    wire N__21171;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21135;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21069;
    wire N__21068;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21041;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20996;
    wire N__20995;
    wire N__20994;
    wire N__20993;
    wire N__20992;
    wire N__20989;
    wire N__20988;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20980;
    wire N__20977;
    wire N__20976;
    wire N__20973;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20962;
    wire N__20961;
    wire N__20958;
    wire N__20957;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20782;
    wire N__20775;
    wire N__20768;
    wire N__20759;
    wire N__20754;
    wire N__20751;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20718;
    wire N__20715;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20670;
    wire N__20669;
    wire N__20666;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20651;
    wire N__20646;
    wire N__20643;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20625;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20617;
    wire N__20612;
    wire N__20607;
    wire N__20604;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20593;
    wire N__20590;
    wire N__20589;
    wire N__20586;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20547;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20496;
    wire N__20493;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20481;
    wire N__20478;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20442;
    wire N__20439;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20221;
    wire N__20216;
    wire N__20215;
    wire N__20214;
    wire N__20213;
    wire N__20212;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20192;
    wire N__20189;
    wire N__20188;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20159;
    wire N__20158;
    wire N__20157;
    wire N__20156;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20144;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20105;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20080;
    wire N__20075;
    wire N__20072;
    wire N__20067;
    wire N__20064;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19897;
    wire N__19896;
    wire N__19891;
    wire N__19886;
    wire N__19881;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19716;
    wire N__19715;
    wire N__19712;
    wire N__19711;
    wire N__19710;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19696;
    wire N__19689;
    wire N__19688;
    wire N__19685;
    wire N__19684;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19673;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19665;
    wire N__19662;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19508;
    wire N__19507;
    wire N__19506;
    wire N__19505;
    wire N__19502;
    wire N__19501;
    wire N__19492;
    wire N__19487;
    wire N__19486;
    wire N__19485;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19470;
    wire N__19469;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19229;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19215;
    wire N__19214;
    wire N__19213;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19183;
    wire N__19182;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19041;
    wire N__19038;
    wire N__19031;
    wire N__19028;
    wire N__19023;
    wire N__19020;
    wire N__19013;
    wire N__19008;
    wire N__18999;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18950;
    wire N__18947;
    wire N__18946;
    wire N__18945;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18922;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18882;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18857;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18849;
    wire N__18846;
    wire N__18841;
    wire N__18838;
    wire N__18831;
    wire N__18830;
    wire N__18829;
    wire N__18828;
    wire N__18827;
    wire N__18826;
    wire N__18823;
    wire N__18816;
    wire N__18811;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18787;
    wire N__18786;
    wire N__18779;
    wire N__18778;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18766;
    wire N__18759;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18662;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18645;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18605;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18582;
    wire N__18581;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18506;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18495;
    wire N__18494;
    wire N__18493;
    wire N__18492;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18481;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18467;
    wire N__18466;
    wire N__18465;
    wire N__18464;
    wire N__18461;
    wire N__18460;
    wire N__18459;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18369;
    wire N__18366;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18338;
    wire N__18333;
    wire N__18330;
    wire N__18329;
    wire N__18328;
    wire N__18327;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18316;
    wire N__18313;
    wire N__18312;
    wire N__18309;
    wire N__18308;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18281;
    wire N__18280;
    wire N__18279;
    wire N__18276;
    wire N__18275;
    wire N__18274;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18226;
    wire N__18221;
    wire N__18218;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18178;
    wire N__18175;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18155;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18137;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18116;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18112;
    wire N__18111;
    wire N__18110;
    wire N__18107;
    wire N__18106;
    wire N__18103;
    wire N__18102;
    wire N__18101;
    wire N__18100;
    wire N__18099;
    wire N__18098;
    wire N__18095;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18082;
    wire N__18079;
    wire N__18076;
    wire N__18073;
    wire N__18070;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17940;
    wire N__17935;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17897;
    wire N__17894;
    wire N__17887;
    wire N__17884;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17834;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17810;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17781;
    wire N__17780;
    wire N__17777;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17760;
    wire N__17759;
    wire N__17758;
    wire N__17757;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17749;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17733;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17697;
    wire N__17688;
    wire N__17687;
    wire N__17686;
    wire N__17685;
    wire N__17684;
    wire N__17683;
    wire N__17682;
    wire N__17681;
    wire N__17678;
    wire N__17677;
    wire N__17676;
    wire N__17675;
    wire N__17674;
    wire N__17673;
    wire N__17672;
    wire N__17671;
    wire N__17670;
    wire N__17669;
    wire N__17664;
    wire N__17659;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17639;
    wire N__17632;
    wire N__17629;
    wire N__17628;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17616;
    wire N__17615;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17601;
    wire N__17596;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17574;
    wire N__17565;
    wire N__17562;
    wire N__17561;
    wire N__17560;
    wire N__17557;
    wire N__17556;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17548;
    wire N__17545;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17522;
    wire N__17517;
    wire N__17516;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17501;
    wire N__17498;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17439;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17423;
    wire N__17422;
    wire N__17421;
    wire N__17418;
    wire N__17413;
    wire N__17412;
    wire N__17411;
    wire N__17408;
    wire N__17407;
    wire N__17406;
    wire N__17401;
    wire N__17396;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17327;
    wire N__17326;
    wire N__17325;
    wire N__17324;
    wire N__17323;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17315;
    wire N__17314;
    wire N__17313;
    wire N__17312;
    wire N__17311;
    wire N__17310;
    wire N__17309;
    wire N__17308;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17303;
    wire N__17302;
    wire N__17299;
    wire N__17294;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17282;
    wire N__17281;
    wire N__17280;
    wire N__17277;
    wire N__17272;
    wire N__17265;
    wire N__17260;
    wire N__17259;
    wire N__17250;
    wire N__17245;
    wire N__17244;
    wire N__17243;
    wire N__17242;
    wire N__17241;
    wire N__17240;
    wire N__17229;
    wire N__17222;
    wire N__17219;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17181;
    wire N__17166;
    wire N__17165;
    wire N__17164;
    wire N__17163;
    wire N__17162;
    wire N__17161;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17153;
    wire N__17144;
    wire N__17143;
    wire N__17142;
    wire N__17141;
    wire N__17140;
    wire N__17139;
    wire N__17138;
    wire N__17135;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17119;
    wire N__17118;
    wire N__17115;
    wire N__17114;
    wire N__17109;
    wire N__17106;
    wire N__17101;
    wire N__17094;
    wire N__17091;
    wire N__17086;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17063;
    wire N__17062;
    wire N__17059;
    wire N__17058;
    wire N__17053;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17029;
    wire N__17028;
    wire N__17027;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17012;
    wire N__17009;
    wire N__17004;
    wire N__17001;
    wire N__16986;
    wire N__16985;
    wire N__16984;
    wire N__16983;
    wire N__16982;
    wire N__16981;
    wire N__16980;
    wire N__16977;
    wire N__16974;
    wire N__16973;
    wire N__16972;
    wire N__16971;
    wire N__16970;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16962;
    wire N__16961;
    wire N__16958;
    wire N__16957;
    wire N__16954;
    wire N__16953;
    wire N__16952;
    wire N__16949;
    wire N__16948;
    wire N__16947;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16932;
    wire N__16931;
    wire N__16924;
    wire N__16919;
    wire N__16914;
    wire N__16911;
    wire N__16910;
    wire N__16909;
    wire N__16908;
    wire N__16903;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16871;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16848;
    wire N__16843;
    wire N__16832;
    wire N__16821;
    wire N__16820;
    wire N__16819;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16811;
    wire N__16810;
    wire N__16809;
    wire N__16806;
    wire N__16799;
    wire N__16796;
    wire N__16795;
    wire N__16794;
    wire N__16793;
    wire N__16792;
    wire N__16791;
    wire N__16790;
    wire N__16789;
    wire N__16788;
    wire N__16785;
    wire N__16784;
    wire N__16783;
    wire N__16780;
    wire N__16779;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16767;
    wire N__16766;
    wire N__16765;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16757;
    wire N__16756;
    wire N__16755;
    wire N__16754;
    wire N__16751;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16738;
    wire N__16733;
    wire N__16732;
    wire N__16729;
    wire N__16722;
    wire N__16721;
    wire N__16720;
    wire N__16719;
    wire N__16718;
    wire N__16711;
    wire N__16708;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16690;
    wire N__16683;
    wire N__16676;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16640;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16619;
    wire N__16608;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16592;
    wire N__16591;
    wire N__16590;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16582;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16563;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16506;
    wire N__16505;
    wire N__16502;
    wire N__16501;
    wire N__16500;
    wire N__16499;
    wire N__16496;
    wire N__16495;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16478;
    wire N__16477;
    wire N__16476;
    wire N__16473;
    wire N__16472;
    wire N__16469;
    wire N__16468;
    wire N__16467;
    wire N__16466;
    wire N__16461;
    wire N__16456;
    wire N__16453;
    wire N__16448;
    wire N__16447;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16432;
    wire N__16427;
    wire N__16418;
    wire N__16411;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16377;
    wire N__16376;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16368;
    wire N__16367;
    wire N__16366;
    wire N__16365;
    wire N__16364;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16339;
    wire N__16336;
    wire N__16335;
    wire N__16332;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16303;
    wire N__16302;
    wire N__16301;
    wire N__16298;
    wire N__16291;
    wire N__16284;
    wire N__16279;
    wire N__16274;
    wire N__16271;
    wire N__16260;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16250;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16235;
    wire N__16234;
    wire N__16233;
    wire N__16230;
    wire N__16225;
    wire N__16224;
    wire N__16223;
    wire N__16222;
    wire N__16219;
    wire N__16218;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16170;
    wire N__16167;
    wire N__16166;
    wire N__16165;
    wire N__16162;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16148;
    wire N__16143;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16125;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16121;
    wire N__16116;
    wire N__16115;
    wire N__16114;
    wire N__16111;
    wire N__16110;
    wire N__16109;
    wire N__16108;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16094;
    wire N__16093;
    wire N__16092;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16080;
    wire N__16075;
    wire N__16068;
    wire N__16065;
    wire N__16060;
    wire N__16055;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16029;
    wire N__16028;
    wire N__16027;
    wire N__16026;
    wire N__16023;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16002;
    wire N__15999;
    wire N__15996;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15992;
    wire N__15989;
    wire N__15988;
    wire N__15987;
    wire N__15986;
    wire N__15985;
    wire N__15978;
    wire N__15975;
    wire N__15972;
    wire N__15969;
    wire N__15962;
    wire N__15951;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15908;
    wire N__15907;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15882;
    wire N__15877;
    wire N__15870;
    wire N__15867;
    wire N__15864;
    wire N__15861;
    wire N__15860;
    wire N__15859;
    wire N__15856;
    wire N__15851;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15827;
    wire N__15826;
    wire N__15825;
    wire N__15822;
    wire N__15819;
    wire N__15818;
    wire N__15815;
    wire N__15814;
    wire N__15811;
    wire N__15810;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15798;
    wire N__15795;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15785;
    wire N__15780;
    wire N__15775;
    wire N__15772;
    wire N__15759;
    wire N__15756;
    wire N__15753;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15728;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15703;
    wire N__15698;
    wire N__15695;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15677;
    wire N__15674;
    wire N__15673;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15656;
    wire N__15655;
    wire N__15654;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15636;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15622;
    wire N__15617;
    wire N__15614;
    wire N__15603;
    wire N__15600;
    wire N__15599;
    wire N__15598;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15581;
    wire N__15580;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15568;
    wire N__15567;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15552;
    wire N__15549;
    wire N__15544;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15518;
    wire N__15517;
    wire N__15516;
    wire N__15513;
    wire N__15508;
    wire N__15505;
    wire N__15498;
    wire N__15495;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15468;
    wire N__15465;
    wire N__15464;
    wire N__15461;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15428;
    wire N__15427;
    wire N__15426;
    wire N__15423;
    wire N__15418;
    wire N__15415;
    wire N__15408;
    wire N__15407;
    wire N__15406;
    wire N__15405;
    wire N__15398;
    wire N__15395;
    wire N__15394;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15386;
    wire N__15385;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15362;
    wire N__15351;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15332;
    wire N__15331;
    wire N__15328;
    wire N__15327;
    wire N__15326;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15318;
    wire N__15317;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15299;
    wire N__15294;
    wire N__15291;
    wire N__15276;
    wire N__15273;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15265;
    wire N__15264;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15256;
    wire N__15255;
    wire N__15254;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15239;
    wire N__15236;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15220;
    wire N__15215;
    wire N__15212;
    wire N__15201;
    wire N__15198;
    wire N__15197;
    wire N__15196;
    wire N__15195;
    wire N__15192;
    wire N__15191;
    wire N__15190;
    wire N__15187;
    wire N__15182;
    wire N__15181;
    wire N__15180;
    wire N__15179;
    wire N__15178;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15129;
    wire N__15126;
    wire N__15125;
    wire N__15124;
    wire N__15121;
    wire N__15120;
    wire N__15119;
    wire N__15116;
    wire N__15115;
    wire N__15114;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15097;
    wire N__15092;
    wire N__15083;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15065;
    wire N__15064;
    wire N__15063;
    wire N__15060;
    wire N__15059;
    wire N__15058;
    wire N__15057;
    wire N__15056;
    wire N__15055;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15037;
    wire N__15028;
    wire N__15023;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14987;
    wire N__14986;
    wire N__14985;
    wire N__14982;
    wire N__14981;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14973;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14948;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14944;
    wire N__14939;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14901;
    wire N__14896;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14876;
    wire N__14875;
    wire N__14874;
    wire N__14873;
    wire N__14872;
    wire N__14869;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14847;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14826;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14798;
    wire N__14797;
    wire N__14794;
    wire N__14793;
    wire N__14792;
    wire N__14791;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14772;
    wire N__14771;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14759;
    wire N__14754;
    wire N__14753;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14742;
    wire N__14741;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14721;
    wire N__14718;
    wire N__14713;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14673;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14646;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14630;
    wire N__14627;
    wire N__14626;
    wire N__14625;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14610;
    wire N__14605;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14537;
    wire N__14536;
    wire N__14533;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14499;
    wire N__14498;
    wire N__14497;
    wire N__14496;
    wire N__14495;
    wire N__14494;
    wire N__14493;
    wire N__14492;
    wire N__14489;
    wire N__14488;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14474;
    wire N__14467;
    wire N__14462;
    wire N__14459;
    wire N__14454;
    wire N__14439;
    wire N__14436;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14418;
    wire N__14415;
    wire N__14412;
    wire N__14409;
    wire N__14406;
    wire N__14403;
    wire N__14400;
    wire N__14397;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14385;
    wire N__14382;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14367;
    wire N__14366;
    wire N__14365;
    wire N__14364;
    wire N__14361;
    wire N__14356;
    wire N__14355;
    wire N__14354;
    wire N__14353;
    wire N__14350;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14334;
    wire N__14331;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14313;
    wire N__14310;
    wire N__14307;
    wire N__14304;
    wire N__14301;
    wire N__14300;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14255;
    wire N__14254;
    wire N__14251;
    wire N__14246;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14234;
    wire N__14229;
    wire N__14226;
    wire N__14221;
    wire N__14214;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14206;
    wire N__14205;
    wire N__14200;
    wire N__14197;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14185;
    wire N__14178;
    wire N__14177;
    wire N__14172;
    wire N__14169;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14157;
    wire N__14156;
    wire N__14155;
    wire N__14154;
    wire N__14151;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14122;
    wire N__14119;
    wire N__14114;
    wire N__14109;
    wire N__14108;
    wire N__14107;
    wire N__14106;
    wire N__14105;
    wire N__14104;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14033;
    wire N__14032;
    wire N__14027;
    wire N__14024;
    wire N__14019;
    wire N__14016;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14008;
    wire N__14007;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13992;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13952;
    wire N__13951;
    wire N__13948;
    wire N__13943;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13922;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13908;
    wire N__13905;
    wire N__13900;
    wire N__13899;
    wire N__13898;
    wire N__13897;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13880;
    wire N__13877;
    wire N__13866;
    wire N__13865;
    wire N__13860;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13811;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13794;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13779;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13771;
    wire N__13770;
    wire N__13769;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13757;
    wire N__13752;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13724;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13694;
    wire N__13693;
    wire N__13690;
    wire N__13685;
    wire N__13680;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13668;
    wire N__13667;
    wire N__13666;
    wire N__13665;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13651;
    wire N__13644;
    wire N__13641;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13629;
    wire N__13628;
    wire N__13627;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13615;
    wire N__13608;
    wire N__13607;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13597;
    wire N__13590;
    wire N__13589;
    wire N__13588;
    wire N__13587;
    wire N__13580;
    wire N__13577;
    wire N__13572;
    wire N__13569;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13557;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13545;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13521;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13499;
    wire N__13498;
    wire N__13497;
    wire N__13496;
    wire N__13495;
    wire N__13494;
    wire N__13489;
    wire N__13486;
    wire N__13483;
    wire N__13478;
    wire N__13475;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13434;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13406;
    wire N__13405;
    wire N__13404;
    wire N__13403;
    wire N__13398;
    wire N__13393;
    wire N__13390;
    wire N__13383;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13375;
    wire N__13370;
    wire N__13367;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13355;
    wire N__13354;
    wire N__13351;
    wire N__13346;
    wire N__13343;
    wire N__13338;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13262;
    wire N__13261;
    wire N__13260;
    wire N__13259;
    wire N__13258;
    wire N__13255;
    wire N__13250;
    wire N__13243;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13208;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13127;
    wire N__13126;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13118;
    wire N__13117;
    wire N__13114;
    wire N__13113;
    wire N__13112;
    wire N__13111;
    wire N__13108;
    wire N__13107;
    wire N__13106;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13086;
    wire N__13083;
    wire N__13082;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13037;
    wire N__13036;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13014;
    wire N__13009;
    wire N__13006;
    wire N__13003;
    wire N__13000;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12979;
    wire N__12972;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12953;
    wire N__12948;
    wire N__12945;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12896;
    wire N__12895;
    wire N__12894;
    wire N__12893;
    wire N__12892;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12880;
    wire N__12877;
    wire N__12872;
    wire N__12861;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12843;
    wire N__12840;
    wire N__12839;
    wire N__12836;
    wire N__12835;
    wire N__12832;
    wire N__12825;
    wire N__12822;
    wire N__12821;
    wire N__12820;
    wire N__12817;
    wire N__12812;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12719;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12704;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12632;
    wire N__12631;
    wire N__12628;
    wire N__12623;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12468;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12456;
    wire N__12453;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12441;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12433;
    wire N__12432;
    wire N__12431;
    wire N__12430;
    wire N__12425;
    wire N__12416;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12404;
    wire N__12403;
    wire N__12400;
    wire N__12399;
    wire N__12398;
    wire N__12397;
    wire N__12392;
    wire N__12383;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12371;
    wire N__12370;
    wire N__12369;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12357;
    wire N__12350;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12338;
    wire N__12337;
    wire N__12336;
    wire N__12335;
    wire N__12334;
    wire N__12329;
    wire N__12320;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12302;
    wire N__12297;
    wire N__12294;
    wire N__12293;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12276;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12268;
    wire N__12263;
    wire N__12262;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12244;
    wire N__12241;
    wire N__12236;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12174;
    wire N__12171;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11861;
    wire N__11858;
    wire N__11855;
    wire N__11852;
    wire N__11847;
    wire N__11844;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire VCCG0;
    wire GNDG0;
    wire port_data_rw_i_i;
    wire port_nmib_0_i;
    wire this_vga_signals_vvisibility_i;
    wire rgb_c_2;
    wire rgb_c_1;
    wire rgb_c_4;
    wire M_this_map_ram_write_data_4;
    wire N_393_0;
    wire rgb_c_3;
    wire M_this_map_address_qZ0Z_0;
    wire bfn_10_27_0_;
    wire M_this_map_address_qZ0Z_1;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire un1_M_this_map_address_q_cry_1;
    wire M_this_map_address_qZ0Z_3;
    wire un1_M_this_map_address_q_cry_2;
    wire M_this_map_address_qZ0Z_4;
    wire un1_M_this_map_address_q_cry_3;
    wire M_this_map_address_qZ0Z_5;
    wire un1_M_this_map_address_q_cry_4;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_5;
    wire M_this_map_address_qZ0Z_7;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire M_this_map_address_qZ0Z_8;
    wire bfn_10_28_0_;
    wire un1_M_this_map_address_q_cry_8;
    wire M_this_map_address_qZ0Z_9;
    wire rgb_c_0;
    wire \this_vga_ramdac.i2_mux_cascade_ ;
    wire \this_vga_ramdac.N_3300_reto ;
    wire \this_vga_ramdac.m6_cascade_ ;
    wire \this_vga_ramdac.N_3299_reto ;
    wire rgb_c_5;
    wire \this_vga_signals.N_729 ;
    wire N_495;
    wire \this_vga_signals.un2_vsynclt8_cascade_ ;
    wire this_vga_signals_vsync_1_i;
    wire \this_vga_signals.vsync_1_2 ;
    wire \this_vga_signals.vsync_1_3 ;
    wire \this_vga_signals.mult1_un47_sum_c3_1_1_0_cascade_ ;
    wire \this_vga_signals.vaddress_5_0_6 ;
    wire \this_vga_signals.N_5 ;
    wire \this_vga_signals.if_m8_0_a3_1_1_0 ;
    wire \this_vga_signals.g2_5 ;
    wire \this_vga_signals.N_18_0 ;
    wire \this_vga_signals.g0_7_0_cascade_ ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire \this_vga_signals.N_4_0_0_cascade_ ;
    wire \this_vga_signals.if_m8_0_a3_1_1_1 ;
    wire \this_vga_signals.if_N_5_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3_1_1_0 ;
    wire \this_vga_ramdac.N_3301_reto ;
    wire \this_vga_signals.vvisibility_1_cascade_ ;
    wire \this_vga_ramdac.m16 ;
    wire \this_vga_ramdac.m19_cascade_ ;
    wire \this_vga_ramdac.N_3302_reto ;
    wire \this_vga_ramdac.N_3303_reto ;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_3;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_1;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire this_pixel_clk_M_counter_q_i_1;
    wire this_pixel_clk_M_counter_q_0;
    wire \this_vga_ramdac.N_880_i_reto ;
    wire N_880_0_cascade_;
    wire M_this_vga_signals_address_5;
    wire M_this_vga_signals_address_3;
    wire M_this_vga_signals_address_4;
    wire port_clk_c;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire M_this_map_ram_write_data_1;
    wire M_this_map_ram_write_data_5;
    wire bfn_13_12_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_13_13_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_0 ;
    wire \this_vga_signals.if_i1_mux_0_cascade_ ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.N_5_i_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3 ;
    wire \this_vga_signals.N_3_2_0_1 ;
    wire \this_vga_signals.g0_i_x4_0_0_cascade_ ;
    wire \this_vga_signals.N_3_3_0_0 ;
    wire \this_vga_signals.g0_0_2_0_0_cascade_ ;
    wire \this_vga_signals.g0_6_2 ;
    wire \this_vga_signals.g1_1_0_0_0_cascade_ ;
    wire \this_vga_signals.N_5_i_1_0_0 ;
    wire \this_vga_signals.g0_2_1_cascade_ ;
    wire \this_vga_signals.N_5_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_x1 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_x0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_ns_cascade_ ;
    wire \this_vga_signals.g0_31_N_4L6 ;
    wire \this_vga_signals.g0_31_N_2L1_cascade_ ;
    wire \this_vga_signals.g0_31_N_5L8 ;
    wire \this_vga_signals.M_pcounter_q_3_0_cascade_ ;
    wire \this_vga_signals.N_2_0_cascade_ ;
    wire \this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_d7lt3_cascade_ ;
    wire \this_vga_ramdac.N_24_mux ;
    wire M_pcounter_q_ret_2_RNIH7PG8;
    wire \this_vga_ramdac.N_3298_reto ;
    wire \this_vga_signals.M_pcounter_q_3_1_cascade_ ;
    wire \this_vga_signals.M_pcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_1_cascade_ ;
    wire M_this_vga_signals_address_0;
    wire N_880_0;
    wire M_this_vga_signals_address_2;
    wire \this_vga_signals.mult1_un82_sum_c2_0 ;
    wire \this_vga_signals.mult1_un82_sum_c2_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_c3_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_2_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_2_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1 ;
    wire M_this_oam_ram_read_data_4;
    wire M_this_map_ram_read_data_4;
    wire M_this_ppu_sprites_addr_10;
    wire M_this_map_ram_write_data_0;
    wire M_this_map_ram_write_data_7;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.N_1_4_1_cascade_ ;
    wire \this_vga_signals.SUM_2_i_1_2_3_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.g0_0_0_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0 ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0 ;
    wire \this_vga_signals.if_i2_mux ;
    wire \this_vga_signals.g0_1_1_x0_cascade_ ;
    wire \this_vga_signals.g0_1_1_cascade_ ;
    wire \this_vga_signals.N_4_0_0_0 ;
    wire \this_vga_signals.g0_0_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_x0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0 ;
    wire \this_vga_signals.g1_5_cascade_ ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_x1 ;
    wire \this_vga_signals.g1_2 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_ns ;
    wire \this_vga_signals.mult1_un68_sum_axb1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c2_0 ;
    wire \this_vga_signals.N_3_0 ;
    wire \this_vga_signals.M_pcounter_q_i_3_1 ;
    wire \this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_ ;
    wire \this_vga_signals.N_2_0 ;
    wire \this_vga_signals.M_pcounter_q_i_3_0 ;
    wire \this_vga_signals.M_hcounter_d7lt7_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_d7_0_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un89_sum_c3 ;
    wire \this_vga_signals.mult1_un75_sum_c2_0 ;
    wire \this_vga_signals.mult1_un75_sum_c2_0_cascade_ ;
    wire \this_vga_signals.if_N_9_1 ;
    wire \this_vga_signals.if_m7_0_x4_0 ;
    wire \this_vga_signals.mult1_un75_sum_c3 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_2 ;
    wire \this_vga_signals.mult1_un75_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire \this_vga_signals.SUM_3_i_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_0_1_cascade_ ;
    wire \this_vga_signals.if_N_8_i_0 ;
    wire \this_vga_signals.M_hcounter_d7lto7_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0 ;
    wire M_hcounter_q_esr_RNIR18F4_9;
    wire \this_vga_signals.N_473_0_cascade_ ;
    wire \this_vga_signals.N_554 ;
    wire \this_vga_signals.SUM_3_i_1_0 ;
    wire \this_vga_signals.N_735_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_2_cascade_ ;
    wire \this_vga_signals.N_735_0 ;
    wire \this_vga_signals.mult1_un61_sum_0_3 ;
    wire \this_vga_signals.hsync_1_i_0_1 ;
    wire \this_vga_signals.N_507_0 ;
    wire M_this_map_ram_write_data_6;
    wire \this_vga_signals.M_lcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_lcounter_d_0_sqmuxa ;
    wire \this_vga_signals.M_hcounter_d7_0 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.N_966_0 ;
    wire \this_vga_signals.N_1332_g ;
    wire \this_vga_signals.g1_0_0_0_0 ;
    wire \this_vga_signals.g0_2_2_1 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_2 ;
    wire \this_vga_signals.vaddress_3_6 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_2_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3_2 ;
    wire \this_vga_signals.mult1_un47_sum_c3_2_cascade_ ;
    wire \this_vga_signals.g0_1 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.vaddress_6_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_i ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un47_sum_c3 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_654_x0 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_654_x1 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_654_ns_cascade_ ;
    wire \this_vga_signals.if_m1_3 ;
    wire \this_vga_signals.if_m1_3_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1 ;
    wire \this_vga_signals.vaddress_0_6 ;
    wire \this_vga_signals.mult1_un47_sum_c3_1_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.g0_2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0_1 ;
    wire \this_vga_signals.N_3_1_0 ;
    wire \this_vga_signals.N_11_0_0_cascade_ ;
    wire \this_vga_signals.N_4_1_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.mult1_un68_sum_axb1 ;
    wire \this_vga_signals.if_m5_s ;
    wire \this_vga_signals.M_vcounter_d7lto8_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ;
    wire \this_vga_signals.M_hcounter_d7lto4_0 ;
    wire \this_sprites_ram.mem_out_bus7_0 ;
    wire \this_sprites_ram.mem_out_bus3_0 ;
    wire bfn_15_20_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_15_21_0_;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.N_966_1 ;
    wire \this_sprites_ram.mem_WE_8 ;
    wire M_this_map_ram_write_data_2;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.g0_0_0_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.g2_0_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.g0_2_0 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_0 ;
    wire \this_vga_signals.SUM_2_i_1_0_3 ;
    wire \this_vga_signals.SUM_2_i_1_2_3 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.vaddress_0_0_6_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i ;
    wire \this_vga_signals.mult1_un54_sum_c3_1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1_654_ns ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ;
    wire \this_vga_signals.g0_i_i_a5_1_0_0_0 ;
    wire \this_vga_signals.g0_i_i_0_0_0 ;
    wire \this_vga_signals.vaddress_2_6_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0_0 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.mult1_un47_sum_c3_0 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i_0_0 ;
    wire \this_vga_signals.N_7_1_0 ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.vaddress_0_0_6 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_1 ;
    wire \this_vga_signals.g0_0_0 ;
    wire \this_ppu.un13_0_cascade_ ;
    wire \this_ppu.M_line_clk_out_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_d7lt9_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.un4_lvisibility_1 ;
    wire \this_vga_signals.line_clk_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire \this_vga_signals.un4_lvisibility_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire M_this_vga_signals_line_clk_0_cascade_;
    wire bfn_16_17_0_;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_6_s1 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_7 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_2 ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_4 ;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.GZ0Z_394 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_vcounter_q_501_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_sprites_ram.mem_WE_10 ;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_7_cascade_ ;
    wire N_597_cascade_;
    wire M_this_sprites_address_qc_7_0;
    wire N_1298_tz_0;
    wire N_1294_tz_0;
    wire N_602_cascade_;
    wire M_this_sprites_address_qc_8_0;
    wire M_this_map_ram_write_data_3;
    wire M_this_oam_ram_read_data_2;
    wire M_this_map_ram_read_data_2;
    wire M_this_ppu_sprites_addr_8;
    wire M_this_ppu_sprites_addr_5;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire M_this_ppu_sprites_addr_4;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_ppu.M_state_q_srsts_i_2_1_cascade_ ;
    wire \this_ppu.M_count_qZ0Z_6 ;
    wire \this_ppu.M_count_qZ0Z_7 ;
    wire \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5_cascade_ ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_5 ;
    wire \this_ppu.M_count_qZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_8 ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5 ;
    wire \this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4 ;
    wire \this_ppu.M_count_d_0_sqmuxa_1 ;
    wire \this_ppu.M_count_d_0_sqmuxa_1_cascade_ ;
    wire \this_ppu.M_line_clk_out_0 ;
    wire \this_ppu.N_1417_0 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ;
    wire \this_ppu.N_1417_0_cascade_ ;
    wire \this_ppu.un13_0 ;
    wire \this_ppu.M_count_qZ0Z_3 ;
    wire \this_sprites_ram.mem_out_bus6_2 ;
    wire \this_sprites_ram.mem_out_bus2_2 ;
    wire \this_reset_cond.M_stage_qZ0Z_3 ;
    wire \this_reset_cond.M_stage_qZ0Z_6 ;
    wire \this_reset_cond.M_stage_qZ0Z_7 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_4 ;
    wire \this_reset_cond.M_stage_qZ0Z_5 ;
    wire \this_sprites_ram.mem_out_bus6_0 ;
    wire \this_sprites_ram.mem_out_bus2_0 ;
    wire M_this_map_ram_read_data_5;
    wire M_this_oam_ram_read_data_5;
    wire M_this_map_ram_read_data_7;
    wire M_this_oam_ram_read_data_7;
    wire \this_sprites_ram.mem_out_bus4_2 ;
    wire \this_sprites_ram.mem_out_bus0_2 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ;
    wire M_this_oam_ram_read_data_3;
    wire M_this_map_ram_read_data_3;
    wire M_this_ppu_sprites_addr_9;
    wire \this_sprites_ram.mem_out_bus7_2 ;
    wire \this_sprites_ram.mem_out_bus3_2 ;
    wire M_this_substate_q_s_1;
    wire M_this_sprites_address_q_0_0_i_480_cascade_;
    wire M_this_sprites_address_qc_4_0;
    wire N_511_1;
    wire this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_4;
    wire this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_5;
    wire \this_vga_signals.N_659_cascade_ ;
    wire N_572_cascade_;
    wire M_this_sprites_address_qc_2_0;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_2 ;
    wire this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_3;
    wire M_this_sprites_address_q_0_0_i_484;
    wire M_this_sprites_address_qc_3_0_cascade_;
    wire N_1318_tz_0;
    wire \this_ppu.M_this_oam_ram_read_data_i_16 ;
    wire bfn_18_11_0_;
    wire \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ;
    wire \this_ppu.un2_vscroll_cry_0 ;
    wire \this_ppu.un2_vscroll_cry_1 ;
    wire \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ;
    wire M_this_oam_ram_read_data_i_17;
    wire \this_ppu.N_124 ;
    wire \this_ppu.N_124_cascade_ ;
    wire \this_ppu.un1_M_vaddress_q_2_c5_cascade_ ;
    wire \this_ppu.un1_M_vaddress_q_2_c5 ;
    wire \this_ppu.M_last_q ;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire M_this_vga_signals_line_clk_0;
    wire \this_sprites_ram.mem_out_bus4_0 ;
    wire \this_sprites_ram.mem_out_bus0_0 ;
    wire \this_ppu.vram_en_i_a2Z0Z_0 ;
    wire \this_ppu.vram_en_i_a2Z0Z_0_cascade_ ;
    wire M_this_ppu_vram_en_0_cascade_;
    wire \this_ppu.un1_M_haddress_q_3_c2_cascade_ ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2 ;
    wire M_this_ppu_vram_data_2;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_ ;
    wire M_this_ppu_vram_data_0;
    wire \this_sprites_ram.mem_out_bus5_2 ;
    wire \this_sprites_ram.mem_out_bus1_2 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ;
    wire dma_0_i;
    wire \this_sprites_ram.mem_out_bus4_3 ;
    wire \this_sprites_ram.mem_out_bus0_3 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0_cascade_ ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ;
    wire M_this_ppu_vram_data_3;
    wire \this_sprites_ram.mem_out_bus5_3 ;
    wire \this_sprites_ram.mem_out_bus1_3 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus7_3 ;
    wire \this_sprites_ram.mem_out_bus3_3 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ;
    wire \this_vga_signals.N_419_0_cascade_ ;
    wire N_440_0_cascade_;
    wire \this_vga_signals.N_467_0_cascade_ ;
    wire \this_vga_signals.N_467_0 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_6 ;
    wire N_510_0;
    wire M_this_sprites_address_qc_5_0;
    wire N_562_cascade_;
    wire M_this_sprites_address_q_0_0_i_476;
    wire M_this_sprites_address_q_0_0_i_496_cascade_;
    wire M_this_sprites_address_qc_0_1;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_0 ;
    wire N_773_cascade_;
    wire M_this_sprites_address_q_0_0_i_492;
    wire M_this_sprites_address_qc_1_0_cascade_;
    wire N_896_0;
    wire N_512_0;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_8 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1Z0Z_5 ;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_11_cascade_ ;
    wire this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_1;
    wire M_this_sprites_address_qc_10_0;
    wire N_1286_tz_0_cascade_;
    wire N_617;
    wire M_this_sprites_address_qc_11_0;
    wire bfn_19_5_0_;
    wire \this_ppu.un1_M_haddress_q_cry_0 ;
    wire \this_ppu.un1_M_haddress_q_cry_1 ;
    wire \this_ppu.un1_M_haddress_q_cry_2 ;
    wire \this_ppu.un1_M_haddress_q_cry_3 ;
    wire \this_ppu.un1_M_haddress_q_cry_4 ;
    wire \this_ppu.un1_M_haddress_q_cry_5 ;
    wire \this_ppu.un1_M_haddress_q_cry_6 ;
    wire \this_ppu.un1_M_haddress_q_cry_7 ;
    wire bfn_19_6_0_;
    wire \this_ppu.M_this_ppu_vram_addr_i_0 ;
    wire bfn_19_7_0_;
    wire \this_ppu.M_this_ppu_vram_addr_i_1 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_0 ;
    wire \this_ppu.M_this_ppu_vram_addr_i_2 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_1 ;
    wire \this_ppu.M_this_ppu_map_addr_i_0 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_2 ;
    wire \this_ppu.M_this_ppu_map_addr_i_1 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_3 ;
    wire \this_ppu.M_this_ppu_map_addr_i_2 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_4 ;
    wire \this_ppu.M_this_ppu_map_addr_i_3 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_5 ;
    wire \this_ppu.M_this_ppu_map_addr_i_4 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_6 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_7 ;
    wire bfn_19_8_0_;
    wire \this_ppu.M_state_qZ0Z_2 ;
    wire \this_ppu.M_state_qZ0Z_3 ;
    wire \this_ppu.N_122 ;
    wire \this_ppu.un1_M_vaddress_q_2_c2 ;
    wire this_vga_signals_vvisibility;
    wire \this_ppu.M_count_d_0_sqmuxa ;
    wire \this_ppu.M_last_q_RNIQRTEB ;
    wire M_this_ppu_map_addr_1;
    wire \this_ppu.un1_M_haddress_q_3_c2 ;
    wire M_this_ppu_map_addr_0;
    wire M_this_ppu_map_addr_4;
    wire \this_ppu.un1_M_haddress_q_3_c5 ;
    wire M_this_ppu_map_addr_2;
    wire M_this_ppu_map_addr_3;
    wire M_this_ppu_vram_en_0;
    wire \this_ppu.M_last_q_RNI3BB75 ;
    wire M_this_oam_ram_read_data_1;
    wire M_this_map_ram_read_data_1;
    wire M_this_ppu_sprites_addr_7;
    wire \this_sprites_ram.mem_out_bus4_1 ;
    wire \this_sprites_ram.mem_out_bus0_1 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_ ;
    wire \this_sprites_ram.mem_radregZ0Z_11 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ;
    wire M_this_ppu_vram_data_1;
    wire M_this_oam_ram_read_data_6;
    wire M_this_map_ram_read_data_6;
    wire \this_sprites_ram.mem_radregZ0Z_12 ;
    wire \this_sprites_ram.mem_out_bus6_1 ;
    wire \this_sprites_ram.mem_out_bus2_1 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus5_1 ;
    wire \this_sprites_ram.mem_out_bus1_1 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus7_1 ;
    wire \this_sprites_ram.mem_out_bus3_1 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_sprites_ram.mem_out_bus6_3 ;
    wire \this_sprites_ram.mem_out_bus2_3 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ;
    wire \this_vga_signals.N_746_cascade_ ;
    wire \this_vga_signals.N_505 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2Z0Z_0 ;
    wire \this_vga_signals.N_459_0 ;
    wire N_440_0;
    wire M_this_sprites_address_qZ0Z_0;
    wire un1_M_this_state_q_6_0;
    wire M_this_sprites_address_q_RNIRO0N6Z0Z_0;
    wire bfn_19_22_0_;
    wire M_this_sprites_address_qZ0Z_1;
    wire un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0;
    wire un1_M_this_sprites_address_q_cry_0;
    wire M_this_sprites_address_qZ0Z_2;
    wire un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0;
    wire un1_M_this_sprites_address_q_cry_1;
    wire M_this_sprites_address_qZ0Z_3;
    wire un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0;
    wire un1_M_this_sprites_address_q_cry_2;
    wire M_this_sprites_address_qZ0Z_4;
    wire un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0;
    wire un1_M_this_sprites_address_q_cry_3;
    wire M_this_sprites_address_qZ0Z_5;
    wire un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0;
    wire un1_M_this_sprites_address_q_cry_4;
    wire un1_M_this_sprites_address_q_cry_5;
    wire M_this_sprites_address_qZ0Z_7;
    wire un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0;
    wire un1_M_this_sprites_address_q_cry_6;
    wire un1_M_this_sprites_address_q_cry_7;
    wire M_this_sprites_address_qZ0Z_8;
    wire un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0;
    wire bfn_19_23_0_;
    wire un1_M_this_sprites_address_q_cry_8;
    wire un1_M_this_sprites_address_q_cry_9;
    wire un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0;
    wire un1_M_this_sprites_address_q_cry_10;
    wire un1_M_this_sprites_address_q_cry_11;
    wire un1_M_this_sprites_address_q_cry_12;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_9 ;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_13 ;
    wire un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0;
    wire N_627;
    wire N_509_0_cascade_;
    wire \this_vga_signals.N_415_0 ;
    wire un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0;
    wire M_this_sprites_address_q_0_0_i_472;
    wire this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_6;
    wire N_773;
    wire M_this_sprites_address_qZ0Z_6;
    wire M_this_sprites_address_qc_6_0;
    wire N_1282_tz_0;
    wire un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0;
    wire N_1290_tz_0_cascade_;
    wire N_607;
    wire M_this_sprites_address_qZ0Z_10;
    wire un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_10_cascade_ ;
    wire N_612;
    wire \this_ppu.un1_M_haddress_q_2_4 ;
    wire bfn_20_6_0_;
    wire \this_ppu.un1_M_vaddress_q_cry_0 ;
    wire \this_ppu.un1_M_vaddress_q_cry_1 ;
    wire \this_ppu.un1_M_vaddress_q_cry_2 ;
    wire \this_ppu.un1_M_vaddress_q_cry_3 ;
    wire \this_ppu.un1_M_vaddress_q_cry_4 ;
    wire \this_ppu.un1_M_vaddress_q_cry_5 ;
    wire \this_ppu.un1_M_vaddress_q_cry_6 ;
    wire \this_ppu.un1_M_vaddress_q_cry_7 ;
    wire \this_ppu.un1_M_haddress_q_2_cry_7_THRU_CO ;
    wire \this_ppu.un1_M_haddress_q_cry_7_THRU_CO ;
    wire bfn_20_7_0_;
    wire \this_ppu.vscroll8 ;
    wire M_this_oam_ram_read_data_i_11;
    wire \this_ppu.un2_vscroll_axb_0 ;
    wire M_this_ppu_sprites_addr_3;
    wire M_this_state_q_RNI0A0EZ0Z_6;
    wire M_this_state_q_RNI244K2Z0Z_6_cascade_;
    wire dma_0;
    wire M_this_state_q_fastZ0Z_9;
    wire N_861;
    wire N_861_cascade_;
    wire dma_c4_1;
    wire this_vga_signals_un20_i_a2_4_a3_0_a4_2_1;
    wire N_460_0_cascade_;
    wire N_560;
    wire M_this_map_ram_write_en_0;
    wire N_888_0_cascade_;
    wire \this_vga_signals.N_779 ;
    wire this_start_data_delay_M_last_q;
    wire port_enb_c;
    wire M_this_delay_clk_out_0;
    wire GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO;
    wire port_address_in_2;
    wire port_address_in_7;
    wire port_rw_in;
    wire \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5LZ0Z8_cascade_ ;
    wire M_this_substate_d_0_sqmuxa;
    wire M_this_substate_d_0_sqmuxa_cascade_;
    wire dma_c4_1_0;
    wire \this_vga_signals.N_732 ;
    wire un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0;
    wire N_622_cascade_;
    wire N_1278_tz_0;
    wire \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_12 ;
    wire M_this_sprites_address_qc_12_0;
    wire \this_vga_signals.N_427_0 ;
    wire M_this_state_qZ0Z_1;
    wire \this_vga_signals.N_427_0_cascade_ ;
    wire N_1274_tz_0;
    wire M_this_sprites_address_qc_0_2;
    wire \this_vga_signals.N_889_0 ;
    wire \this_vga_signals.N_889_0_cascade_ ;
    wire N_750;
    wire N_762;
    wire M_this_sprites_address_qZ0Z_9;
    wire N_750_cascade_;
    wire M_this_sprites_address_qc_9_0;
    wire port_address_in_0;
    wire \this_vga_signals.N_648 ;
    wire port_address_in_1;
    wire N_460_0;
    wire M_this_state_qZ0Z_8;
    wire M_this_state_qZ0Z_3;
    wire \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_2 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1 ;
    wire M_this_state_qZ0Z_2;
    wire N_250;
    wire \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3Z0Z_0_cascade_ ;
    wire \this_vga_signals.N_743 ;
    wire N_228;
    wire N_248;
    wire M_this_oam_ram_read_data_16;
    wire M_this_ppu_vram_addr_7;
    wire \this_ppu.M_this_ppu_vram_addr_i_7 ;
    wire bfn_21_6_0_;
    wire \this_ppu.M_vaddress_qZ0Z_1 ;
    wire M_this_oam_ram_read_data_17;
    wire \this_ppu.M_vaddress_q_i_1 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_0 ;
    wire \this_ppu.M_vaddress_qZ0Z_2 ;
    wire M_this_oam_ram_read_data_18;
    wire \this_ppu.M_vaddress_q_i_2 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_1 ;
    wire M_this_ppu_map_addr_5;
    wire \this_ppu.M_this_ppu_map_addr_i_5 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_2 ;
    wire M_this_ppu_map_addr_6;
    wire \this_ppu.M_this_ppu_map_addr_i_6 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_3 ;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.M_this_ppu_map_addr_i_7 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_4 ;
    wire M_this_ppu_map_addr_8;
    wire \this_ppu.M_this_ppu_map_addr_i_8 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_5 ;
    wire M_this_ppu_map_addr_9;
    wire \this_ppu.M_this_ppu_map_addr_i_9 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_6 ;
    wire \this_ppu.un1_M_vaddress_q_3_cry_7 ;
    wire bfn_21_7_0_;
    wire \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ;
    wire M_this_oam_ram_write_data_16;
    wire M_this_oam_ram_read_data_i_19;
    wire M_this_data_tmp_qZ0Z_16;
    wire this_vga_signals_un20_i_a2_0_a3_0_a4_2_2;
    wire \this_sprites_ram.mem_out_bus5_0 ;
    wire \this_sprites_ram.mem_out_bus1_0 ;
    wire \this_sprites_ram.mem_radregZ0Z_13 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ;
    wire M_this_state_qZ0Z_10;
    wire \this_vga_signals.N_433_0_cascade_ ;
    wire \this_vga_signals.N_442_0_cascade_ ;
    wire \this_vga_signals.N_719_cascade_ ;
    wire this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2;
    wire this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2_cascade_;
    wire N_307_0_cascade_;
    wire M_this_state_qZ0Z_5;
    wire \this_vga_signals.N_665_1_cascade_ ;
    wire M_this_data_count_q_3_0_13_cascade_;
    wire N_755;
    wire bfn_21_22_0_;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_q_s_2;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire M_this_data_count_q_s_8;
    wire bfn_21_23_0_;
    wire M_this_data_count_q_s_9;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_q_cry_9_THRU_CO;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_q_s_11;
    wire M_this_data_count_q_cry_10;
    wire M_this_data_count_q_s_12;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_q_cry_12_THRU_CO;
    wire M_this_data_count_q_cry_12;
    wire CONSTANT_ONE_NET;
    wire M_this_data_count_q_s_14;
    wire M_this_data_count_q_cry_13;
    wire M_this_data_count_q_cry_14;
    wire M_this_data_count_q_s_15;
    wire \this_vga_signals.N_431_0 ;
    wire \this_vga_signals.N_428_0 ;
    wire N_226;
    wire M_this_data_tmp_qZ0Z_6;
    wire M_this_oam_ram_write_data_6;
    wire M_this_data_tmp_qZ0Z_2;
    wire M_this_oam_ram_write_data_2;
    wire M_this_data_tmp_qZ0Z_1;
    wire M_this_oam_ram_write_data_1;
    wire \this_ppu.un1_oam_data_c2_cascade_ ;
    wire \this_ppu.un1_M_vaddress_q_3_6 ;
    wire M_this_data_tmp_qZ0Z_23;
    wire M_this_oam_ram_write_data_23;
    wire M_this_oam_ram_read_data_22;
    wire M_this_oam_ram_read_data_23;
    wire \this_ppu.un1_oam_data_c2 ;
    wire \this_ppu.un1_M_vaddress_q_3_7 ;
    wire M_this_oam_ram_write_data_25;
    wire M_this_data_tmp_qZ0Z_17;
    wire M_this_oam_ram_write_data_17;
    wire \this_ppu.un1_M_vaddress_q_3_4 ;
    wire M_this_oam_ram_write_data_24;
    wire M_this_state_qZ0Z_12;
    wire M_this_state_qZ0Z_11;
    wire \this_vga_signals.N_469_0_cascade_ ;
    wire \this_vga_signals.N_506_cascade_ ;
    wire M_this_state_qZ0Z_6;
    wire M_this_data_count_qZ0Z_14;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_qZ0Z_15;
    wire M_this_data_count_qZ0Z_12;
    wire \this_vga_signals.N_745 ;
    wire \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2 ;
    wire \this_vga_signals.N_442_0 ;
    wire M_this_reset_cond_out_0;
    wire \this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2_cascade_ ;
    wire \this_vga_signals.M_this_data_count_qlde_iZ0Z_1 ;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_qZ0Z_0;
    wire M_this_state_d62_11;
    wire M_this_state_d62_8_cascade_;
    wire un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2;
    wire M_this_state_d62_cascade_;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_qZ0Z_9;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_state_d62_10;
    wire M_this_state_d62_9;
    wire M_this_data_count_q_cry_0_THRU_CO;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_q_cry_2_THRU_CO;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_q_cry_3_THRU_CO;
    wire M_this_data_count_qZ0Z_4;
    wire M_this_data_count_q_cry_4_THRU_CO;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_q_cry_5_THRU_CO;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_oam_ram_write_data_4;
    wire M_this_data_tmp_qZ0Z_7;
    wire M_this_oam_ram_write_data_7;
    wire M_this_oam_ram_write_data_8;
    wire M_this_oam_ram_write_data_0;
    wire M_this_data_tmp_qZ0Z_4;
    wire M_this_data_tmp_qZ0Z_0;
    wire N_1412_0;
    wire M_this_data_tmp_qZ0Z_3;
    wire M_this_oam_ram_write_data_3;
    wire M_this_oam_ram_write_data_10;
    wire M_this_data_tmp_qZ0Z_10;
    wire M_this_oam_ram_write_data_11;
    wire M_this_oam_address_qZ0Z_5;
    wire M_this_oam_address_qZ0Z_4;
    wire M_this_data_tmp_qZ0Z_11;
    wire M_this_data_tmp_qZ0Z_8;
    wire N_413_0;
    wire un1_M_this_oam_address_q_c4;
    wire M_this_oam_address_qZ0Z_3;
    wire M_this_oam_address_qZ0Z_2;
    wire M_this_oam_address_qZ0Z_0;
    wire M_this_state_qZ0Z_13;
    wire M_this_oam_address_qZ0Z_1;
    wire un1_M_this_oam_address_q_c2;
    wire \this_vga_signals.N_461_0 ;
    wire \this_vga_signals.N_747 ;
    wire M_this_state_qZ0Z_9;
    wire M_this_state_qZ0Z_7;
    wire \this_vga_signals.N_433_0 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_i_1Z0Z_0 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4Z0Z_0 ;
    wire M_this_state_d62;
    wire \this_vga_signals.N_746 ;
    wire \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12 ;
    wire M_this_oam_address_q_0_i_o3_0_a2_5;
    wire \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12_cascade_ ;
    wire led_c_1;
    wire M_this_substate_qZ0;
    wire \this_vga_signals.N_419_0 ;
    wire M_this_data_count_q_cry_6_THRU_CO;
    wire N_716_i;
    wire M_this_data_count_qZ0Z_7;
    wire N_364;
    wire port_data_c_0;
    wire M_this_state_qZ0Z_4;
    wire N_888_0;
    wire N_760_cascade_;
    wire M_this_external_address_q_3_0_12;
    wire \this_sprites_ram.mem_WE_4 ;
    wire \this_ppu.un1_M_haddress_q_2_5 ;
    wire M_this_oam_ram_write_data_13;
    wire M_this_oam_ram_write_data_15;
    wire M_this_oam_ram_read_data_15;
    wire \this_ppu.un1_M_haddress_q_2_7 ;
    wire M_this_oam_ram_read_data_12;
    wire M_this_oam_ram_read_data_11;
    wire \this_ppu.un1_oam_data_1_c2 ;
    wire M_this_oam_ram_read_data_14;
    wire \this_ppu.un1_oam_data_1_c2_cascade_ ;
    wire M_this_oam_ram_read_data_13;
    wire \this_ppu.un1_M_haddress_q_2_6 ;
    wire M_this_data_tmp_qZ0Z_12;
    wire M_this_oam_ram_write_data_12;
    wire M_this_oam_ram_read_data_21;
    wire M_this_oam_ram_read_data_20;
    wire M_this_oam_ram_read_data_19;
    wire \this_ppu.un1_M_vaddress_q_3_5 ;
    wire M_this_data_tmp_qZ0Z_5;
    wire M_this_oam_ram_write_data_5;
    wire M_this_oam_ram_read_data_9;
    wire M_this_oam_ram_write_data_9;
    wire M_this_oam_ram_write_data_18;
    wire M_this_oam_ram_write_data_20;
    wire M_this_oam_ram_write_data_29;
    wire M_this_oam_ram_write_data_30;
    wire M_this_data_tmp_qZ0Z_22;
    wire M_this_oam_ram_write_data_22;
    wire M_this_oam_ram_write_data_31;
    wire M_this_data_tmp_qZ0Z_18;
    wire M_this_data_tmp_qZ0Z_20;
    wire port_data_c_4;
    wire M_this_oam_ram_write_data_28;
    wire M_this_data_tmp_qZ0Z_21;
    wire M_this_oam_ram_write_data_21;
    wire M_this_oam_address_qZ0Z_6;
    wire un1_M_this_oam_address_q_c6;
    wire M_this_oam_address_qZ0Z_7;
    wire N_404_g;
    wire M_this_data_tmp_qZ0Z_9;
    wire \this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ;
    wire bfn_24_11_0_;
    wire M_this_oam_ram_read_data_i_9;
    wire \this_ppu.un2_hscroll_cry_0 ;
    wire M_this_oam_ram_read_data_10;
    wire \this_ppu.un2_hscroll_cry_1 ;
    wire M_this_oam_ram_write_data_26;
    wire M_this_oam_ram_write_data_19;
    wire M_this_ppu_vram_addr_1;
    wire \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ;
    wire M_this_ppu_sprites_addr_1;
    wire M_this_oam_ram_read_data_8;
    wire M_this_ppu_vram_addr_2;
    wire \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ;
    wire M_this_ppu_sprites_addr_2;
    wire \this_ppu.un2_hscroll_axb_0 ;
    wire M_this_ppu_vram_addr_0;
    wire M_this_ppu_sprites_addr_0;
    wire M_this_data_tmp_qZ0Z_19;
    wire N_1396_0;
    wire M_this_oam_ram_read_data_0;
    wire M_this_map_ram_read_data_0;
    wire \this_ppu.M_state_qZ0Z_4 ;
    wire \this_ppu.M_state_qZ0Z_5 ;
    wire M_this_ppu_sprites_addr_6;
    wire \this_sprites_ram.mem_WE_14 ;
    wire \this_sprites_ram.mem_WE_12 ;
    wire \this_sprites_ram.mem_WE_0 ;
    wire port_data_c_1;
    wire this_vga_signals_M_this_external_address_q_3_i_0_0_15;
    wire N_661;
    wire \this_sprites_ram.mem_WE_2 ;
    wire \this_vga_signals.N_665_1 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3LZ0Z4 ;
    wire \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4LZ0Z6 ;
    wire port_address_in_3;
    wire port_address_in_5;
    wire port_address_in_6;
    wire port_address_in_4;
    wire \this_vga_signals.un1_M_this_state_q_19_i_0_o2Z0Z_4 ;
    wire port_data_c_2;
    wire N_760;
    wire M_this_sprites_address_qZ0Z_12;
    wire N_25_0;
    wire M_this_sprites_address_qZ0Z_13;
    wire M_this_sprites_address_qZ0Z_11;
    wire \this_sprites_ram.mem_WE_6 ;
    wire M_this_oam_ram_write_data_14;
    wire port_data_c_7;
    wire M_this_data_tmp_qZ0Z_15;
    wire port_data_c_6;
    wire M_this_data_tmp_qZ0Z_14;
    wire port_data_c_5;
    wire M_this_data_tmp_qZ0Z_13;
    wire N_1404_0;
    wire M_this_reset_cond_out_g_0;
    wire port_data_c_3;
    wire M_this_oam_ram_write_data_0_sqmuxa;
    wire M_this_oam_ram_write_data_27;
    wire M_this_external_address_q_3_0_13;
    wire N_312_0;
    wire M_this_external_address_qZ0Z_0;
    wire bfn_26_21_0_;
    wire M_this_external_address_qZ0Z_1;
    wire M_this_external_address_q_cry_0;
    wire M_this_external_address_qZ0Z_2;
    wire M_this_external_address_q_cry_1;
    wire M_this_external_address_qZ0Z_3;
    wire M_this_external_address_q_cry_2;
    wire M_this_external_address_qZ0Z_4;
    wire M_this_external_address_q_cry_3;
    wire M_this_external_address_qZ0Z_5;
    wire M_this_external_address_q_cry_4;
    wire M_this_external_address_qZ0Z_6;
    wire M_this_external_address_q_cry_5;
    wire N_49;
    wire M_this_external_address_qZ0Z_7;
    wire M_this_external_address_q_cry_6;
    wire M_this_external_address_q_cry_7;
    wire clk_0_c_g;
    wire N_47;
    wire M_this_external_address_qZ0Z_8;
    wire M_this_external_address_q_s_8;
    wire bfn_26_22_0_;
    wire M_this_external_address_qZ0Z_9;
    wire M_this_external_address_q_s_9;
    wire M_this_external_address_q_cry_8;
    wire M_this_external_address_qZ0Z_10;
    wire M_this_external_address_q_s_10;
    wire M_this_external_address_q_cry_9;
    wire M_this_external_address_qZ0Z_11;
    wire M_this_external_address_q_s_11;
    wire M_this_external_address_q_cry_10;
    wire M_this_external_address_qZ0Z_12;
    wire M_this_external_address_q_cry_11_THRU_CO;
    wire M_this_external_address_q_cry_11;
    wire M_this_external_address_qZ0Z_13;
    wire M_this_external_address_q_cry_12_THRU_CO;
    wire M_this_external_address_q_cry_12;
    wire M_this_external_address_qZ0Z_14;
    wire M_this_external_address_q_cry_13_THRU_CO;
    wire M_this_external_address_q_cry_13;
    wire M_this_external_address_qZ0Z_15;
    wire M_this_external_address_q_cry_14;
    wire M_this_external_address_q_s_15;
    wire _gnd_net_;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_map_ram_read_data_3,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_map_ram_read_data_2,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_map_ram_read_data_1,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_map_ram_read_data_0,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__27978,N__27276,N__27342,N__27417,N__27486,N__21303,N__21174,N__21246,N__21447,N__21374}),
            .WADDR({dangling_wire_13,N__11781,N__11814,N__11844,N__11874,N__11904,N__11934,N__11964,N__11610,N__11640,N__11667}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__18555,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__15723,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__12507,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__13314,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__36969),
            .RE(N__28934),
            .WCLKE(N__25299),
            .WCLK(N__36970),
            .WE(N__28851));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__27972,N__27269,N__27336,N__27411,N__27480,N__21297,N__21167,N__21236,N__21437,N__21362}),
            .WADDR({dangling_wire_55,N__11775,N__11808,N__11838,N__11868,N__11898,N__11928,N__11958,N__11604,N__11634,N__11661}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__13305,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__13968,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__12495,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__11709,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__36973),
            .RE(N__28935),
            .WCLKE(N__25292),
            .WCLK(N__36974),
            .WE(N__28852));
    defparam \this_oam_ram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_0_physical  (
            .RDATA({M_this_oam_ram_read_data_15,M_this_oam_ram_read_data_14,M_this_oam_ram_read_data_13,M_this_oam_ram_read_data_12,M_this_oam_ram_read_data_11,M_this_oam_ram_read_data_10,M_this_oam_ram_read_data_9,M_this_oam_ram_read_data_8,M_this_oam_ram_read_data_7,M_this_oam_ram_read_data_6,M_this_oam_ram_read_data_5,M_this_oam_ram_read_data_4,M_this_oam_ram_read_data_3,M_this_oam_ram_read_data_2,M_this_oam_ram_read_data_1,M_this_oam_ram_read_data_0}),
            .RADDR({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .WADDR({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,N__32241,N__32274,N__30120,N__30084,N__30747,N__30708}),
            .MASK({dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115}),
            .WDATA({N__31881,N__34590,N__31887,N__32148,N__30132,N__30150,N__31968,N__29859,N__29871,N__28395,N__32007,N__29898,N__30162,N__28371,N__28353,N__29850}),
            .RCLKE(),
            .RCLK(N__36859),
            .RE(N__29117),
            .WCLKE(N__35709),
            .WCLK(N__36860),
            .WE(N__29102));
    defparam \this_oam_ram.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,M_this_oam_ram_read_data_23,M_this_oam_ram_read_data_22,M_this_oam_ram_read_data_21,M_this_oam_ram_read_data_20,M_this_oam_ram_read_data_19,M_this_oam_ram_read_data_18,M_this_oam_ram_read_data_17,M_this_oam_ram_read_data_16}),
            .RADDR({dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134}),
            .WADDR({dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,N__32234,N__32268,N__30114,N__30078,N__30741,N__30702}),
            .MASK({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155}),
            .WDATA({N__32466,N__31944,N__31950,N__32298,N__35511,N__33090,N__29172,N__29430,N__29253,N__32475,N__32280,N__31956,N__33078,N__31962,N__29154,N__27894}),
            .RCLKE(),
            .RCLK(N__36874),
            .RE(N__29081),
            .WCLKE(N__35708),
            .WCLK(N__36875),
            .WE(N__29098));
    defparam \this_sprites_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,\this_sprites_ram.mem_out_bus0_1 ,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,\this_sprites_ram.mem_out_bus0_0 ,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .RADDR({N__13111,N__19232,N__18480,N__20987,N__33601,N__18279,N__18100,N__24773,N__32621,N__32878,N__34135}),
            .WADDR({N__24615,N__26076,N__23688,N__23937,N__24232,N__22110,N__22358,N__22608,N__22857,N__23087,N__23351}),
            .MASK({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185}),
            .WDATA({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,N__26754,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,N__28493,dangling_wire_197,dangling_wire_198,dangling_wire_199}),
            .RCLKE(),
            .RCLK(N__36891),
            .RE(N__29068),
            .WCLKE(N__33483),
            .WCLK(N__36890),
            .WE(N__29025));
    defparam \this_sprites_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,\this_sprites_ram.mem_out_bus0_3 ,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,\this_sprites_ram.mem_out_bus0_2 ,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .RADDR({N__13125,N__19233,N__18459,N__20997,N__33600,N__18194,N__18101,N__24802,N__32566,N__32842,N__34085}),
            .WADDR({N__24605,N__26072,N__23683,N__23961,N__24233,N__22106,N__22367,N__22604,N__22800,N__23110,N__23330}),
            .MASK({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229}),
            .WDATA({dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,N__26883,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,N__26653,dangling_wire_241,dangling_wire_242,dangling_wire_243}),
            .RCLKE(),
            .RCLK(N__36901),
            .RE(N__29023),
            .WCLKE(N__33482),
            .WCLK(N__36902),
            .WE(N__29024));
    defparam \this_sprites_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,\this_sprites_ram.mem_out_bus1_1 ,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,\this_sprites_ram.mem_out_bus1_0 ,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .RADDR({N__13107,N__19182,N__18460,N__20961,N__33550,N__18274,N__18024,N__24772,N__32534,N__32843,N__34062}),
            .WADDR({N__24589,N__26065,N__23682,N__23893,N__24205,N__22099,N__22368,N__22603,N__22858,N__23109,N__23329}),
            .MASK({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273}),
            .WDATA({dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,N__26753,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,N__28485,dangling_wire_285,dangling_wire_286,dangling_wire_287}),
            .RCLKE(),
            .RCLK(N__36917),
            .RE(N__29011),
            .WCLKE(N__33458),
            .WCLK(N__36918),
            .WE(N__28939));
    defparam \this_sprites_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,\this_sprites_ram.mem_out_bus1_3 ,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,\this_sprites_ram.mem_out_bus1_2 ,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .RADDR({N__13105,N__19228,N__18491,N__20992,N__33524,N__18275,N__18099,N__24768,N__32567,N__32882,N__34111}),
            .WADDR({N__24588,N__26055,N__23667,N__23970,N__24206,N__22088,N__22345,N__22592,N__22859,N__23094,N__23328}),
            .MASK({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317}),
            .WDATA({dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,N__26879,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,N__26662,dangling_wire_329,dangling_wire_330,dangling_wire_331}),
            .RCLKE(),
            .RCLK(N__36929),
            .RE(N__28937),
            .WCLKE(N__33459),
            .WCLK(N__36930),
            .WE(N__28938));
    defparam \this_sprites_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,\this_sprites_ram.mem_out_bus2_1 ,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,\this_sprites_ram.mem_out_bus2_0 ,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .RADDR({N__13081,N__19146,N__18481,N__20993,N__33646,N__18316,N__18102,N__24809,N__32648,N__32971,N__34203}),
            .WADDR({N__24627,N__26019,N__23687,N__23963,N__24240,N__22046,N__22357,N__22557,N__22856,N__23111,N__23355}),
            .MASK({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361}),
            .WDATA({dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,N__26744,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,N__28494,dangling_wire_373,dangling_wire_374,dangling_wire_375}),
            .RCLKE(),
            .RCLK(N__36945),
            .RE(N__28717),
            .WCLKE(N__17450),
            .WCLK(N__36946),
            .WE(N__28778));
    defparam \this_sprites_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,\this_sprites_ram.mem_out_bus2_3 ,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,\this_sprites_ram.mem_out_bus2_2 ,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .RADDR({N__13036,N__19230,N__18505,N__20995,N__33658,N__18328,N__18113,N__24810,N__32649,N__32983,N__34213}),
            .WADDR({N__24623,N__26018,N__23677,N__23942,N__24237,N__22041,N__22352,N__22556,N__22855,N__23011,N__23317}),
            .MASK({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405}),
            .WDATA({dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,N__26854,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,N__26664,dangling_wire_417,dangling_wire_418,dangling_wire_419}),
            .RCLKE(),
            .RCLK(N__36952),
            .RE(N__28736),
            .WCLKE(N__17451),
            .WCLK(N__36953),
            .WE(N__28779));
    defparam \this_sprites_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,\this_sprites_ram.mem_out_bus3_1 ,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,\this_sprites_ram.mem_out_bus3_0 ,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .RADDR({N__13082,N__19231,N__18506,N__20988,N__33665,N__18329,N__18114,N__24811,N__32650,N__32984,N__34214}),
            .WADDR({N__24616,N__25980,N__23654,N__23906,N__24238,N__22042,N__22356,N__22554,N__22853,N__23101,N__23353}),
            .MASK({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449}),
            .WDATA({dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,N__26745,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,N__28489,dangling_wire_461,dangling_wire_462,dangling_wire_463}),
            .RCLKE(),
            .RCLK(N__36959),
            .RE(N__28737),
            .WCLKE(N__15753),
            .WCLK(N__36960),
            .WE(N__28842));
    defparam \this_sprites_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,\this_sprites_ram.mem_out_bus3_3 ,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,\this_sprites_ram.mem_out_bus3_2 ,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .RADDR({N__13112,N__19183,N__18510,N__20994,N__33666,N__18333,N__18112,N__24812,N__32651,N__32988,N__34215}),
            .WADDR({N__24593,N__26017,N__23681,N__23946,N__24236,N__22070,N__22366,N__22555,N__22854,N__23112,N__23354}),
            .MASK({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493}),
            .WDATA({dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,N__26855,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,N__26663,dangling_wire_505,dangling_wire_506,dangling_wire_507}),
            .RCLKE(),
            .RCLK(N__36964),
            .RE(N__28850),
            .WCLKE(N__15752),
            .WCLK(N__36965),
            .WE(N__28843));
    defparam \this_sprites_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,\this_sprites_ram.mem_out_bus4_1 ,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,\this_sprites_ram.mem_out_bus4_0 ,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .RADDR({N__13127,N__19214,N__18494,N__20957,N__33656,N__18326,N__18117,N__24808,N__32660,N__32981,N__34175}),
            .WADDR({N__24582,N__26042,N__23665,N__23968,N__24222,N__22084,N__22279,N__22587,N__22863,N__23089,N__23335}),
            .MASK({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537}),
            .WDATA({dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,N__26748,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,N__28460,dangling_wire_549,dangling_wire_550,dangling_wire_551}),
            .RCLKE(),
            .RCLK(N__36975),
            .RE(N__29121),
            .WCLKE(N__34607),
            .WCLK(N__36976),
            .WE(N__29122));
    defparam \this_sprites_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,\this_sprites_ram.mem_out_bus4_3 ,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,\this_sprites_ram.mem_out_bus4_2 ,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .RADDR({N__13131,N__19193,N__18495,N__20956,N__33657,N__18327,N__18116,N__24813,N__32661,N__32982,N__34190}),
            .WADDR({N__24583,N__26041,N__23653,N__23969,N__24223,N__22098,N__22348,N__22602,N__22817,N__23108,N__23336}),
            .MASK({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581}),
            .WDATA({dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,N__26877,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,N__26660,dangling_wire_593,dangling_wire_594,dangling_wire_595}),
            .RCLKE(),
            .RCLK(N__36977),
            .RE(N__28936),
            .WCLKE(N__34608),
            .WCLK(N__36978),
            .WE(N__29123));
    defparam \this_sprites_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,\this_sprites_ram.mem_out_bus5_1 ,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,\this_sprites_ram.mem_out_bus5_0 ,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .RADDR({N__13106,N__19213,N__18493,N__20916,N__33639,N__18312,N__18106,N__24804,N__32653,N__32964,N__34174}),
            .WADDR({N__24581,N__26020,N__23664,N__23954,N__24224,N__22083,N__22365,N__22586,N__22869,N__23088,N__23334}),
            .MASK({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625}),
            .WDATA({dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,N__26749,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,N__28445,dangling_wire_637,dangling_wire_638,dangling_wire_639}),
            .RCLKE(),
            .RCLK(N__36971),
            .RE(N__28853),
            .WCLKE(N__31929),
            .WCLK(N__36972),
            .WE(N__29107));
    defparam \this_sprites_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,\this_sprites_ram.mem_out_bus5_3 ,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,\this_sprites_ram.mem_out_bus5_2 ,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .RADDR({N__13118,N__19181,N__18492,N__20980,N__33638,N__18308,N__18110,N__24780,N__32652,N__32963,N__34157}),
            .WADDR({N__24580,N__26024,N__23629,N__23883,N__24225,N__22060,N__22335,N__22559,N__22864,N__23055,N__23352}),
            .MASK({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669}),
            .WDATA({dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,N__26856,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,N__26651,dangling_wire_681,dangling_wire_682,dangling_wire_683}),
            .RCLKE(),
            .RCLK(N__36967),
            .RE(N__29061),
            .WCLKE(N__31925),
            .WCLK(N__36968),
            .WE(N__29106));
    defparam \this_sprites_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,\this_sprites_ram.mem_out_bus6_1 ,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,\this_sprites_ram.mem_out_bus6_0 ,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .RADDR({N__13117,N__19215,N__18467,N__20976,N__33613,N__18288,N__18111,N__24803,N__32635,N__32938,N__34156}),
            .WADDR({N__24584,N__25990,N__23628,N__23947,N__24149,N__22059,N__22334,N__22558,N__22801,N__23054,N__23337}),
            .MASK({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713}),
            .WDATA({dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,N__26747,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,dangling_wire_723,dangling_wire_724,N__28444,dangling_wire_725,dangling_wire_726,dangling_wire_727}),
            .RCLKE(),
            .RCLK(N__36961),
            .RE(N__29082),
            .WCLKE(N__33174),
            .WCLK(N__36962),
            .WE(N__29083));
    defparam \this_sprites_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,\this_sprites_ram.mem_out_bus6_3 ,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,\this_sprites_ram.mem_out_bus6_2 ,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .RADDR({N__13086,N__19212,N__18466,N__20996,N__33612,N__18281,N__18115,N__24776,N__32634,N__32937,N__34137}),
            .WADDR({N__24585,N__26028,N__23636,N__23938,N__24239,N__22014,N__22347,N__22569,N__22845,N__22974,N__23307}),
            .MASK({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,dangling_wire_753,dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757}),
            .WDATA({dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,N__26853,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,dangling_wire_767,dangling_wire_768,N__26652,dangling_wire_769,dangling_wire_770,dangling_wire_771}),
            .RCLKE(),
            .RCLK(N__36955),
            .RE(N__29066),
            .WCLKE(N__33170),
            .WCLK(N__36956),
            .WE(N__29067));
    defparam \this_sprites_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,\this_sprites_ram.mem_out_bus7_1 ,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,\this_sprites_ram.mem_out_bus7_0 ,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .RADDR({N__13113,N__19165,N__18465,N__20972,N__33582,N__18280,N__18094,N__24775,N__32603,N__32909,N__34136}),
            .WADDR({N__24586,N__26029,N__23637,N__23964,N__24235,N__22047,N__22346,N__22570,N__22852,N__23065,N__23341}),
            .MASK({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801}),
            .WDATA({dangling_wire_802,dangling_wire_803,dangling_wire_804,dangling_wire_805,N__26746,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,dangling_wire_811,dangling_wire_812,N__28461,dangling_wire_813,dangling_wire_814,dangling_wire_815}),
            .RCLKE(),
            .RCLK(N__36949),
            .RE(N__29042),
            .WCLKE(N__33432),
            .WCLK(N__36950),
            .WE(N__29016));
    defparam \this_sprites_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,\this_sprites_ram.mem_out_bus7_3 ,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,\this_sprites_ram.mem_out_bus7_2 ,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .RADDR({N__13126,N__19229,N__18464,N__20962,N__33581,N__18307,N__18098,N__24774,N__32602,N__32908,N__34112}),
            .WADDR({N__24587,N__26043,N__23666,N__23962,N__24234,N__22071,N__22309,N__22591,N__22868,N__23093,N__23327}),
            .MASK({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,dangling_wire_841,dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845}),
            .WDATA({dangling_wire_846,dangling_wire_847,dangling_wire_848,dangling_wire_849,N__26878,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,dangling_wire_855,dangling_wire_856,N__26661,dangling_wire_857,dangling_wire_858,dangling_wire_859}),
            .RCLKE(),
            .RCLK(N__36939),
            .RE(N__29065),
            .WCLKE(N__33428),
            .WCLK(N__36940),
            .WE(N__29015));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_872,dangling_wire_873,dangling_wire_874,N__12696,N__11700,N__12570,N__12540,N__12555,N__13236,N__12807,N__12786}),
            .WADDR({dangling_wire_875,dangling_wire_876,dangling_wire_877,N__27824,N__21170,N__21245,N__21446,N__21375,N__32754,N__33065,N__34314}),
            .MASK({dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,dangling_wire_892,dangling_wire_893}),
            .WDATA({dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,dangling_wire_899,dangling_wire_900,dangling_wire_901,dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,N__20013,N__19803,N__21720,N__19758}),
            .RCLKE(),
            .RCLK(N__36934),
            .RE(N__28652),
            .WCLKE(N__21102),
            .WCLK(N__36935),
            .WE(N__28660));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__37831),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__37833),
            .DIN(N__37832),
            .DOUT(N__37831),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__37833),
            .PADOUT(N__37832),
            .PADIN(N__37831),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__37822),
            .DIN(N__37821),
            .DOUT(N__37820),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__37822),
            .PADOUT(N__37821),
            .PADIN(N__37820),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__37813),
            .DIN(N__37812),
            .DOUT(N__37811),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__37813),
            .PADOUT(N__37812),
            .PADIN(N__37811),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__37804),
            .DIN(N__37803),
            .DOUT(N__37802),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__37804),
            .PADOUT(N__37803),
            .PADIN(N__37802),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12114),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__37795),
            .DIN(N__37794),
            .DOUT(N__37793),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__37795),
            .PADOUT(N__37794),
            .PADIN(N__37793),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13743),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__37786),
            .DIN(N__37785),
            .DOUT(N__37784),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__37786),
            .PADOUT(N__37785),
            .PADIN(N__37784),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29124),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__37777),
            .DIN(N__37776),
            .DOUT(N__37775),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__37777),
            .PADOUT(N__37776),
            .PADIN(N__37775),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__31653),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__37768),
            .DIN(N__37767),
            .DOUT(N__37766),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__37768),
            .PADOUT(N__37767),
            .PADIN(N__37766),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__37759),
            .DIN(N__37758),
            .DOUT(N__37757),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__37759),
            .PADOUT(N__37758),
            .PADIN(N__37757),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__37750),
            .DIN(N__37749),
            .DOUT(N__37748),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__37750),
            .PADOUT(N__37749),
            .PADIN(N__37748),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__37741),
            .DIN(N__37740),
            .DOUT(N__37739),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__37741),
            .PADOUT(N__37740),
            .PADIN(N__37739),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__37732),
            .DIN(N__37731),
            .DOUT(N__37730),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__37732),
            .PADOUT(N__37731),
            .PADIN(N__37730),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__37723),
            .DIN(N__37722),
            .DOUT(N__37721),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__37723),
            .PADOUT(N__37722),
            .PADIN(N__37721),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__37714),
            .DIN(N__37713),
            .DOUT(N__37712),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__37714),
            .PADOUT(N__37713),
            .PADIN(N__37712),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__35484),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20157));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__37705),
            .DIN(N__37704),
            .DOUT(N__37703),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__37705),
            .PADOUT(N__37704),
            .PADIN(N__37703),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__35457),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20211));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__37696),
            .DIN(N__37695),
            .DOUT(N__37694),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__37696),
            .PADOUT(N__37695),
            .PADIN(N__37694),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__35436),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20187));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__37687),
            .DIN(N__37686),
            .DOUT(N__37685),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__37687),
            .PADOUT(N__37686),
            .PADIN(N__37685),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__35409),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20155));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__37678),
            .DIN(N__37677),
            .DOUT(N__37676),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__37678),
            .PADOUT(N__37677),
            .PADIN(N__37676),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__35382),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20214));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__37669),
            .DIN(N__37668),
            .DOUT(N__37667),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__37669),
            .PADOUT(N__37668),
            .PADIN(N__37667),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__37158),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20212));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__37660),
            .DIN(N__37659),
            .DOUT(N__37658),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__37660),
            .PADOUT(N__37659),
            .PADIN(N__37658),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__37140),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20192));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__37651),
            .DIN(N__37650),
            .DOUT(N__37649),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__37651),
            .PADOUT(N__37650),
            .PADIN(N__37649),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__37008),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20229));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__37642),
            .DIN(N__37641),
            .DOUT(N__37640),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__37642),
            .PADOUT(N__37641),
            .PADIN(N__37640),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36438),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20159));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__37633),
            .DIN(N__37632),
            .DOUT(N__37631),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__37633),
            .PADOUT(N__37632),
            .PADIN(N__37631),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36399),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20156));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__37624),
            .DIN(N__37623),
            .DOUT(N__37622),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__37624),
            .PADOUT(N__37623),
            .PADIN(N__37622),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37353),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20215));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__37615),
            .DIN(N__37614),
            .DOUT(N__37613),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__37615),
            .PADOUT(N__37614),
            .PADIN(N__37613),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37305),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20213));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__37606),
            .DIN(N__37605),
            .DOUT(N__37604),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__37606),
            .PADOUT(N__37605),
            .PADIN(N__37604),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37260),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20151));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__37597),
            .DIN(N__37596),
            .DOUT(N__37595),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__37597),
            .PADOUT(N__37596),
            .PADIN(N__37595),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37215),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20228));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__37588),
            .DIN(N__37587),
            .DOUT(N__37586),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__37588),
            .PADOUT(N__37587),
            .PADIN(N__37586),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36525),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20158));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__37579),
            .DIN(N__37578),
            .DOUT(N__37577),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__37579),
            .PADOUT(N__37578),
            .PADIN(N__37577),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36483),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20188));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__37570),
            .DIN(N__37569),
            .DOUT(N__37568),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__37570),
            .PADOUT(N__37569),
            .PADIN(N__37568),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__37561),
            .DIN(N__37560),
            .DOUT(N__37559),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__37561),
            .PADOUT(N__37560),
            .PADIN(N__37559),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__37552),
            .DIN(N__37551),
            .DOUT(N__37550),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__37552),
            .PADOUT(N__37551),
            .PADIN(N__37550),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__37543),
            .DIN(N__37542),
            .DOUT(N__37541),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__37543),
            .PADOUT(N__37542),
            .PADIN(N__37541),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__37534),
            .DIN(N__37533),
            .DOUT(N__37532),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__37534),
            .PADOUT(N__37533),
            .PADIN(N__37532),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__37525),
            .DIN(N__37524),
            .DOUT(N__37523),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__37525),
            .PADOUT(N__37524),
            .PADIN(N__37523),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__37516),
            .DIN(N__37515),
            .DOUT(N__37514),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__37516),
            .PADOUT(N__37515),
            .PADIN(N__37514),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__37507),
            .DIN(N__37506),
            .DOUT(N__37505),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__37507),
            .PADOUT(N__37506),
            .PADIN(N__37505),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__37498),
            .DIN(N__37497),
            .DOUT(N__37496),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__37498),
            .PADOUT(N__37497),
            .PADIN(N__37496),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__37489),
            .DIN(N__37488),
            .DOUT(N__37487),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__37489),
            .PADOUT(N__37488),
            .PADIN(N__37487),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11583),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__37480),
            .DIN(N__37479),
            .DOUT(N__37478),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__37480),
            .PADOUT(N__37479),
            .PADIN(N__37478),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24984),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__37471),
            .DIN(N__37470),
            .DOUT(N__37469),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__37471),
            .PADOUT(N__37470),
            .PADIN(N__37469),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__37462),
            .DIN(N__37461),
            .DOUT(N__37460),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__37462),
            .PADOUT(N__37461),
            .PADIN(N__37460),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11577),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__37453),
            .DIN(N__37452),
            .DOUT(N__37451),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__37453),
            .PADOUT(N__37452),
            .PADIN(N__37451),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__28777),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__20221));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__37444),
            .DIN(N__37443),
            .DOUT(N__37442),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__37444),
            .PADOUT(N__37443),
            .PADIN(N__37442),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12051),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__37435),
            .DIN(N__37434),
            .DOUT(N__37433),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__37435),
            .PADOUT(N__37434),
            .PADIN(N__37433),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11742),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__37426),
            .DIN(N__37425),
            .DOUT(N__37424),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__37426),
            .PADOUT(N__37425),
            .PADIN(N__37424),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11754),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__37417),
            .DIN(N__37416),
            .DOUT(N__37415),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__37417),
            .PADOUT(N__37416),
            .PADIN(N__37415),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11688),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__37408),
            .DIN(N__37407),
            .DOUT(N__37406),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__37408),
            .PADOUT(N__37407),
            .PADIN(N__37406),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11733),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__37399),
            .DIN(N__37398),
            .DOUT(N__37397),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__37399),
            .PADOUT(N__37398),
            .PADIN(N__37397),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12000),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__37390),
            .DIN(N__37389),
            .DOUT(N__37388),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__37390),
            .PADOUT(N__37389),
            .PADIN(N__37388),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__37381),
            .DIN(N__37380),
            .DOUT(N__37379),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__37381),
            .PADOUT(N__37380),
            .PADIN(N__37379),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__11568),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__37372),
            .DIN(N__37371),
            .DOUT(N__37370),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__37372),
            .PADOUT(N__37371),
            .PADIN(N__37370),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12090),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__9454 (
            .O(N__37353),
            .I(N__37350));
    LocalMux I__9453 (
            .O(N__37350),
            .I(N__37347));
    Span4Mux_s1_h I__9452 (
            .O(N__37347),
            .I(N__37344));
    Span4Mux_h I__9451 (
            .O(N__37344),
            .I(N__37339));
    CascadeMux I__9450 (
            .O(N__37343),
            .I(N__37336));
    InMux I__9449 (
            .O(N__37342),
            .I(N__37333));
    Span4Mux_h I__9448 (
            .O(N__37339),
            .I(N__37330));
    InMux I__9447 (
            .O(N__37336),
            .I(N__37327));
    LocalMux I__9446 (
            .O(N__37333),
            .I(N__37324));
    Odrv4 I__9445 (
            .O(N__37330),
            .I(M_this_external_address_qZ0Z_12));
    LocalMux I__9444 (
            .O(N__37327),
            .I(M_this_external_address_qZ0Z_12));
    Odrv12 I__9443 (
            .O(N__37324),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__9442 (
            .O(N__37317),
            .I(N__37314));
    LocalMux I__9441 (
            .O(N__37314),
            .I(N__37311));
    Odrv4 I__9440 (
            .O(N__37311),
            .I(M_this_external_address_q_cry_11_THRU_CO));
    InMux I__9439 (
            .O(N__37308),
            .I(M_this_external_address_q_cry_11));
    IoInMux I__9438 (
            .O(N__37305),
            .I(N__37302));
    LocalMux I__9437 (
            .O(N__37302),
            .I(N__37299));
    IoSpan4Mux I__9436 (
            .O(N__37299),
            .I(N__37294));
    CascadeMux I__9435 (
            .O(N__37298),
            .I(N__37291));
    InMux I__9434 (
            .O(N__37297),
            .I(N__37288));
    Sp12to4 I__9433 (
            .O(N__37294),
            .I(N__37285));
    InMux I__9432 (
            .O(N__37291),
            .I(N__37282));
    LocalMux I__9431 (
            .O(N__37288),
            .I(N__37279));
    Odrv12 I__9430 (
            .O(N__37285),
            .I(M_this_external_address_qZ0Z_13));
    LocalMux I__9429 (
            .O(N__37282),
            .I(M_this_external_address_qZ0Z_13));
    Odrv12 I__9428 (
            .O(N__37279),
            .I(M_this_external_address_qZ0Z_13));
    InMux I__9427 (
            .O(N__37272),
            .I(N__37269));
    LocalMux I__9426 (
            .O(N__37269),
            .I(N__37266));
    Odrv4 I__9425 (
            .O(N__37266),
            .I(M_this_external_address_q_cry_12_THRU_CO));
    InMux I__9424 (
            .O(N__37263),
            .I(M_this_external_address_q_cry_12));
    IoInMux I__9423 (
            .O(N__37260),
            .I(N__37257));
    LocalMux I__9422 (
            .O(N__37257),
            .I(N__37254));
    Span4Mux_s3_h I__9421 (
            .O(N__37254),
            .I(N__37249));
    CascadeMux I__9420 (
            .O(N__37253),
            .I(N__37246));
    InMux I__9419 (
            .O(N__37252),
            .I(N__37243));
    Span4Mux_v I__9418 (
            .O(N__37249),
            .I(N__37240));
    InMux I__9417 (
            .O(N__37246),
            .I(N__37237));
    LocalMux I__9416 (
            .O(N__37243),
            .I(N__37234));
    Odrv4 I__9415 (
            .O(N__37240),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__9414 (
            .O(N__37237),
            .I(M_this_external_address_qZ0Z_14));
    Odrv4 I__9413 (
            .O(N__37234),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__9412 (
            .O(N__37227),
            .I(N__37224));
    LocalMux I__9411 (
            .O(N__37224),
            .I(N__37221));
    Odrv4 I__9410 (
            .O(N__37221),
            .I(M_this_external_address_q_cry_13_THRU_CO));
    InMux I__9409 (
            .O(N__37218),
            .I(M_this_external_address_q_cry_13));
    IoInMux I__9408 (
            .O(N__37215),
            .I(N__37212));
    LocalMux I__9407 (
            .O(N__37212),
            .I(N__37209));
    IoSpan4Mux I__9406 (
            .O(N__37209),
            .I(N__37206));
    Span4Mux_s3_h I__9405 (
            .O(N__37206),
            .I(N__37203));
    Span4Mux_v I__9404 (
            .O(N__37203),
            .I(N__37199));
    InMux I__9403 (
            .O(N__37202),
            .I(N__37196));
    Span4Mux_v I__9402 (
            .O(N__37199),
            .I(N__37193));
    LocalMux I__9401 (
            .O(N__37196),
            .I(N__37190));
    Span4Mux_h I__9400 (
            .O(N__37193),
            .I(N__37187));
    Span4Mux_h I__9399 (
            .O(N__37190),
            .I(N__37184));
    Odrv4 I__9398 (
            .O(N__37187),
            .I(M_this_external_address_qZ0Z_15));
    Odrv4 I__9397 (
            .O(N__37184),
            .I(M_this_external_address_qZ0Z_15));
    InMux I__9396 (
            .O(N__37179),
            .I(M_this_external_address_q_cry_14));
    CascadeMux I__9395 (
            .O(N__37176),
            .I(N__37173));
    InMux I__9394 (
            .O(N__37173),
            .I(N__37170));
    LocalMux I__9393 (
            .O(N__37170),
            .I(N__37167));
    Span4Mux_h I__9392 (
            .O(N__37167),
            .I(N__37164));
    Odrv4 I__9391 (
            .O(N__37164),
            .I(M_this_external_address_q_s_15));
    InMux I__9390 (
            .O(N__37161),
            .I(M_this_external_address_q_cry_3));
    IoInMux I__9389 (
            .O(N__37158),
            .I(N__37155));
    LocalMux I__9388 (
            .O(N__37155),
            .I(N__37151));
    InMux I__9387 (
            .O(N__37154),
            .I(N__37148));
    Odrv12 I__9386 (
            .O(N__37151),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__9385 (
            .O(N__37148),
            .I(M_this_external_address_qZ0Z_5));
    InMux I__9384 (
            .O(N__37143),
            .I(M_this_external_address_q_cry_4));
    IoInMux I__9383 (
            .O(N__37140),
            .I(N__37137));
    LocalMux I__9382 (
            .O(N__37137),
            .I(N__37134));
    Span4Mux_s3_h I__9381 (
            .O(N__37134),
            .I(N__37131));
    Span4Mux_v I__9380 (
            .O(N__37131),
            .I(N__37127));
    InMux I__9379 (
            .O(N__37130),
            .I(N__37124));
    Odrv4 I__9378 (
            .O(N__37127),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__9377 (
            .O(N__37124),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__9376 (
            .O(N__37119),
            .I(M_this_external_address_q_cry_5));
    InMux I__9375 (
            .O(N__37116),
            .I(N__37100));
    InMux I__9374 (
            .O(N__37115),
            .I(N__37100));
    InMux I__9373 (
            .O(N__37114),
            .I(N__37097));
    InMux I__9372 (
            .O(N__37113),
            .I(N__37092));
    InMux I__9371 (
            .O(N__37112),
            .I(N__37092));
    InMux I__9370 (
            .O(N__37111),
            .I(N__37083));
    InMux I__9369 (
            .O(N__37110),
            .I(N__37083));
    InMux I__9368 (
            .O(N__37109),
            .I(N__37083));
    InMux I__9367 (
            .O(N__37108),
            .I(N__37083));
    InMux I__9366 (
            .O(N__37107),
            .I(N__37072));
    InMux I__9365 (
            .O(N__37106),
            .I(N__37072));
    InMux I__9364 (
            .O(N__37105),
            .I(N__37072));
    LocalMux I__9363 (
            .O(N__37100),
            .I(N__37069));
    LocalMux I__9362 (
            .O(N__37097),
            .I(N__37066));
    LocalMux I__9361 (
            .O(N__37092),
            .I(N__37063));
    LocalMux I__9360 (
            .O(N__37083),
            .I(N__37060));
    InMux I__9359 (
            .O(N__37082),
            .I(N__37051));
    InMux I__9358 (
            .O(N__37081),
            .I(N__37051));
    InMux I__9357 (
            .O(N__37080),
            .I(N__37051));
    InMux I__9356 (
            .O(N__37079),
            .I(N__37051));
    LocalMux I__9355 (
            .O(N__37072),
            .I(N__37048));
    Span4Mux_v I__9354 (
            .O(N__37069),
            .I(N__37045));
    Span4Mux_v I__9353 (
            .O(N__37066),
            .I(N__37042));
    Span4Mux_h I__9352 (
            .O(N__37063),
            .I(N__37039));
    Span4Mux_v I__9351 (
            .O(N__37060),
            .I(N__37034));
    LocalMux I__9350 (
            .O(N__37051),
            .I(N__37034));
    Span4Mux_h I__9349 (
            .O(N__37048),
            .I(N__37031));
    Span4Mux_h I__9348 (
            .O(N__37045),
            .I(N__37024));
    Span4Mux_h I__9347 (
            .O(N__37042),
            .I(N__37024));
    Span4Mux_h I__9346 (
            .O(N__37039),
            .I(N__37024));
    Sp12to4 I__9345 (
            .O(N__37034),
            .I(N__37021));
    Span4Mux_h I__9344 (
            .O(N__37031),
            .I(N__37018));
    Span4Mux_h I__9343 (
            .O(N__37024),
            .I(N__37015));
    Odrv12 I__9342 (
            .O(N__37021),
            .I(N_49));
    Odrv4 I__9341 (
            .O(N__37018),
            .I(N_49));
    Odrv4 I__9340 (
            .O(N__37015),
            .I(N_49));
    IoInMux I__9339 (
            .O(N__37008),
            .I(N__37005));
    LocalMux I__9338 (
            .O(N__37005),
            .I(N__37002));
    Span4Mux_s2_h I__9337 (
            .O(N__37002),
            .I(N__36999));
    Span4Mux_h I__9336 (
            .O(N__36999),
            .I(N__36996));
    Sp12to4 I__9335 (
            .O(N__36996),
            .I(N__36993));
    Span12Mux_v I__9334 (
            .O(N__36993),
            .I(N__36989));
    InMux I__9333 (
            .O(N__36992),
            .I(N__36986));
    Odrv12 I__9332 (
            .O(N__36989),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__9331 (
            .O(N__36986),
            .I(M_this_external_address_qZ0Z_7));
    InMux I__9330 (
            .O(N__36981),
            .I(M_this_external_address_q_cry_6));
    ClkMux I__9329 (
            .O(N__36978),
            .I(N__36582));
    ClkMux I__9328 (
            .O(N__36977),
            .I(N__36582));
    ClkMux I__9327 (
            .O(N__36976),
            .I(N__36582));
    ClkMux I__9326 (
            .O(N__36975),
            .I(N__36582));
    ClkMux I__9325 (
            .O(N__36974),
            .I(N__36582));
    ClkMux I__9324 (
            .O(N__36973),
            .I(N__36582));
    ClkMux I__9323 (
            .O(N__36972),
            .I(N__36582));
    ClkMux I__9322 (
            .O(N__36971),
            .I(N__36582));
    ClkMux I__9321 (
            .O(N__36970),
            .I(N__36582));
    ClkMux I__9320 (
            .O(N__36969),
            .I(N__36582));
    ClkMux I__9319 (
            .O(N__36968),
            .I(N__36582));
    ClkMux I__9318 (
            .O(N__36967),
            .I(N__36582));
    ClkMux I__9317 (
            .O(N__36966),
            .I(N__36582));
    ClkMux I__9316 (
            .O(N__36965),
            .I(N__36582));
    ClkMux I__9315 (
            .O(N__36964),
            .I(N__36582));
    ClkMux I__9314 (
            .O(N__36963),
            .I(N__36582));
    ClkMux I__9313 (
            .O(N__36962),
            .I(N__36582));
    ClkMux I__9312 (
            .O(N__36961),
            .I(N__36582));
    ClkMux I__9311 (
            .O(N__36960),
            .I(N__36582));
    ClkMux I__9310 (
            .O(N__36959),
            .I(N__36582));
    ClkMux I__9309 (
            .O(N__36958),
            .I(N__36582));
    ClkMux I__9308 (
            .O(N__36957),
            .I(N__36582));
    ClkMux I__9307 (
            .O(N__36956),
            .I(N__36582));
    ClkMux I__9306 (
            .O(N__36955),
            .I(N__36582));
    ClkMux I__9305 (
            .O(N__36954),
            .I(N__36582));
    ClkMux I__9304 (
            .O(N__36953),
            .I(N__36582));
    ClkMux I__9303 (
            .O(N__36952),
            .I(N__36582));
    ClkMux I__9302 (
            .O(N__36951),
            .I(N__36582));
    ClkMux I__9301 (
            .O(N__36950),
            .I(N__36582));
    ClkMux I__9300 (
            .O(N__36949),
            .I(N__36582));
    ClkMux I__9299 (
            .O(N__36948),
            .I(N__36582));
    ClkMux I__9298 (
            .O(N__36947),
            .I(N__36582));
    ClkMux I__9297 (
            .O(N__36946),
            .I(N__36582));
    ClkMux I__9296 (
            .O(N__36945),
            .I(N__36582));
    ClkMux I__9295 (
            .O(N__36944),
            .I(N__36582));
    ClkMux I__9294 (
            .O(N__36943),
            .I(N__36582));
    ClkMux I__9293 (
            .O(N__36942),
            .I(N__36582));
    ClkMux I__9292 (
            .O(N__36941),
            .I(N__36582));
    ClkMux I__9291 (
            .O(N__36940),
            .I(N__36582));
    ClkMux I__9290 (
            .O(N__36939),
            .I(N__36582));
    ClkMux I__9289 (
            .O(N__36938),
            .I(N__36582));
    ClkMux I__9288 (
            .O(N__36937),
            .I(N__36582));
    ClkMux I__9287 (
            .O(N__36936),
            .I(N__36582));
    ClkMux I__9286 (
            .O(N__36935),
            .I(N__36582));
    ClkMux I__9285 (
            .O(N__36934),
            .I(N__36582));
    ClkMux I__9284 (
            .O(N__36933),
            .I(N__36582));
    ClkMux I__9283 (
            .O(N__36932),
            .I(N__36582));
    ClkMux I__9282 (
            .O(N__36931),
            .I(N__36582));
    ClkMux I__9281 (
            .O(N__36930),
            .I(N__36582));
    ClkMux I__9280 (
            .O(N__36929),
            .I(N__36582));
    ClkMux I__9279 (
            .O(N__36928),
            .I(N__36582));
    ClkMux I__9278 (
            .O(N__36927),
            .I(N__36582));
    ClkMux I__9277 (
            .O(N__36926),
            .I(N__36582));
    ClkMux I__9276 (
            .O(N__36925),
            .I(N__36582));
    ClkMux I__9275 (
            .O(N__36924),
            .I(N__36582));
    ClkMux I__9274 (
            .O(N__36923),
            .I(N__36582));
    ClkMux I__9273 (
            .O(N__36922),
            .I(N__36582));
    ClkMux I__9272 (
            .O(N__36921),
            .I(N__36582));
    ClkMux I__9271 (
            .O(N__36920),
            .I(N__36582));
    ClkMux I__9270 (
            .O(N__36919),
            .I(N__36582));
    ClkMux I__9269 (
            .O(N__36918),
            .I(N__36582));
    ClkMux I__9268 (
            .O(N__36917),
            .I(N__36582));
    ClkMux I__9267 (
            .O(N__36916),
            .I(N__36582));
    ClkMux I__9266 (
            .O(N__36915),
            .I(N__36582));
    ClkMux I__9265 (
            .O(N__36914),
            .I(N__36582));
    ClkMux I__9264 (
            .O(N__36913),
            .I(N__36582));
    ClkMux I__9263 (
            .O(N__36912),
            .I(N__36582));
    ClkMux I__9262 (
            .O(N__36911),
            .I(N__36582));
    ClkMux I__9261 (
            .O(N__36910),
            .I(N__36582));
    ClkMux I__9260 (
            .O(N__36909),
            .I(N__36582));
    ClkMux I__9259 (
            .O(N__36908),
            .I(N__36582));
    ClkMux I__9258 (
            .O(N__36907),
            .I(N__36582));
    ClkMux I__9257 (
            .O(N__36906),
            .I(N__36582));
    ClkMux I__9256 (
            .O(N__36905),
            .I(N__36582));
    ClkMux I__9255 (
            .O(N__36904),
            .I(N__36582));
    ClkMux I__9254 (
            .O(N__36903),
            .I(N__36582));
    ClkMux I__9253 (
            .O(N__36902),
            .I(N__36582));
    ClkMux I__9252 (
            .O(N__36901),
            .I(N__36582));
    ClkMux I__9251 (
            .O(N__36900),
            .I(N__36582));
    ClkMux I__9250 (
            .O(N__36899),
            .I(N__36582));
    ClkMux I__9249 (
            .O(N__36898),
            .I(N__36582));
    ClkMux I__9248 (
            .O(N__36897),
            .I(N__36582));
    ClkMux I__9247 (
            .O(N__36896),
            .I(N__36582));
    ClkMux I__9246 (
            .O(N__36895),
            .I(N__36582));
    ClkMux I__9245 (
            .O(N__36894),
            .I(N__36582));
    ClkMux I__9244 (
            .O(N__36893),
            .I(N__36582));
    ClkMux I__9243 (
            .O(N__36892),
            .I(N__36582));
    ClkMux I__9242 (
            .O(N__36891),
            .I(N__36582));
    ClkMux I__9241 (
            .O(N__36890),
            .I(N__36582));
    ClkMux I__9240 (
            .O(N__36889),
            .I(N__36582));
    ClkMux I__9239 (
            .O(N__36888),
            .I(N__36582));
    ClkMux I__9238 (
            .O(N__36887),
            .I(N__36582));
    ClkMux I__9237 (
            .O(N__36886),
            .I(N__36582));
    ClkMux I__9236 (
            .O(N__36885),
            .I(N__36582));
    ClkMux I__9235 (
            .O(N__36884),
            .I(N__36582));
    ClkMux I__9234 (
            .O(N__36883),
            .I(N__36582));
    ClkMux I__9233 (
            .O(N__36882),
            .I(N__36582));
    ClkMux I__9232 (
            .O(N__36881),
            .I(N__36582));
    ClkMux I__9231 (
            .O(N__36880),
            .I(N__36582));
    ClkMux I__9230 (
            .O(N__36879),
            .I(N__36582));
    ClkMux I__9229 (
            .O(N__36878),
            .I(N__36582));
    ClkMux I__9228 (
            .O(N__36877),
            .I(N__36582));
    ClkMux I__9227 (
            .O(N__36876),
            .I(N__36582));
    ClkMux I__9226 (
            .O(N__36875),
            .I(N__36582));
    ClkMux I__9225 (
            .O(N__36874),
            .I(N__36582));
    ClkMux I__9224 (
            .O(N__36873),
            .I(N__36582));
    ClkMux I__9223 (
            .O(N__36872),
            .I(N__36582));
    ClkMux I__9222 (
            .O(N__36871),
            .I(N__36582));
    ClkMux I__9221 (
            .O(N__36870),
            .I(N__36582));
    ClkMux I__9220 (
            .O(N__36869),
            .I(N__36582));
    ClkMux I__9219 (
            .O(N__36868),
            .I(N__36582));
    ClkMux I__9218 (
            .O(N__36867),
            .I(N__36582));
    ClkMux I__9217 (
            .O(N__36866),
            .I(N__36582));
    ClkMux I__9216 (
            .O(N__36865),
            .I(N__36582));
    ClkMux I__9215 (
            .O(N__36864),
            .I(N__36582));
    ClkMux I__9214 (
            .O(N__36863),
            .I(N__36582));
    ClkMux I__9213 (
            .O(N__36862),
            .I(N__36582));
    ClkMux I__9212 (
            .O(N__36861),
            .I(N__36582));
    ClkMux I__9211 (
            .O(N__36860),
            .I(N__36582));
    ClkMux I__9210 (
            .O(N__36859),
            .I(N__36582));
    ClkMux I__9209 (
            .O(N__36858),
            .I(N__36582));
    ClkMux I__9208 (
            .O(N__36857),
            .I(N__36582));
    ClkMux I__9207 (
            .O(N__36856),
            .I(N__36582));
    ClkMux I__9206 (
            .O(N__36855),
            .I(N__36582));
    ClkMux I__9205 (
            .O(N__36854),
            .I(N__36582));
    ClkMux I__9204 (
            .O(N__36853),
            .I(N__36582));
    ClkMux I__9203 (
            .O(N__36852),
            .I(N__36582));
    ClkMux I__9202 (
            .O(N__36851),
            .I(N__36582));
    ClkMux I__9201 (
            .O(N__36850),
            .I(N__36582));
    ClkMux I__9200 (
            .O(N__36849),
            .I(N__36582));
    ClkMux I__9199 (
            .O(N__36848),
            .I(N__36582));
    ClkMux I__9198 (
            .O(N__36847),
            .I(N__36582));
    GlobalMux I__9197 (
            .O(N__36582),
            .I(N__36579));
    gio2CtrlBuf I__9196 (
            .O(N__36579),
            .I(clk_0_c_g));
    CEMux I__9195 (
            .O(N__36576),
            .I(N__36571));
    CEMux I__9194 (
            .O(N__36575),
            .I(N__36568));
    CEMux I__9193 (
            .O(N__36574),
            .I(N__36565));
    LocalMux I__9192 (
            .O(N__36571),
            .I(N__36562));
    LocalMux I__9191 (
            .O(N__36568),
            .I(N__36557));
    LocalMux I__9190 (
            .O(N__36565),
            .I(N__36554));
    Span4Mux_h I__9189 (
            .O(N__36562),
            .I(N__36551));
    CEMux I__9188 (
            .O(N__36561),
            .I(N__36548));
    CEMux I__9187 (
            .O(N__36560),
            .I(N__36545));
    Span4Mux_v I__9186 (
            .O(N__36557),
            .I(N__36540));
    Span4Mux_v I__9185 (
            .O(N__36554),
            .I(N__36540));
    Span4Mux_h I__9184 (
            .O(N__36551),
            .I(N__36535));
    LocalMux I__9183 (
            .O(N__36548),
            .I(N__36535));
    LocalMux I__9182 (
            .O(N__36545),
            .I(N__36532));
    Odrv4 I__9181 (
            .O(N__36540),
            .I(N_47));
    Odrv4 I__9180 (
            .O(N__36535),
            .I(N_47));
    Odrv12 I__9179 (
            .O(N__36532),
            .I(N_47));
    IoInMux I__9178 (
            .O(N__36525),
            .I(N__36522));
    LocalMux I__9177 (
            .O(N__36522),
            .I(N__36519));
    IoSpan4Mux I__9176 (
            .O(N__36519),
            .I(N__36516));
    Span4Mux_s3_v I__9175 (
            .O(N__36516),
            .I(N__36513));
    Span4Mux_h I__9174 (
            .O(N__36513),
            .I(N__36509));
    InMux I__9173 (
            .O(N__36512),
            .I(N__36506));
    Span4Mux_v I__9172 (
            .O(N__36509),
            .I(N__36503));
    LocalMux I__9171 (
            .O(N__36506),
            .I(N__36500));
    Odrv4 I__9170 (
            .O(N__36503),
            .I(M_this_external_address_qZ0Z_8));
    Odrv4 I__9169 (
            .O(N__36500),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__9168 (
            .O(N__36495),
            .I(N__36492));
    LocalMux I__9167 (
            .O(N__36492),
            .I(N__36489));
    Odrv12 I__9166 (
            .O(N__36489),
            .I(M_this_external_address_q_s_8));
    InMux I__9165 (
            .O(N__36486),
            .I(bfn_26_22_0_));
    IoInMux I__9164 (
            .O(N__36483),
            .I(N__36480));
    LocalMux I__9163 (
            .O(N__36480),
            .I(N__36477));
    IoSpan4Mux I__9162 (
            .O(N__36477),
            .I(N__36473));
    InMux I__9161 (
            .O(N__36476),
            .I(N__36470));
    Span4Mux_s1_v I__9160 (
            .O(N__36473),
            .I(N__36467));
    LocalMux I__9159 (
            .O(N__36470),
            .I(N__36464));
    Sp12to4 I__9158 (
            .O(N__36467),
            .I(N__36461));
    Span4Mux_h I__9157 (
            .O(N__36464),
            .I(N__36458));
    Odrv12 I__9156 (
            .O(N__36461),
            .I(M_this_external_address_qZ0Z_9));
    Odrv4 I__9155 (
            .O(N__36458),
            .I(M_this_external_address_qZ0Z_9));
    InMux I__9154 (
            .O(N__36453),
            .I(N__36450));
    LocalMux I__9153 (
            .O(N__36450),
            .I(N__36447));
    Span4Mux_h I__9152 (
            .O(N__36447),
            .I(N__36444));
    Odrv4 I__9151 (
            .O(N__36444),
            .I(M_this_external_address_q_s_9));
    InMux I__9150 (
            .O(N__36441),
            .I(M_this_external_address_q_cry_8));
    IoInMux I__9149 (
            .O(N__36438),
            .I(N__36435));
    LocalMux I__9148 (
            .O(N__36435),
            .I(N__36432));
    IoSpan4Mux I__9147 (
            .O(N__36432),
            .I(N__36429));
    Span4Mux_s3_v I__9146 (
            .O(N__36429),
            .I(N__36425));
    InMux I__9145 (
            .O(N__36428),
            .I(N__36422));
    Span4Mux_v I__9144 (
            .O(N__36425),
            .I(N__36419));
    LocalMux I__9143 (
            .O(N__36422),
            .I(N__36416));
    Odrv4 I__9142 (
            .O(N__36419),
            .I(M_this_external_address_qZ0Z_10));
    Odrv4 I__9141 (
            .O(N__36416),
            .I(M_this_external_address_qZ0Z_10));
    InMux I__9140 (
            .O(N__36411),
            .I(N__36408));
    LocalMux I__9139 (
            .O(N__36408),
            .I(N__36405));
    Odrv4 I__9138 (
            .O(N__36405),
            .I(M_this_external_address_q_s_10));
    InMux I__9137 (
            .O(N__36402),
            .I(M_this_external_address_q_cry_9));
    IoInMux I__9136 (
            .O(N__36399),
            .I(N__36396));
    LocalMux I__9135 (
            .O(N__36396),
            .I(N__36393));
    Span4Mux_s2_v I__9134 (
            .O(N__36393),
            .I(N__36390));
    Span4Mux_v I__9133 (
            .O(N__36390),
            .I(N__36387));
    Span4Mux_v I__9132 (
            .O(N__36387),
            .I(N__36383));
    InMux I__9131 (
            .O(N__36386),
            .I(N__36380));
    Sp12to4 I__9130 (
            .O(N__36383),
            .I(N__36375));
    LocalMux I__9129 (
            .O(N__36380),
            .I(N__36375));
    Odrv12 I__9128 (
            .O(N__36375),
            .I(M_this_external_address_qZ0Z_11));
    InMux I__9127 (
            .O(N__36372),
            .I(N__36369));
    LocalMux I__9126 (
            .O(N__36369),
            .I(N__36366));
    Odrv4 I__9125 (
            .O(N__36366),
            .I(M_this_external_address_q_s_11));
    InMux I__9124 (
            .O(N__36363),
            .I(M_this_external_address_q_cry_10));
    InMux I__9123 (
            .O(N__36360),
            .I(N__36357));
    LocalMux I__9122 (
            .O(N__36357),
            .I(N__36352));
    CascadeMux I__9121 (
            .O(N__36356),
            .I(N__36349));
    InMux I__9120 (
            .O(N__36355),
            .I(N__36345));
    Span4Mux_v I__9119 (
            .O(N__36352),
            .I(N__36341));
    InMux I__9118 (
            .O(N__36349),
            .I(N__36338));
    CascadeMux I__9117 (
            .O(N__36348),
            .I(N__36335));
    LocalMux I__9116 (
            .O(N__36345),
            .I(N__36329));
    InMux I__9115 (
            .O(N__36344),
            .I(N__36326));
    Span4Mux_h I__9114 (
            .O(N__36341),
            .I(N__36318));
    LocalMux I__9113 (
            .O(N__36338),
            .I(N__36318));
    InMux I__9112 (
            .O(N__36335),
            .I(N__36315));
    InMux I__9111 (
            .O(N__36334),
            .I(N__36310));
    InMux I__9110 (
            .O(N__36333),
            .I(N__36307));
    CascadeMux I__9109 (
            .O(N__36332),
            .I(N__36304));
    Span4Mux_v I__9108 (
            .O(N__36329),
            .I(N__36297));
    LocalMux I__9107 (
            .O(N__36326),
            .I(N__36294));
    InMux I__9106 (
            .O(N__36325),
            .I(N__36291));
    InMux I__9105 (
            .O(N__36324),
            .I(N__36288));
    InMux I__9104 (
            .O(N__36323),
            .I(N__36285));
    Span4Mux_v I__9103 (
            .O(N__36318),
            .I(N__36281));
    LocalMux I__9102 (
            .O(N__36315),
            .I(N__36278));
    InMux I__9101 (
            .O(N__36314),
            .I(N__36275));
    InMux I__9100 (
            .O(N__36313),
            .I(N__36272));
    LocalMux I__9099 (
            .O(N__36310),
            .I(N__36267));
    LocalMux I__9098 (
            .O(N__36307),
            .I(N__36267));
    InMux I__9097 (
            .O(N__36304),
            .I(N__36260));
    InMux I__9096 (
            .O(N__36303),
            .I(N__36260));
    InMux I__9095 (
            .O(N__36302),
            .I(N__36260));
    InMux I__9094 (
            .O(N__36301),
            .I(N__36256));
    InMux I__9093 (
            .O(N__36300),
            .I(N__36253));
    Span4Mux_v I__9092 (
            .O(N__36297),
            .I(N__36249));
    Span4Mux_v I__9091 (
            .O(N__36294),
            .I(N__36244));
    LocalMux I__9090 (
            .O(N__36291),
            .I(N__36244));
    LocalMux I__9089 (
            .O(N__36288),
            .I(N__36241));
    LocalMux I__9088 (
            .O(N__36285),
            .I(N__36238));
    InMux I__9087 (
            .O(N__36284),
            .I(N__36235));
    Span4Mux_h I__9086 (
            .O(N__36281),
            .I(N__36222));
    Span4Mux_v I__9085 (
            .O(N__36278),
            .I(N__36222));
    LocalMux I__9084 (
            .O(N__36275),
            .I(N__36222));
    LocalMux I__9083 (
            .O(N__36272),
            .I(N__36222));
    Span4Mux_v I__9082 (
            .O(N__36267),
            .I(N__36222));
    LocalMux I__9081 (
            .O(N__36260),
            .I(N__36222));
    InMux I__9080 (
            .O(N__36259),
            .I(N__36219));
    LocalMux I__9079 (
            .O(N__36256),
            .I(N__36214));
    LocalMux I__9078 (
            .O(N__36253),
            .I(N__36214));
    InMux I__9077 (
            .O(N__36252),
            .I(N__36211));
    Span4Mux_v I__9076 (
            .O(N__36249),
            .I(N__36204));
    Span4Mux_v I__9075 (
            .O(N__36244),
            .I(N__36204));
    Span4Mux_v I__9074 (
            .O(N__36241),
            .I(N__36204));
    Span4Mux_h I__9073 (
            .O(N__36238),
            .I(N__36199));
    LocalMux I__9072 (
            .O(N__36235),
            .I(N__36199));
    Span4Mux_v I__9071 (
            .O(N__36222),
            .I(N__36196));
    LocalMux I__9070 (
            .O(N__36219),
            .I(N__36193));
    Span12Mux_h I__9069 (
            .O(N__36214),
            .I(N__36190));
    LocalMux I__9068 (
            .O(N__36211),
            .I(N__36187));
    Span4Mux_h I__9067 (
            .O(N__36204),
            .I(N__36182));
    Span4Mux_v I__9066 (
            .O(N__36199),
            .I(N__36182));
    Span4Mux_h I__9065 (
            .O(N__36196),
            .I(N__36177));
    Span4Mux_v I__9064 (
            .O(N__36193),
            .I(N__36177));
    Span12Mux_v I__9063 (
            .O(N__36190),
            .I(N__36174));
    Span12Mux_v I__9062 (
            .O(N__36187),
            .I(N__36169));
    Sp12to4 I__9061 (
            .O(N__36182),
            .I(N__36169));
    Span4Mux_h I__9060 (
            .O(N__36177),
            .I(N__36166));
    Odrv12 I__9059 (
            .O(N__36174),
            .I(port_data_c_5));
    Odrv12 I__9058 (
            .O(N__36169),
            .I(port_data_c_5));
    Odrv4 I__9057 (
            .O(N__36166),
            .I(port_data_c_5));
    InMux I__9056 (
            .O(N__36159),
            .I(N__36156));
    LocalMux I__9055 (
            .O(N__36156),
            .I(N__36153));
    Span4Mux_h I__9054 (
            .O(N__36153),
            .I(N__36150));
    Odrv4 I__9053 (
            .O(N__36150),
            .I(M_this_data_tmp_qZ0Z_13));
    CEMux I__9052 (
            .O(N__36147),
            .I(N__36144));
    LocalMux I__9051 (
            .O(N__36144),
            .I(N__36138));
    CEMux I__9050 (
            .O(N__36143),
            .I(N__36135));
    CEMux I__9049 (
            .O(N__36142),
            .I(N__36132));
    CEMux I__9048 (
            .O(N__36141),
            .I(N__36129));
    Span4Mux_h I__9047 (
            .O(N__36138),
            .I(N__36119));
    LocalMux I__9046 (
            .O(N__36135),
            .I(N__36119));
    LocalMux I__9045 (
            .O(N__36132),
            .I(N__36119));
    LocalMux I__9044 (
            .O(N__36129),
            .I(N__36119));
    CEMux I__9043 (
            .O(N__36128),
            .I(N__36116));
    Span4Mux_v I__9042 (
            .O(N__36119),
            .I(N__36113));
    LocalMux I__9041 (
            .O(N__36116),
            .I(N__36110));
    Odrv4 I__9040 (
            .O(N__36113),
            .I(N_1404_0));
    Odrv12 I__9039 (
            .O(N__36110),
            .I(N_1404_0));
    InMux I__9038 (
            .O(N__36105),
            .I(N__36083));
    InMux I__9037 (
            .O(N__36104),
            .I(N__36080));
    InMux I__9036 (
            .O(N__36103),
            .I(N__36077));
    InMux I__9035 (
            .O(N__36102),
            .I(N__36074));
    InMux I__9034 (
            .O(N__36101),
            .I(N__36071));
    InMux I__9033 (
            .O(N__36100),
            .I(N__36068));
    InMux I__9032 (
            .O(N__36099),
            .I(N__36065));
    InMux I__9031 (
            .O(N__36098),
            .I(N__36062));
    InMux I__9030 (
            .O(N__36097),
            .I(N__36059));
    InMux I__9029 (
            .O(N__36096),
            .I(N__36056));
    InMux I__9028 (
            .O(N__36095),
            .I(N__36053));
    InMux I__9027 (
            .O(N__36094),
            .I(N__36048));
    InMux I__9026 (
            .O(N__36093),
            .I(N__36048));
    InMux I__9025 (
            .O(N__36092),
            .I(N__36045));
    InMux I__9024 (
            .O(N__36091),
            .I(N__36042));
    InMux I__9023 (
            .O(N__36090),
            .I(N__36035));
    InMux I__9022 (
            .O(N__36089),
            .I(N__36035));
    InMux I__9021 (
            .O(N__36088),
            .I(N__36035));
    InMux I__9020 (
            .O(N__36087),
            .I(N__36030));
    InMux I__9019 (
            .O(N__36086),
            .I(N__36030));
    LocalMux I__9018 (
            .O(N__36083),
            .I(N__36002));
    LocalMux I__9017 (
            .O(N__36080),
            .I(N__35999));
    LocalMux I__9016 (
            .O(N__36077),
            .I(N__35996));
    LocalMux I__9015 (
            .O(N__36074),
            .I(N__35993));
    LocalMux I__9014 (
            .O(N__36071),
            .I(N__35990));
    LocalMux I__9013 (
            .O(N__36068),
            .I(N__35987));
    LocalMux I__9012 (
            .O(N__36065),
            .I(N__35984));
    LocalMux I__9011 (
            .O(N__36062),
            .I(N__35981));
    LocalMux I__9010 (
            .O(N__36059),
            .I(N__35978));
    LocalMux I__9009 (
            .O(N__36056),
            .I(N__35975));
    LocalMux I__9008 (
            .O(N__36053),
            .I(N__35972));
    LocalMux I__9007 (
            .O(N__36048),
            .I(N__35969));
    LocalMux I__9006 (
            .O(N__36045),
            .I(N__35966));
    LocalMux I__9005 (
            .O(N__36042),
            .I(N__35963));
    LocalMux I__9004 (
            .O(N__36035),
            .I(N__35960));
    LocalMux I__9003 (
            .O(N__36030),
            .I(N__35957));
    SRMux I__9002 (
            .O(N__36029),
            .I(N__35874));
    SRMux I__9001 (
            .O(N__36028),
            .I(N__35874));
    SRMux I__9000 (
            .O(N__36027),
            .I(N__35874));
    SRMux I__8999 (
            .O(N__36026),
            .I(N__35874));
    SRMux I__8998 (
            .O(N__36025),
            .I(N__35874));
    SRMux I__8997 (
            .O(N__36024),
            .I(N__35874));
    SRMux I__8996 (
            .O(N__36023),
            .I(N__35874));
    SRMux I__8995 (
            .O(N__36022),
            .I(N__35874));
    SRMux I__8994 (
            .O(N__36021),
            .I(N__35874));
    SRMux I__8993 (
            .O(N__36020),
            .I(N__35874));
    SRMux I__8992 (
            .O(N__36019),
            .I(N__35874));
    SRMux I__8991 (
            .O(N__36018),
            .I(N__35874));
    SRMux I__8990 (
            .O(N__36017),
            .I(N__35874));
    SRMux I__8989 (
            .O(N__36016),
            .I(N__35874));
    SRMux I__8988 (
            .O(N__36015),
            .I(N__35874));
    SRMux I__8987 (
            .O(N__36014),
            .I(N__35874));
    SRMux I__8986 (
            .O(N__36013),
            .I(N__35874));
    SRMux I__8985 (
            .O(N__36012),
            .I(N__35874));
    SRMux I__8984 (
            .O(N__36011),
            .I(N__35874));
    SRMux I__8983 (
            .O(N__36010),
            .I(N__35874));
    SRMux I__8982 (
            .O(N__36009),
            .I(N__35874));
    SRMux I__8981 (
            .O(N__36008),
            .I(N__35874));
    SRMux I__8980 (
            .O(N__36007),
            .I(N__35874));
    SRMux I__8979 (
            .O(N__36006),
            .I(N__35874));
    SRMux I__8978 (
            .O(N__36005),
            .I(N__35874));
    Glb2LocalMux I__8977 (
            .O(N__36002),
            .I(N__35874));
    Glb2LocalMux I__8976 (
            .O(N__35999),
            .I(N__35874));
    Glb2LocalMux I__8975 (
            .O(N__35996),
            .I(N__35874));
    Glb2LocalMux I__8974 (
            .O(N__35993),
            .I(N__35874));
    Glb2LocalMux I__8973 (
            .O(N__35990),
            .I(N__35874));
    Glb2LocalMux I__8972 (
            .O(N__35987),
            .I(N__35874));
    Glb2LocalMux I__8971 (
            .O(N__35984),
            .I(N__35874));
    Glb2LocalMux I__8970 (
            .O(N__35981),
            .I(N__35874));
    Glb2LocalMux I__8969 (
            .O(N__35978),
            .I(N__35874));
    Glb2LocalMux I__8968 (
            .O(N__35975),
            .I(N__35874));
    Glb2LocalMux I__8967 (
            .O(N__35972),
            .I(N__35874));
    Glb2LocalMux I__8966 (
            .O(N__35969),
            .I(N__35874));
    Glb2LocalMux I__8965 (
            .O(N__35966),
            .I(N__35874));
    Glb2LocalMux I__8964 (
            .O(N__35963),
            .I(N__35874));
    Glb2LocalMux I__8963 (
            .O(N__35960),
            .I(N__35874));
    Glb2LocalMux I__8962 (
            .O(N__35957),
            .I(N__35874));
    GlobalMux I__8961 (
            .O(N__35874),
            .I(N__35871));
    gio2CtrlBuf I__8960 (
            .O(N__35871),
            .I(M_this_reset_cond_out_g_0));
    InMux I__8959 (
            .O(N__35868),
            .I(N__35865));
    LocalMux I__8958 (
            .O(N__35865),
            .I(N__35860));
    InMux I__8957 (
            .O(N__35864),
            .I(N__35857));
    CascadeMux I__8956 (
            .O(N__35863),
            .I(N__35854));
    Span4Mux_h I__8955 (
            .O(N__35860),
            .I(N__35849));
    LocalMux I__8954 (
            .O(N__35857),
            .I(N__35849));
    InMux I__8953 (
            .O(N__35854),
            .I(N__35843));
    Span4Mux_h I__8952 (
            .O(N__35849),
            .I(N__35840));
    InMux I__8951 (
            .O(N__35848),
            .I(N__35835));
    CascadeMux I__8950 (
            .O(N__35847),
            .I(N__35832));
    CascadeMux I__8949 (
            .O(N__35846),
            .I(N__35827));
    LocalMux I__8948 (
            .O(N__35843),
            .I(N__35823));
    Span4Mux_v I__8947 (
            .O(N__35840),
            .I(N__35820));
    InMux I__8946 (
            .O(N__35839),
            .I(N__35817));
    InMux I__8945 (
            .O(N__35838),
            .I(N__35814));
    LocalMux I__8944 (
            .O(N__35835),
            .I(N__35811));
    InMux I__8943 (
            .O(N__35832),
            .I(N__35808));
    CascadeMux I__8942 (
            .O(N__35831),
            .I(N__35805));
    InMux I__8941 (
            .O(N__35830),
            .I(N__35802));
    InMux I__8940 (
            .O(N__35827),
            .I(N__35797));
    InMux I__8939 (
            .O(N__35826),
            .I(N__35797));
    Span4Mux_v I__8938 (
            .O(N__35823),
            .I(N__35794));
    Span4Mux_v I__8937 (
            .O(N__35820),
            .I(N__35791));
    LocalMux I__8936 (
            .O(N__35817),
            .I(N__35788));
    LocalMux I__8935 (
            .O(N__35814),
            .I(N__35785));
    Span4Mux_v I__8934 (
            .O(N__35811),
            .I(N__35782));
    LocalMux I__8933 (
            .O(N__35808),
            .I(N__35779));
    InMux I__8932 (
            .O(N__35805),
            .I(N__35776));
    LocalMux I__8931 (
            .O(N__35802),
            .I(N__35773));
    LocalMux I__8930 (
            .O(N__35797),
            .I(N__35770));
    Span4Mux_h I__8929 (
            .O(N__35794),
            .I(N__35767));
    Span4Mux_v I__8928 (
            .O(N__35791),
            .I(N__35762));
    Span4Mux_h I__8927 (
            .O(N__35788),
            .I(N__35762));
    Span4Mux_h I__8926 (
            .O(N__35785),
            .I(N__35759));
    Span4Mux_v I__8925 (
            .O(N__35782),
            .I(N__35754));
    Span4Mux_h I__8924 (
            .O(N__35779),
            .I(N__35754));
    LocalMux I__8923 (
            .O(N__35776),
            .I(N__35751));
    Span4Mux_h I__8922 (
            .O(N__35773),
            .I(N__35746));
    Span4Mux_v I__8921 (
            .O(N__35770),
            .I(N__35746));
    Span4Mux_h I__8920 (
            .O(N__35767),
            .I(N__35741));
    Span4Mux_v I__8919 (
            .O(N__35762),
            .I(N__35741));
    Sp12to4 I__8918 (
            .O(N__35759),
            .I(N__35738));
    Span4Mux_h I__8917 (
            .O(N__35754),
            .I(N__35735));
    Span12Mux_v I__8916 (
            .O(N__35751),
            .I(N__35730));
    Sp12to4 I__8915 (
            .O(N__35746),
            .I(N__35730));
    Span4Mux_v I__8914 (
            .O(N__35741),
            .I(N__35727));
    Span12Mux_v I__8913 (
            .O(N__35738),
            .I(N__35722));
    Sp12to4 I__8912 (
            .O(N__35735),
            .I(N__35722));
    Span12Mux_h I__8911 (
            .O(N__35730),
            .I(N__35719));
    IoSpan4Mux I__8910 (
            .O(N__35727),
            .I(N__35716));
    Odrv12 I__8909 (
            .O(N__35722),
            .I(port_data_c_3));
    Odrv12 I__8908 (
            .O(N__35719),
            .I(port_data_c_3));
    Odrv4 I__8907 (
            .O(N__35716),
            .I(port_data_c_3));
    CEMux I__8906 (
            .O(N__35709),
            .I(N__35685));
    CEMux I__8905 (
            .O(N__35708),
            .I(N__35682));
    InMux I__8904 (
            .O(N__35707),
            .I(N__35679));
    InMux I__8903 (
            .O(N__35706),
            .I(N__35674));
    InMux I__8902 (
            .O(N__35705),
            .I(N__35674));
    InMux I__8901 (
            .O(N__35704),
            .I(N__35667));
    InMux I__8900 (
            .O(N__35703),
            .I(N__35667));
    InMux I__8899 (
            .O(N__35702),
            .I(N__35667));
    InMux I__8898 (
            .O(N__35701),
            .I(N__35658));
    InMux I__8897 (
            .O(N__35700),
            .I(N__35658));
    InMux I__8896 (
            .O(N__35699),
            .I(N__35658));
    InMux I__8895 (
            .O(N__35698),
            .I(N__35658));
    InMux I__8894 (
            .O(N__35697),
            .I(N__35645));
    InMux I__8893 (
            .O(N__35696),
            .I(N__35645));
    InMux I__8892 (
            .O(N__35695),
            .I(N__35645));
    InMux I__8891 (
            .O(N__35694),
            .I(N__35645));
    InMux I__8890 (
            .O(N__35693),
            .I(N__35645));
    InMux I__8889 (
            .O(N__35692),
            .I(N__35645));
    InMux I__8888 (
            .O(N__35691),
            .I(N__35638));
    InMux I__8887 (
            .O(N__35690),
            .I(N__35631));
    InMux I__8886 (
            .O(N__35689),
            .I(N__35631));
    InMux I__8885 (
            .O(N__35688),
            .I(N__35631));
    LocalMux I__8884 (
            .O(N__35685),
            .I(N__35622));
    LocalMux I__8883 (
            .O(N__35682),
            .I(N__35619));
    LocalMux I__8882 (
            .O(N__35679),
            .I(N__35616));
    LocalMux I__8881 (
            .O(N__35674),
            .I(N__35609));
    LocalMux I__8880 (
            .O(N__35667),
            .I(N__35609));
    LocalMux I__8879 (
            .O(N__35658),
            .I(N__35609));
    LocalMux I__8878 (
            .O(N__35645),
            .I(N__35606));
    InMux I__8877 (
            .O(N__35644),
            .I(N__35601));
    InMux I__8876 (
            .O(N__35643),
            .I(N__35601));
    InMux I__8875 (
            .O(N__35642),
            .I(N__35598));
    InMux I__8874 (
            .O(N__35641),
            .I(N__35595));
    LocalMux I__8873 (
            .O(N__35638),
            .I(N__35592));
    LocalMux I__8872 (
            .O(N__35631),
            .I(N__35589));
    InMux I__8871 (
            .O(N__35630),
            .I(N__35584));
    InMux I__8870 (
            .O(N__35629),
            .I(N__35584));
    InMux I__8869 (
            .O(N__35628),
            .I(N__35577));
    InMux I__8868 (
            .O(N__35627),
            .I(N__35577));
    InMux I__8867 (
            .O(N__35626),
            .I(N__35577));
    InMux I__8866 (
            .O(N__35625),
            .I(N__35574));
    Span4Mux_v I__8865 (
            .O(N__35622),
            .I(N__35571));
    Span4Mux_h I__8864 (
            .O(N__35619),
            .I(N__35568));
    Span4Mux_h I__8863 (
            .O(N__35616),
            .I(N__35559));
    Span4Mux_v I__8862 (
            .O(N__35609),
            .I(N__35559));
    Span4Mux_h I__8861 (
            .O(N__35606),
            .I(N__35559));
    LocalMux I__8860 (
            .O(N__35601),
            .I(N__35559));
    LocalMux I__8859 (
            .O(N__35598),
            .I(N__35554));
    LocalMux I__8858 (
            .O(N__35595),
            .I(N__35554));
    Span4Mux_h I__8857 (
            .O(N__35592),
            .I(N__35545));
    Span4Mux_h I__8856 (
            .O(N__35589),
            .I(N__35545));
    LocalMux I__8855 (
            .O(N__35584),
            .I(N__35545));
    LocalMux I__8854 (
            .O(N__35577),
            .I(N__35545));
    LocalMux I__8853 (
            .O(N__35574),
            .I(N__35542));
    Span4Mux_v I__8852 (
            .O(N__35571),
            .I(N__35535));
    Span4Mux_v I__8851 (
            .O(N__35568),
            .I(N__35535));
    Span4Mux_v I__8850 (
            .O(N__35559),
            .I(N__35532));
    Span4Mux_h I__8849 (
            .O(N__35554),
            .I(N__35525));
    Span4Mux_v I__8848 (
            .O(N__35545),
            .I(N__35525));
    Span4Mux_h I__8847 (
            .O(N__35542),
            .I(N__35525));
    InMux I__8846 (
            .O(N__35541),
            .I(N__35520));
    InMux I__8845 (
            .O(N__35540),
            .I(N__35520));
    Odrv4 I__8844 (
            .O(N__35535),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv4 I__8843 (
            .O(N__35532),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv4 I__8842 (
            .O(N__35525),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    LocalMux I__8841 (
            .O(N__35520),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    InMux I__8840 (
            .O(N__35511),
            .I(N__35508));
    LocalMux I__8839 (
            .O(N__35508),
            .I(N__35505));
    Odrv4 I__8838 (
            .O(N__35505),
            .I(M_this_oam_ram_write_data_27));
    InMux I__8837 (
            .O(N__35502),
            .I(N__35499));
    LocalMux I__8836 (
            .O(N__35499),
            .I(N__35496));
    Odrv4 I__8835 (
            .O(N__35496),
            .I(M_this_external_address_q_3_0_13));
    InMux I__8834 (
            .O(N__35493),
            .I(N__35490));
    LocalMux I__8833 (
            .O(N__35490),
            .I(N__35487));
    Odrv4 I__8832 (
            .O(N__35487),
            .I(N_312_0));
    IoInMux I__8831 (
            .O(N__35484),
            .I(N__35481));
    LocalMux I__8830 (
            .O(N__35481),
            .I(N__35478));
    Span4Mux_s3_v I__8829 (
            .O(N__35478),
            .I(N__35475));
    Sp12to4 I__8828 (
            .O(N__35475),
            .I(N__35472));
    Span12Mux_h I__8827 (
            .O(N__35472),
            .I(N__35468));
    InMux I__8826 (
            .O(N__35471),
            .I(N__35465));
    Odrv12 I__8825 (
            .O(N__35468),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__8824 (
            .O(N__35465),
            .I(M_this_external_address_qZ0Z_0));
    InMux I__8823 (
            .O(N__35460),
            .I(bfn_26_21_0_));
    IoInMux I__8822 (
            .O(N__35457),
            .I(N__35454));
    LocalMux I__8821 (
            .O(N__35454),
            .I(N__35451));
    Span12Mux_s2_v I__8820 (
            .O(N__35451),
            .I(N__35447));
    InMux I__8819 (
            .O(N__35450),
            .I(N__35444));
    Odrv12 I__8818 (
            .O(N__35447),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__8817 (
            .O(N__35444),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__8816 (
            .O(N__35439),
            .I(M_this_external_address_q_cry_0));
    IoInMux I__8815 (
            .O(N__35436),
            .I(N__35433));
    LocalMux I__8814 (
            .O(N__35433),
            .I(N__35430));
    Span4Mux_s1_v I__8813 (
            .O(N__35430),
            .I(N__35427));
    Span4Mux_h I__8812 (
            .O(N__35427),
            .I(N__35424));
    Sp12to4 I__8811 (
            .O(N__35424),
            .I(N__35420));
    InMux I__8810 (
            .O(N__35423),
            .I(N__35417));
    Odrv12 I__8809 (
            .O(N__35420),
            .I(M_this_external_address_qZ0Z_2));
    LocalMux I__8808 (
            .O(N__35417),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__8807 (
            .O(N__35412),
            .I(M_this_external_address_q_cry_1));
    IoInMux I__8806 (
            .O(N__35409),
            .I(N__35406));
    LocalMux I__8805 (
            .O(N__35406),
            .I(N__35403));
    Span4Mux_s2_h I__8804 (
            .O(N__35403),
            .I(N__35400));
    Span4Mux_h I__8803 (
            .O(N__35400),
            .I(N__35397));
    Span4Mux_v I__8802 (
            .O(N__35397),
            .I(N__35393));
    InMux I__8801 (
            .O(N__35396),
            .I(N__35390));
    Odrv4 I__8800 (
            .O(N__35393),
            .I(M_this_external_address_qZ0Z_3));
    LocalMux I__8799 (
            .O(N__35390),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__8798 (
            .O(N__35385),
            .I(M_this_external_address_q_cry_2));
    IoInMux I__8797 (
            .O(N__35382),
            .I(N__35379));
    LocalMux I__8796 (
            .O(N__35379),
            .I(N__35376));
    Span4Mux_s2_h I__8795 (
            .O(N__35376),
            .I(N__35373));
    Span4Mux_h I__8794 (
            .O(N__35373),
            .I(N__35369));
    InMux I__8793 (
            .O(N__35372),
            .I(N__35366));
    Odrv4 I__8792 (
            .O(N__35369),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__8791 (
            .O(N__35366),
            .I(M_this_external_address_qZ0Z_4));
    InMux I__8790 (
            .O(N__35361),
            .I(N__35358));
    LocalMux I__8789 (
            .O(N__35358),
            .I(N__35355));
    Odrv4 I__8788 (
            .O(N__35355),
            .I(\this_vga_signals.N_665_1 ));
    InMux I__8787 (
            .O(N__35352),
            .I(N__35349));
    LocalMux I__8786 (
            .O(N__35349),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3LZ0Z4 ));
    InMux I__8785 (
            .O(N__35346),
            .I(N__35343));
    LocalMux I__8784 (
            .O(N__35343),
            .I(N__35340));
    Odrv12 I__8783 (
            .O(N__35340),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4LZ0Z6 ));
    InMux I__8782 (
            .O(N__35337),
            .I(N__35334));
    LocalMux I__8781 (
            .O(N__35334),
            .I(N__35331));
    Span4Mux_v I__8780 (
            .O(N__35331),
            .I(N__35328));
    Span4Mux_h I__8779 (
            .O(N__35328),
            .I(N__35324));
    InMux I__8778 (
            .O(N__35327),
            .I(N__35321));
    Span4Mux_v I__8777 (
            .O(N__35324),
            .I(N__35318));
    LocalMux I__8776 (
            .O(N__35321),
            .I(N__35315));
    Sp12to4 I__8775 (
            .O(N__35318),
            .I(N__35310));
    Span12Mux_v I__8774 (
            .O(N__35315),
            .I(N__35310));
    Odrv12 I__8773 (
            .O(N__35310),
            .I(port_address_in_3));
    CascadeMux I__8772 (
            .O(N__35307),
            .I(N__35303));
    InMux I__8771 (
            .O(N__35306),
            .I(N__35300));
    InMux I__8770 (
            .O(N__35303),
            .I(N__35297));
    LocalMux I__8769 (
            .O(N__35300),
            .I(N__35292));
    LocalMux I__8768 (
            .O(N__35297),
            .I(N__35292));
    Odrv12 I__8767 (
            .O(N__35292),
            .I(port_address_in_5));
    CascadeMux I__8766 (
            .O(N__35289),
            .I(N__35286));
    InMux I__8765 (
            .O(N__35286),
            .I(N__35280));
    InMux I__8764 (
            .O(N__35285),
            .I(N__35280));
    LocalMux I__8763 (
            .O(N__35280),
            .I(N__35277));
    Span12Mux_v I__8762 (
            .O(N__35277),
            .I(N__35274));
    Odrv12 I__8761 (
            .O(N__35274),
            .I(port_address_in_6));
    InMux I__8760 (
            .O(N__35271),
            .I(N__35265));
    InMux I__8759 (
            .O(N__35270),
            .I(N__35265));
    LocalMux I__8758 (
            .O(N__35265),
            .I(N__35262));
    Span4Mux_v I__8757 (
            .O(N__35262),
            .I(N__35259));
    Span4Mux_h I__8756 (
            .O(N__35259),
            .I(N__35256));
    Odrv4 I__8755 (
            .O(N__35256),
            .I(port_address_in_4));
    InMux I__8754 (
            .O(N__35253),
            .I(N__35250));
    LocalMux I__8753 (
            .O(N__35250),
            .I(N__35247));
    Span4Mux_h I__8752 (
            .O(N__35247),
            .I(N__35244));
    Span4Mux_h I__8751 (
            .O(N__35244),
            .I(N__35241));
    Odrv4 I__8750 (
            .O(N__35241),
            .I(\this_vga_signals.un1_M_this_state_q_19_i_0_o2Z0Z_4 ));
    CascadeMux I__8749 (
            .O(N__35238),
            .I(N__35235));
    InMux I__8748 (
            .O(N__35235),
            .I(N__35230));
    InMux I__8747 (
            .O(N__35234),
            .I(N__35225));
    InMux I__8746 (
            .O(N__35233),
            .I(N__35221));
    LocalMux I__8745 (
            .O(N__35230),
            .I(N__35215));
    InMux I__8744 (
            .O(N__35229),
            .I(N__35212));
    CascadeMux I__8743 (
            .O(N__35228),
            .I(N__35208));
    LocalMux I__8742 (
            .O(N__35225),
            .I(N__35204));
    CascadeMux I__8741 (
            .O(N__35224),
            .I(N__35200));
    LocalMux I__8740 (
            .O(N__35221),
            .I(N__35197));
    InMux I__8739 (
            .O(N__35220),
            .I(N__35194));
    InMux I__8738 (
            .O(N__35219),
            .I(N__35189));
    InMux I__8737 (
            .O(N__35218),
            .I(N__35189));
    Span4Mux_v I__8736 (
            .O(N__35215),
            .I(N__35184));
    LocalMux I__8735 (
            .O(N__35212),
            .I(N__35184));
    InMux I__8734 (
            .O(N__35211),
            .I(N__35179));
    InMux I__8733 (
            .O(N__35208),
            .I(N__35179));
    CascadeMux I__8732 (
            .O(N__35207),
            .I(N__35176));
    Span4Mux_v I__8731 (
            .O(N__35204),
            .I(N__35173));
    InMux I__8730 (
            .O(N__35203),
            .I(N__35169));
    InMux I__8729 (
            .O(N__35200),
            .I(N__35165));
    Span4Mux_v I__8728 (
            .O(N__35197),
            .I(N__35153));
    LocalMux I__8727 (
            .O(N__35194),
            .I(N__35153));
    LocalMux I__8726 (
            .O(N__35189),
            .I(N__35153));
    Span4Mux_h I__8725 (
            .O(N__35184),
            .I(N__35153));
    LocalMux I__8724 (
            .O(N__35179),
            .I(N__35153));
    InMux I__8723 (
            .O(N__35176),
            .I(N__35150));
    Span4Mux_v I__8722 (
            .O(N__35173),
            .I(N__35147));
    CascadeMux I__8721 (
            .O(N__35172),
            .I(N__35144));
    LocalMux I__8720 (
            .O(N__35169),
            .I(N__35141));
    InMux I__8719 (
            .O(N__35168),
            .I(N__35138));
    LocalMux I__8718 (
            .O(N__35165),
            .I(N__35133));
    InMux I__8717 (
            .O(N__35164),
            .I(N__35130));
    Span4Mux_v I__8716 (
            .O(N__35153),
            .I(N__35125));
    LocalMux I__8715 (
            .O(N__35150),
            .I(N__35125));
    Span4Mux_v I__8714 (
            .O(N__35147),
            .I(N__35122));
    InMux I__8713 (
            .O(N__35144),
            .I(N__35119));
    Span4Mux_v I__8712 (
            .O(N__35141),
            .I(N__35114));
    LocalMux I__8711 (
            .O(N__35138),
            .I(N__35114));
    InMux I__8710 (
            .O(N__35137),
            .I(N__35111));
    InMux I__8709 (
            .O(N__35136),
            .I(N__35108));
    Span4Mux_v I__8708 (
            .O(N__35133),
            .I(N__35105));
    LocalMux I__8707 (
            .O(N__35130),
            .I(N__35102));
    Span4Mux_v I__8706 (
            .O(N__35125),
            .I(N__35099));
    Span4Mux_v I__8705 (
            .O(N__35122),
            .I(N__35094));
    LocalMux I__8704 (
            .O(N__35119),
            .I(N__35094));
    Span4Mux_h I__8703 (
            .O(N__35114),
            .I(N__35091));
    LocalMux I__8702 (
            .O(N__35111),
            .I(N__35088));
    LocalMux I__8701 (
            .O(N__35108),
            .I(N__35085));
    Span4Mux_h I__8700 (
            .O(N__35105),
            .I(N__35080));
    Span4Mux_v I__8699 (
            .O(N__35102),
            .I(N__35080));
    Span4Mux_h I__8698 (
            .O(N__35099),
            .I(N__35075));
    Span4Mux_v I__8697 (
            .O(N__35094),
            .I(N__35075));
    Sp12to4 I__8696 (
            .O(N__35091),
            .I(N__35072));
    Span12Mux_s7_v I__8695 (
            .O(N__35088),
            .I(N__35069));
    Span12Mux_h I__8694 (
            .O(N__35085),
            .I(N__35066));
    Span4Mux_h I__8693 (
            .O(N__35080),
            .I(N__35063));
    Span4Mux_v I__8692 (
            .O(N__35075),
            .I(N__35060));
    Span12Mux_v I__8691 (
            .O(N__35072),
            .I(N__35055));
    Span12Mux_h I__8690 (
            .O(N__35069),
            .I(N__35055));
    Span12Mux_v I__8689 (
            .O(N__35066),
            .I(N__35050));
    Sp12to4 I__8688 (
            .O(N__35063),
            .I(N__35050));
    IoSpan4Mux I__8687 (
            .O(N__35060),
            .I(N__35047));
    Odrv12 I__8686 (
            .O(N__35055),
            .I(port_data_c_2));
    Odrv12 I__8685 (
            .O(N__35050),
            .I(port_data_c_2));
    Odrv4 I__8684 (
            .O(N__35047),
            .I(port_data_c_2));
    InMux I__8683 (
            .O(N__35040),
            .I(N__35032));
    InMux I__8682 (
            .O(N__35039),
            .I(N__35029));
    InMux I__8681 (
            .O(N__35038),
            .I(N__35026));
    InMux I__8680 (
            .O(N__35037),
            .I(N__35023));
    InMux I__8679 (
            .O(N__35036),
            .I(N__35020));
    InMux I__8678 (
            .O(N__35035),
            .I(N__35017));
    LocalMux I__8677 (
            .O(N__35032),
            .I(N__35014));
    LocalMux I__8676 (
            .O(N__35029),
            .I(N__35007));
    LocalMux I__8675 (
            .O(N__35026),
            .I(N__35007));
    LocalMux I__8674 (
            .O(N__35023),
            .I(N__35007));
    LocalMux I__8673 (
            .O(N__35020),
            .I(N_760));
    LocalMux I__8672 (
            .O(N__35017),
            .I(N_760));
    Odrv4 I__8671 (
            .O(N__35014),
            .I(N_760));
    Odrv4 I__8670 (
            .O(N__35007),
            .I(N_760));
    InMux I__8669 (
            .O(N__34998),
            .I(N__34988));
    InMux I__8668 (
            .O(N__34997),
            .I(N__34983));
    InMux I__8667 (
            .O(N__34996),
            .I(N__34983));
    InMux I__8666 (
            .O(N__34995),
            .I(N__34980));
    InMux I__8665 (
            .O(N__34994),
            .I(N__34977));
    InMux I__8664 (
            .O(N__34993),
            .I(N__34974));
    InMux I__8663 (
            .O(N__34992),
            .I(N__34971));
    InMux I__8662 (
            .O(N__34991),
            .I(N__34968));
    LocalMux I__8661 (
            .O(N__34988),
            .I(N__34963));
    LocalMux I__8660 (
            .O(N__34983),
            .I(N__34963));
    LocalMux I__8659 (
            .O(N__34980),
            .I(N__34960));
    LocalMux I__8658 (
            .O(N__34977),
            .I(N__34957));
    LocalMux I__8657 (
            .O(N__34974),
            .I(N__34948));
    LocalMux I__8656 (
            .O(N__34971),
            .I(N__34948));
    LocalMux I__8655 (
            .O(N__34968),
            .I(N__34943));
    Span4Mux_v I__8654 (
            .O(N__34963),
            .I(N__34943));
    Span4Mux_v I__8653 (
            .O(N__34960),
            .I(N__34938));
    Span4Mux_v I__8652 (
            .O(N__34957),
            .I(N__34938));
    InMux I__8651 (
            .O(N__34956),
            .I(N__34931));
    InMux I__8650 (
            .O(N__34955),
            .I(N__34931));
    InMux I__8649 (
            .O(N__34954),
            .I(N__34931));
    InMux I__8648 (
            .O(N__34953),
            .I(N__34928));
    Span4Mux_v I__8647 (
            .O(N__34948),
            .I(N__34921));
    Span4Mux_v I__8646 (
            .O(N__34943),
            .I(N__34921));
    Span4Mux_h I__8645 (
            .O(N__34938),
            .I(N__34921));
    LocalMux I__8644 (
            .O(N__34931),
            .I(M_this_sprites_address_qZ0Z_12));
    LocalMux I__8643 (
            .O(N__34928),
            .I(M_this_sprites_address_qZ0Z_12));
    Odrv4 I__8642 (
            .O(N__34921),
            .I(M_this_sprites_address_qZ0Z_12));
    InMux I__8641 (
            .O(N__34914),
            .I(N__34907));
    CascadeMux I__8640 (
            .O(N__34913),
            .I(N__34902));
    InMux I__8639 (
            .O(N__34912),
            .I(N__34899));
    InMux I__8638 (
            .O(N__34911),
            .I(N__34896));
    InMux I__8637 (
            .O(N__34910),
            .I(N__34893));
    LocalMux I__8636 (
            .O(N__34907),
            .I(N__34890));
    InMux I__8635 (
            .O(N__34906),
            .I(N__34886));
    InMux I__8634 (
            .O(N__34905),
            .I(N__34881));
    InMux I__8633 (
            .O(N__34902),
            .I(N__34881));
    LocalMux I__8632 (
            .O(N__34899),
            .I(N__34878));
    LocalMux I__8631 (
            .O(N__34896),
            .I(N__34873));
    LocalMux I__8630 (
            .O(N__34893),
            .I(N__34873));
    Span4Mux_h I__8629 (
            .O(N__34890),
            .I(N__34870));
    InMux I__8628 (
            .O(N__34889),
            .I(N__34867));
    LocalMux I__8627 (
            .O(N__34886),
            .I(N__34864));
    LocalMux I__8626 (
            .O(N__34881),
            .I(N__34861));
    Span4Mux_h I__8625 (
            .O(N__34878),
            .I(N__34858));
    Span4Mux_h I__8624 (
            .O(N__34873),
            .I(N__34853));
    Span4Mux_h I__8623 (
            .O(N__34870),
            .I(N__34853));
    LocalMux I__8622 (
            .O(N__34867),
            .I(N__34850));
    Span4Mux_h I__8621 (
            .O(N__34864),
            .I(N__34847));
    Span4Mux_h I__8620 (
            .O(N__34861),
            .I(N__34840));
    Span4Mux_h I__8619 (
            .O(N__34858),
            .I(N__34840));
    Span4Mux_v I__8618 (
            .O(N__34853),
            .I(N__34840));
    Odrv12 I__8617 (
            .O(N__34850),
            .I(N_25_0));
    Odrv4 I__8616 (
            .O(N__34847),
            .I(N_25_0));
    Odrv4 I__8615 (
            .O(N__34840),
            .I(N_25_0));
    CascadeMux I__8614 (
            .O(N__34833),
            .I(N__34825));
    CascadeMux I__8613 (
            .O(N__34832),
            .I(N__34822));
    InMux I__8612 (
            .O(N__34831),
            .I(N__34815));
    CascadeMux I__8611 (
            .O(N__34830),
            .I(N__34812));
    CascadeMux I__8610 (
            .O(N__34829),
            .I(N__34809));
    CascadeMux I__8609 (
            .O(N__34828),
            .I(N__34806));
    InMux I__8608 (
            .O(N__34825),
            .I(N__34803));
    InMux I__8607 (
            .O(N__34822),
            .I(N__34798));
    InMux I__8606 (
            .O(N__34821),
            .I(N__34798));
    CascadeMux I__8605 (
            .O(N__34820),
            .I(N__34795));
    CascadeMux I__8604 (
            .O(N__34819),
            .I(N__34792));
    InMux I__8603 (
            .O(N__34818),
            .I(N__34789));
    LocalMux I__8602 (
            .O(N__34815),
            .I(N__34786));
    InMux I__8601 (
            .O(N__34812),
            .I(N__34783));
    InMux I__8600 (
            .O(N__34809),
            .I(N__34780));
    InMux I__8599 (
            .O(N__34806),
            .I(N__34777));
    LocalMux I__8598 (
            .O(N__34803),
            .I(N__34772));
    LocalMux I__8597 (
            .O(N__34798),
            .I(N__34772));
    InMux I__8596 (
            .O(N__34795),
            .I(N__34768));
    InMux I__8595 (
            .O(N__34792),
            .I(N__34765));
    LocalMux I__8594 (
            .O(N__34789),
            .I(N__34762));
    Span4Mux_v I__8593 (
            .O(N__34786),
            .I(N__34759));
    LocalMux I__8592 (
            .O(N__34783),
            .I(N__34754));
    LocalMux I__8591 (
            .O(N__34780),
            .I(N__34754));
    LocalMux I__8590 (
            .O(N__34777),
            .I(N__34749));
    Span4Mux_v I__8589 (
            .O(N__34772),
            .I(N__34749));
    InMux I__8588 (
            .O(N__34771),
            .I(N__34745));
    LocalMux I__8587 (
            .O(N__34768),
            .I(N__34742));
    LocalMux I__8586 (
            .O(N__34765),
            .I(N__34739));
    Span4Mux_v I__8585 (
            .O(N__34762),
            .I(N__34730));
    Span4Mux_h I__8584 (
            .O(N__34759),
            .I(N__34730));
    Span4Mux_v I__8583 (
            .O(N__34754),
            .I(N__34730));
    Span4Mux_v I__8582 (
            .O(N__34749),
            .I(N__34730));
    InMux I__8581 (
            .O(N__34748),
            .I(N__34727));
    LocalMux I__8580 (
            .O(N__34745),
            .I(N__34724));
    Span4Mux_v I__8579 (
            .O(N__34742),
            .I(N__34717));
    Span4Mux_v I__8578 (
            .O(N__34739),
            .I(N__34717));
    Span4Mux_h I__8577 (
            .O(N__34730),
            .I(N__34717));
    LocalMux I__8576 (
            .O(N__34727),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__8575 (
            .O(N__34724),
            .I(M_this_sprites_address_qZ0Z_13));
    Odrv4 I__8574 (
            .O(N__34717),
            .I(M_this_sprites_address_qZ0Z_13));
    InMux I__8573 (
            .O(N__34710),
            .I(N__34703));
    InMux I__8572 (
            .O(N__34709),
            .I(N__34703));
    InMux I__8571 (
            .O(N__34708),
            .I(N__34700));
    LocalMux I__8570 (
            .O(N__34703),
            .I(N__34694));
    LocalMux I__8569 (
            .O(N__34700),
            .I(N__34694));
    InMux I__8568 (
            .O(N__34699),
            .I(N__34690));
    Span4Mux_v I__8567 (
            .O(N__34694),
            .I(N__34687));
    InMux I__8566 (
            .O(N__34693),
            .I(N__34684));
    LocalMux I__8565 (
            .O(N__34690),
            .I(N__34679));
    Sp12to4 I__8564 (
            .O(N__34687),
            .I(N__34670));
    LocalMux I__8563 (
            .O(N__34684),
            .I(N__34670));
    InMux I__8562 (
            .O(N__34683),
            .I(N__34667));
    InMux I__8561 (
            .O(N__34682),
            .I(N__34664));
    Span4Mux_h I__8560 (
            .O(N__34679),
            .I(N__34661));
    InMux I__8559 (
            .O(N__34678),
            .I(N__34658));
    CascadeMux I__8558 (
            .O(N__34677),
            .I(N__34655));
    CascadeMux I__8557 (
            .O(N__34676),
            .I(N__34652));
    InMux I__8556 (
            .O(N__34675),
            .I(N__34648));
    Span12Mux_h I__8555 (
            .O(N__34670),
            .I(N__34645));
    LocalMux I__8554 (
            .O(N__34667),
            .I(N__34640));
    LocalMux I__8553 (
            .O(N__34664),
            .I(N__34640));
    Span4Mux_v I__8552 (
            .O(N__34661),
            .I(N__34635));
    LocalMux I__8551 (
            .O(N__34658),
            .I(N__34635));
    InMux I__8550 (
            .O(N__34655),
            .I(N__34632));
    InMux I__8549 (
            .O(N__34652),
            .I(N__34629));
    InMux I__8548 (
            .O(N__34651),
            .I(N__34626));
    LocalMux I__8547 (
            .O(N__34648),
            .I(N__34623));
    Odrv12 I__8546 (
            .O(N__34645),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv12 I__8545 (
            .O(N__34640),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__8544 (
            .O(N__34635),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__8543 (
            .O(N__34632),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__8542 (
            .O(N__34629),
            .I(M_this_sprites_address_qZ0Z_11));
    LocalMux I__8541 (
            .O(N__34626),
            .I(M_this_sprites_address_qZ0Z_11));
    Odrv4 I__8540 (
            .O(N__34623),
            .I(M_this_sprites_address_qZ0Z_11));
    CEMux I__8539 (
            .O(N__34608),
            .I(N__34604));
    CEMux I__8538 (
            .O(N__34607),
            .I(N__34601));
    LocalMux I__8537 (
            .O(N__34604),
            .I(N__34596));
    LocalMux I__8536 (
            .O(N__34601),
            .I(N__34596));
    Span4Mux_v I__8535 (
            .O(N__34596),
            .I(N__34593));
    Odrv4 I__8534 (
            .O(N__34593),
            .I(\this_sprites_ram.mem_WE_6 ));
    InMux I__8533 (
            .O(N__34590),
            .I(N__34587));
    LocalMux I__8532 (
            .O(N__34587),
            .I(N__34584));
    Odrv4 I__8531 (
            .O(N__34584),
            .I(M_this_oam_ram_write_data_14));
    InMux I__8530 (
            .O(N__34581),
            .I(N__34578));
    LocalMux I__8529 (
            .O(N__34578),
            .I(N__34574));
    CascadeMux I__8528 (
            .O(N__34577),
            .I(N__34570));
    Span4Mux_v I__8527 (
            .O(N__34574),
            .I(N__34566));
    InMux I__8526 (
            .O(N__34573),
            .I(N__34561));
    InMux I__8525 (
            .O(N__34570),
            .I(N__34561));
    CascadeMux I__8524 (
            .O(N__34569),
            .I(N__34558));
    Span4Mux_h I__8523 (
            .O(N__34566),
            .I(N__34553));
    LocalMux I__8522 (
            .O(N__34561),
            .I(N__34553));
    InMux I__8521 (
            .O(N__34558),
            .I(N__34549));
    Span4Mux_h I__8520 (
            .O(N__34553),
            .I(N__34546));
    InMux I__8519 (
            .O(N__34552),
            .I(N__34543));
    LocalMux I__8518 (
            .O(N__34549),
            .I(N__34539));
    Span4Mux_h I__8517 (
            .O(N__34546),
            .I(N__34536));
    LocalMux I__8516 (
            .O(N__34543),
            .I(N__34533));
    InMux I__8515 (
            .O(N__34542),
            .I(N__34530));
    Span4Mux_v I__8514 (
            .O(N__34539),
            .I(N__34526));
    Span4Mux_v I__8513 (
            .O(N__34536),
            .I(N__34521));
    Span4Mux_h I__8512 (
            .O(N__34533),
            .I(N__34521));
    LocalMux I__8511 (
            .O(N__34530),
            .I(N__34518));
    InMux I__8510 (
            .O(N__34529),
            .I(N__34515));
    Span4Mux_h I__8509 (
            .O(N__34526),
            .I(N__34510));
    Span4Mux_v I__8508 (
            .O(N__34521),
            .I(N__34507));
    Span4Mux_v I__8507 (
            .O(N__34518),
            .I(N__34504));
    LocalMux I__8506 (
            .O(N__34515),
            .I(N__34501));
    InMux I__8505 (
            .O(N__34514),
            .I(N__34498));
    InMux I__8504 (
            .O(N__34513),
            .I(N__34495));
    Sp12to4 I__8503 (
            .O(N__34510),
            .I(N__34490));
    Sp12to4 I__8502 (
            .O(N__34507),
            .I(N__34490));
    Span4Mux_h I__8501 (
            .O(N__34504),
            .I(N__34485));
    Span4Mux_v I__8500 (
            .O(N__34501),
            .I(N__34485));
    LocalMux I__8499 (
            .O(N__34498),
            .I(N__34482));
    LocalMux I__8498 (
            .O(N__34495),
            .I(N__34479));
    Span12Mux_v I__8497 (
            .O(N__34490),
            .I(N__34470));
    Sp12to4 I__8496 (
            .O(N__34485),
            .I(N__34470));
    Span12Mux_h I__8495 (
            .O(N__34482),
            .I(N__34470));
    Span12Mux_s9_v I__8494 (
            .O(N__34479),
            .I(N__34470));
    Odrv12 I__8493 (
            .O(N__34470),
            .I(port_data_c_7));
    InMux I__8492 (
            .O(N__34467),
            .I(N__34464));
    LocalMux I__8491 (
            .O(N__34464),
            .I(N__34461));
    Span4Mux_h I__8490 (
            .O(N__34461),
            .I(N__34458));
    Odrv4 I__8489 (
            .O(N__34458),
            .I(M_this_data_tmp_qZ0Z_15));
    InMux I__8488 (
            .O(N__34455),
            .I(N__34452));
    LocalMux I__8487 (
            .O(N__34452),
            .I(N__34449));
    Span4Mux_h I__8486 (
            .O(N__34449),
            .I(N__34446));
    Span4Mux_h I__8485 (
            .O(N__34446),
            .I(N__34436));
    InMux I__8484 (
            .O(N__34445),
            .I(N__34433));
    InMux I__8483 (
            .O(N__34444),
            .I(N__34428));
    InMux I__8482 (
            .O(N__34443),
            .I(N__34428));
    CascadeMux I__8481 (
            .O(N__34442),
            .I(N__34425));
    InMux I__8480 (
            .O(N__34441),
            .I(N__34421));
    InMux I__8479 (
            .O(N__34440),
            .I(N__34418));
    CascadeMux I__8478 (
            .O(N__34439),
            .I(N__34414));
    Span4Mux_v I__8477 (
            .O(N__34436),
            .I(N__34407));
    LocalMux I__8476 (
            .O(N__34433),
            .I(N__34407));
    LocalMux I__8475 (
            .O(N__34428),
            .I(N__34407));
    InMux I__8474 (
            .O(N__34425),
            .I(N__34404));
    CascadeMux I__8473 (
            .O(N__34424),
            .I(N__34401));
    LocalMux I__8472 (
            .O(N__34421),
            .I(N__34398));
    LocalMux I__8471 (
            .O(N__34418),
            .I(N__34395));
    InMux I__8470 (
            .O(N__34417),
            .I(N__34392));
    InMux I__8469 (
            .O(N__34414),
            .I(N__34388));
    Span4Mux_v I__8468 (
            .O(N__34407),
            .I(N__34385));
    LocalMux I__8467 (
            .O(N__34404),
            .I(N__34382));
    InMux I__8466 (
            .O(N__34401),
            .I(N__34379));
    Span4Mux_v I__8465 (
            .O(N__34398),
            .I(N__34372));
    Span4Mux_v I__8464 (
            .O(N__34395),
            .I(N__34372));
    LocalMux I__8463 (
            .O(N__34392),
            .I(N__34372));
    InMux I__8462 (
            .O(N__34391),
            .I(N__34369));
    LocalMux I__8461 (
            .O(N__34388),
            .I(N__34366));
    Span4Mux_h I__8460 (
            .O(N__34385),
            .I(N__34359));
    Span4Mux_h I__8459 (
            .O(N__34382),
            .I(N__34359));
    LocalMux I__8458 (
            .O(N__34379),
            .I(N__34359));
    Span4Mux_h I__8457 (
            .O(N__34372),
            .I(N__34354));
    LocalMux I__8456 (
            .O(N__34369),
            .I(N__34354));
    Span12Mux_h I__8455 (
            .O(N__34366),
            .I(N__34351));
    Sp12to4 I__8454 (
            .O(N__34359),
            .I(N__34348));
    Span4Mux_h I__8453 (
            .O(N__34354),
            .I(N__34345));
    Span12Mux_v I__8452 (
            .O(N__34351),
            .I(N__34342));
    Span12Mux_v I__8451 (
            .O(N__34348),
            .I(N__34339));
    Span4Mux_v I__8450 (
            .O(N__34345),
            .I(N__34336));
    Odrv12 I__8449 (
            .O(N__34342),
            .I(port_data_c_6));
    Odrv12 I__8448 (
            .O(N__34339),
            .I(port_data_c_6));
    Odrv4 I__8447 (
            .O(N__34336),
            .I(port_data_c_6));
    InMux I__8446 (
            .O(N__34329),
            .I(N__34326));
    LocalMux I__8445 (
            .O(N__34326),
            .I(N__34323));
    Odrv4 I__8444 (
            .O(N__34323),
            .I(M_this_data_tmp_qZ0Z_14));
    InMux I__8443 (
            .O(N__34320),
            .I(N__34317));
    LocalMux I__8442 (
            .O(N__34317),
            .I(\this_ppu.un2_hscroll_axb_0 ));
    CascadeMux I__8441 (
            .O(N__34314),
            .I(N__34311));
    InMux I__8440 (
            .O(N__34311),
            .I(N__34308));
    LocalMux I__8439 (
            .O(N__34308),
            .I(N__34304));
    CascadeMux I__8438 (
            .O(N__34307),
            .I(N__34298));
    Span4Mux_v I__8437 (
            .O(N__34304),
            .I(N__34294));
    InMux I__8436 (
            .O(N__34303),
            .I(N__34291));
    InMux I__8435 (
            .O(N__34302),
            .I(N__34287));
    InMux I__8434 (
            .O(N__34301),
            .I(N__34284));
    InMux I__8433 (
            .O(N__34298),
            .I(N__34280));
    InMux I__8432 (
            .O(N__34297),
            .I(N__34277));
    Sp12to4 I__8431 (
            .O(N__34294),
            .I(N__34274));
    LocalMux I__8430 (
            .O(N__34291),
            .I(N__34271));
    InMux I__8429 (
            .O(N__34290),
            .I(N__34268));
    LocalMux I__8428 (
            .O(N__34287),
            .I(N__34264));
    LocalMux I__8427 (
            .O(N__34284),
            .I(N__34261));
    InMux I__8426 (
            .O(N__34283),
            .I(N__34258));
    LocalMux I__8425 (
            .O(N__34280),
            .I(N__34255));
    LocalMux I__8424 (
            .O(N__34277),
            .I(N__34252));
    Span12Mux_h I__8423 (
            .O(N__34274),
            .I(N__34249));
    Span4Mux_v I__8422 (
            .O(N__34271),
            .I(N__34244));
    LocalMux I__8421 (
            .O(N__34268),
            .I(N__34244));
    InMux I__8420 (
            .O(N__34267),
            .I(N__34241));
    Sp12to4 I__8419 (
            .O(N__34264),
            .I(N__34236));
    Span12Mux_v I__8418 (
            .O(N__34261),
            .I(N__34236));
    LocalMux I__8417 (
            .O(N__34258),
            .I(N__34231));
    Span12Mux_h I__8416 (
            .O(N__34255),
            .I(N__34231));
    Span4Mux_v I__8415 (
            .O(N__34252),
            .I(N__34228));
    Odrv12 I__8414 (
            .O(N__34249),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__8413 (
            .O(N__34244),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__8412 (
            .O(N__34241),
            .I(M_this_ppu_vram_addr_0));
    Odrv12 I__8411 (
            .O(N__34236),
            .I(M_this_ppu_vram_addr_0));
    Odrv12 I__8410 (
            .O(N__34231),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__8409 (
            .O(N__34228),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__8408 (
            .O(N__34215),
            .I(N__34210));
    CascadeMux I__8407 (
            .O(N__34214),
            .I(N__34207));
    CascadeMux I__8406 (
            .O(N__34213),
            .I(N__34204));
    InMux I__8405 (
            .O(N__34210),
            .I(N__34200));
    InMux I__8404 (
            .O(N__34207),
            .I(N__34197));
    InMux I__8403 (
            .O(N__34204),
            .I(N__34194));
    CascadeMux I__8402 (
            .O(N__34203),
            .I(N__34191));
    LocalMux I__8401 (
            .O(N__34200),
            .I(N__34185));
    LocalMux I__8400 (
            .O(N__34197),
            .I(N__34185));
    LocalMux I__8399 (
            .O(N__34194),
            .I(N__34182));
    InMux I__8398 (
            .O(N__34191),
            .I(N__34179));
    CascadeMux I__8397 (
            .O(N__34190),
            .I(N__34176));
    Span4Mux_v I__8396 (
            .O(N__34185),
            .I(N__34167));
    Span4Mux_h I__8395 (
            .O(N__34182),
            .I(N__34167));
    LocalMux I__8394 (
            .O(N__34179),
            .I(N__34167));
    InMux I__8393 (
            .O(N__34176),
            .I(N__34164));
    CascadeMux I__8392 (
            .O(N__34175),
            .I(N__34161));
    CascadeMux I__8391 (
            .O(N__34174),
            .I(N__34158));
    Span4Mux_v I__8390 (
            .O(N__34167),
            .I(N__34153));
    LocalMux I__8389 (
            .O(N__34164),
            .I(N__34150));
    InMux I__8388 (
            .O(N__34161),
            .I(N__34147));
    InMux I__8387 (
            .O(N__34158),
            .I(N__34144));
    CascadeMux I__8386 (
            .O(N__34157),
            .I(N__34141));
    CascadeMux I__8385 (
            .O(N__34156),
            .I(N__34138));
    Span4Mux_h I__8384 (
            .O(N__34153),
            .I(N__34132));
    Span4Mux_s3_v I__8383 (
            .O(N__34150),
            .I(N__34125));
    LocalMux I__8382 (
            .O(N__34147),
            .I(N__34125));
    LocalMux I__8381 (
            .O(N__34144),
            .I(N__34125));
    InMux I__8380 (
            .O(N__34141),
            .I(N__34122));
    InMux I__8379 (
            .O(N__34138),
            .I(N__34119));
    CascadeMux I__8378 (
            .O(N__34137),
            .I(N__34116));
    CascadeMux I__8377 (
            .O(N__34136),
            .I(N__34113));
    CascadeMux I__8376 (
            .O(N__34135),
            .I(N__34108));
    Span4Mux_h I__8375 (
            .O(N__34132),
            .I(N__34105));
    Span4Mux_v I__8374 (
            .O(N__34125),
            .I(N__34098));
    LocalMux I__8373 (
            .O(N__34122),
            .I(N__34098));
    LocalMux I__8372 (
            .O(N__34119),
            .I(N__34098));
    InMux I__8371 (
            .O(N__34116),
            .I(N__34095));
    InMux I__8370 (
            .O(N__34113),
            .I(N__34092));
    CascadeMux I__8369 (
            .O(N__34112),
            .I(N__34089));
    CascadeMux I__8368 (
            .O(N__34111),
            .I(N__34086));
    InMux I__8367 (
            .O(N__34108),
            .I(N__34082));
    Span4Mux_h I__8366 (
            .O(N__34105),
            .I(N__34079));
    Span4Mux_v I__8365 (
            .O(N__34098),
            .I(N__34072));
    LocalMux I__8364 (
            .O(N__34095),
            .I(N__34072));
    LocalMux I__8363 (
            .O(N__34092),
            .I(N__34072));
    InMux I__8362 (
            .O(N__34089),
            .I(N__34069));
    InMux I__8361 (
            .O(N__34086),
            .I(N__34066));
    CascadeMux I__8360 (
            .O(N__34085),
            .I(N__34063));
    LocalMux I__8359 (
            .O(N__34082),
            .I(N__34059));
    Span4Mux_h I__8358 (
            .O(N__34079),
            .I(N__34050));
    Span4Mux_v I__8357 (
            .O(N__34072),
            .I(N__34050));
    LocalMux I__8356 (
            .O(N__34069),
            .I(N__34050));
    LocalMux I__8355 (
            .O(N__34066),
            .I(N__34050));
    InMux I__8354 (
            .O(N__34063),
            .I(N__34047));
    CascadeMux I__8353 (
            .O(N__34062),
            .I(N__34044));
    Span4Mux_h I__8352 (
            .O(N__34059),
            .I(N__34037));
    Span4Mux_v I__8351 (
            .O(N__34050),
            .I(N__34037));
    LocalMux I__8350 (
            .O(N__34047),
            .I(N__34037));
    InMux I__8349 (
            .O(N__34044),
            .I(N__34034));
    Odrv4 I__8348 (
            .O(N__34037),
            .I(M_this_ppu_sprites_addr_0));
    LocalMux I__8347 (
            .O(N__34034),
            .I(M_this_ppu_sprites_addr_0));
    InMux I__8346 (
            .O(N__34029),
            .I(N__34026));
    LocalMux I__8345 (
            .O(N__34026),
            .I(N__34023));
    Odrv12 I__8344 (
            .O(N__34023),
            .I(M_this_data_tmp_qZ0Z_19));
    CEMux I__8343 (
            .O(N__34020),
            .I(N__34015));
    CEMux I__8342 (
            .O(N__34019),
            .I(N__34012));
    CEMux I__8341 (
            .O(N__34018),
            .I(N__34009));
    LocalMux I__8340 (
            .O(N__34015),
            .I(N__34006));
    LocalMux I__8339 (
            .O(N__34012),
            .I(N__34002));
    LocalMux I__8338 (
            .O(N__34009),
            .I(N__33999));
    Span4Mux_v I__8337 (
            .O(N__34006),
            .I(N__33996));
    CEMux I__8336 (
            .O(N__34005),
            .I(N__33993));
    Span4Mux_v I__8335 (
            .O(N__34002),
            .I(N__33990));
    Span4Mux_v I__8334 (
            .O(N__33999),
            .I(N__33987));
    Span4Mux_v I__8333 (
            .O(N__33996),
            .I(N__33982));
    LocalMux I__8332 (
            .O(N__33993),
            .I(N__33982));
    Odrv4 I__8331 (
            .O(N__33990),
            .I(N_1396_0));
    Odrv4 I__8330 (
            .O(N__33987),
            .I(N_1396_0));
    Odrv4 I__8329 (
            .O(N__33982),
            .I(N_1396_0));
    InMux I__8328 (
            .O(N__33975),
            .I(N__33972));
    LocalMux I__8327 (
            .O(N__33972),
            .I(N__33969));
    Span4Mux_v I__8326 (
            .O(N__33969),
            .I(N__33966));
    Span4Mux_v I__8325 (
            .O(N__33966),
            .I(N__33963));
    Odrv4 I__8324 (
            .O(N__33963),
            .I(M_this_oam_ram_read_data_0));
    InMux I__8323 (
            .O(N__33960),
            .I(N__33957));
    LocalMux I__8322 (
            .O(N__33957),
            .I(N__33954));
    Span4Mux_v I__8321 (
            .O(N__33954),
            .I(N__33951));
    Sp12to4 I__8320 (
            .O(N__33951),
            .I(N__33948));
    Span12Mux_h I__8319 (
            .O(N__33948),
            .I(N__33945));
    Span12Mux_v I__8318 (
            .O(N__33945),
            .I(N__33942));
    Odrv12 I__8317 (
            .O(N__33942),
            .I(M_this_map_ram_read_data_0));
    CascadeMux I__8316 (
            .O(N__33939),
            .I(N__33936));
    InMux I__8315 (
            .O(N__33936),
            .I(N__33928));
    CascadeMux I__8314 (
            .O(N__33935),
            .I(N__33924));
    CascadeMux I__8313 (
            .O(N__33934),
            .I(N__33921));
    CascadeMux I__8312 (
            .O(N__33933),
            .I(N__33918));
    CascadeMux I__8311 (
            .O(N__33932),
            .I(N__33914));
    CascadeMux I__8310 (
            .O(N__33931),
            .I(N__33911));
    LocalMux I__8309 (
            .O(N__33928),
            .I(N__33908));
    CascadeMux I__8308 (
            .O(N__33927),
            .I(N__33903));
    InMux I__8307 (
            .O(N__33924),
            .I(N__33898));
    InMux I__8306 (
            .O(N__33921),
            .I(N__33898));
    InMux I__8305 (
            .O(N__33918),
            .I(N__33894));
    InMux I__8304 (
            .O(N__33917),
            .I(N__33889));
    InMux I__8303 (
            .O(N__33914),
            .I(N__33889));
    InMux I__8302 (
            .O(N__33911),
            .I(N__33885));
    Span4Mux_v I__8301 (
            .O(N__33908),
            .I(N__33882));
    InMux I__8300 (
            .O(N__33907),
            .I(N__33875));
    InMux I__8299 (
            .O(N__33906),
            .I(N__33875));
    InMux I__8298 (
            .O(N__33903),
            .I(N__33875));
    LocalMux I__8297 (
            .O(N__33898),
            .I(N__33872));
    CascadeMux I__8296 (
            .O(N__33897),
            .I(N__33869));
    LocalMux I__8295 (
            .O(N__33894),
            .I(N__33864));
    LocalMux I__8294 (
            .O(N__33889),
            .I(N__33864));
    CascadeMux I__8293 (
            .O(N__33888),
            .I(N__33860));
    LocalMux I__8292 (
            .O(N__33885),
            .I(N__33857));
    Span4Mux_h I__8291 (
            .O(N__33882),
            .I(N__33850));
    LocalMux I__8290 (
            .O(N__33875),
            .I(N__33850));
    Span4Mux_h I__8289 (
            .O(N__33872),
            .I(N__33850));
    InMux I__8288 (
            .O(N__33869),
            .I(N__33847));
    Span4Mux_v I__8287 (
            .O(N__33864),
            .I(N__33841));
    InMux I__8286 (
            .O(N__33863),
            .I(N__33836));
    InMux I__8285 (
            .O(N__33860),
            .I(N__33836));
    Span4Mux_h I__8284 (
            .O(N__33857),
            .I(N__33829));
    Span4Mux_v I__8283 (
            .O(N__33850),
            .I(N__33829));
    LocalMux I__8282 (
            .O(N__33847),
            .I(N__33829));
    CascadeMux I__8281 (
            .O(N__33846),
            .I(N__33826));
    CascadeMux I__8280 (
            .O(N__33845),
            .I(N__33823));
    InMux I__8279 (
            .O(N__33844),
            .I(N__33820));
    Span4Mux_h I__8278 (
            .O(N__33841),
            .I(N__33817));
    LocalMux I__8277 (
            .O(N__33836),
            .I(N__33814));
    Span4Mux_h I__8276 (
            .O(N__33829),
            .I(N__33811));
    InMux I__8275 (
            .O(N__33826),
            .I(N__33808));
    InMux I__8274 (
            .O(N__33823),
            .I(N__33805));
    LocalMux I__8273 (
            .O(N__33820),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__8272 (
            .O(N__33817),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__8271 (
            .O(N__33814),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__8270 (
            .O(N__33811),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    LocalMux I__8269 (
            .O(N__33808),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    LocalMux I__8268 (
            .O(N__33805),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    InMux I__8267 (
            .O(N__33792),
            .I(N__33787));
    InMux I__8266 (
            .O(N__33791),
            .I(N__33781));
    InMux I__8265 (
            .O(N__33790),
            .I(N__33778));
    LocalMux I__8264 (
            .O(N__33787),
            .I(N__33768));
    InMux I__8263 (
            .O(N__33786),
            .I(N__33761));
    InMux I__8262 (
            .O(N__33785),
            .I(N__33761));
    InMux I__8261 (
            .O(N__33784),
            .I(N__33761));
    LocalMux I__8260 (
            .O(N__33781),
            .I(N__33757));
    LocalMux I__8259 (
            .O(N__33778),
            .I(N__33754));
    InMux I__8258 (
            .O(N__33777),
            .I(N__33749));
    InMux I__8257 (
            .O(N__33776),
            .I(N__33749));
    InMux I__8256 (
            .O(N__33775),
            .I(N__33743));
    InMux I__8255 (
            .O(N__33774),
            .I(N__33743));
    InMux I__8254 (
            .O(N__33773),
            .I(N__33738));
    InMux I__8253 (
            .O(N__33772),
            .I(N__33738));
    InMux I__8252 (
            .O(N__33771),
            .I(N__33735));
    Span4Mux_v I__8251 (
            .O(N__33768),
            .I(N__33732));
    LocalMux I__8250 (
            .O(N__33761),
            .I(N__33729));
    InMux I__8249 (
            .O(N__33760),
            .I(N__33726));
    Span4Mux_v I__8248 (
            .O(N__33757),
            .I(N__33720));
    Span4Mux_h I__8247 (
            .O(N__33754),
            .I(N__33720));
    LocalMux I__8246 (
            .O(N__33749),
            .I(N__33717));
    InMux I__8245 (
            .O(N__33748),
            .I(N__33714));
    LocalMux I__8244 (
            .O(N__33743),
            .I(N__33710));
    LocalMux I__8243 (
            .O(N__33738),
            .I(N__33707));
    LocalMux I__8242 (
            .O(N__33735),
            .I(N__33704));
    Span4Mux_h I__8241 (
            .O(N__33732),
            .I(N__33697));
    Span4Mux_v I__8240 (
            .O(N__33729),
            .I(N__33697));
    LocalMux I__8239 (
            .O(N__33726),
            .I(N__33697));
    InMux I__8238 (
            .O(N__33725),
            .I(N__33694));
    Span4Mux_h I__8237 (
            .O(N__33720),
            .I(N__33687));
    Span4Mux_v I__8236 (
            .O(N__33717),
            .I(N__33687));
    LocalMux I__8235 (
            .O(N__33714),
            .I(N__33687));
    InMux I__8234 (
            .O(N__33713),
            .I(N__33684));
    Span4Mux_h I__8233 (
            .O(N__33710),
            .I(N__33675));
    Span4Mux_v I__8232 (
            .O(N__33707),
            .I(N__33675));
    Span4Mux_h I__8231 (
            .O(N__33704),
            .I(N__33675));
    Span4Mux_v I__8230 (
            .O(N__33697),
            .I(N__33675));
    LocalMux I__8229 (
            .O(N__33694),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    Odrv4 I__8228 (
            .O(N__33687),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__8227 (
            .O(N__33684),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    Odrv4 I__8226 (
            .O(N__33675),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    CascadeMux I__8225 (
            .O(N__33666),
            .I(N__33662));
    CascadeMux I__8224 (
            .O(N__33665),
            .I(N__33659));
    InMux I__8223 (
            .O(N__33662),
            .I(N__33653));
    InMux I__8222 (
            .O(N__33659),
            .I(N__33650));
    CascadeMux I__8221 (
            .O(N__33658),
            .I(N__33647));
    CascadeMux I__8220 (
            .O(N__33657),
            .I(N__33643));
    CascadeMux I__8219 (
            .O(N__33656),
            .I(N__33640));
    LocalMux I__8218 (
            .O(N__33653),
            .I(N__33635));
    LocalMux I__8217 (
            .O(N__33650),
            .I(N__33632));
    InMux I__8216 (
            .O(N__33647),
            .I(N__33629));
    CascadeMux I__8215 (
            .O(N__33646),
            .I(N__33626));
    InMux I__8214 (
            .O(N__33643),
            .I(N__33623));
    InMux I__8213 (
            .O(N__33640),
            .I(N__33620));
    CascadeMux I__8212 (
            .O(N__33639),
            .I(N__33617));
    CascadeMux I__8211 (
            .O(N__33638),
            .I(N__33614));
    Span4Mux_v I__8210 (
            .O(N__33635),
            .I(N__33605));
    Span4Mux_h I__8209 (
            .O(N__33632),
            .I(N__33605));
    LocalMux I__8208 (
            .O(N__33629),
            .I(N__33605));
    InMux I__8207 (
            .O(N__33626),
            .I(N__33602));
    LocalMux I__8206 (
            .O(N__33623),
            .I(N__33595));
    LocalMux I__8205 (
            .O(N__33620),
            .I(N__33595));
    InMux I__8204 (
            .O(N__33617),
            .I(N__33592));
    InMux I__8203 (
            .O(N__33614),
            .I(N__33589));
    CascadeMux I__8202 (
            .O(N__33613),
            .I(N__33586));
    CascadeMux I__8201 (
            .O(N__33612),
            .I(N__33583));
    Span4Mux_v I__8200 (
            .O(N__33605),
            .I(N__33576));
    LocalMux I__8199 (
            .O(N__33602),
            .I(N__33576));
    CascadeMux I__8198 (
            .O(N__33601),
            .I(N__33573));
    CascadeMux I__8197 (
            .O(N__33600),
            .I(N__33570));
    Span4Mux_v I__8196 (
            .O(N__33595),
            .I(N__33563));
    LocalMux I__8195 (
            .O(N__33592),
            .I(N__33563));
    LocalMux I__8194 (
            .O(N__33589),
            .I(N__33563));
    InMux I__8193 (
            .O(N__33586),
            .I(N__33560));
    InMux I__8192 (
            .O(N__33583),
            .I(N__33557));
    CascadeMux I__8191 (
            .O(N__33582),
            .I(N__33554));
    CascadeMux I__8190 (
            .O(N__33581),
            .I(N__33551));
    Span4Mux_v I__8189 (
            .O(N__33576),
            .I(N__33547));
    InMux I__8188 (
            .O(N__33573),
            .I(N__33544));
    InMux I__8187 (
            .O(N__33570),
            .I(N__33541));
    Span4Mux_v I__8186 (
            .O(N__33563),
            .I(N__33534));
    LocalMux I__8185 (
            .O(N__33560),
            .I(N__33534));
    LocalMux I__8184 (
            .O(N__33557),
            .I(N__33534));
    InMux I__8183 (
            .O(N__33554),
            .I(N__33531));
    InMux I__8182 (
            .O(N__33551),
            .I(N__33528));
    CascadeMux I__8181 (
            .O(N__33550),
            .I(N__33525));
    Sp12to4 I__8180 (
            .O(N__33547),
            .I(N__33521));
    LocalMux I__8179 (
            .O(N__33544),
            .I(N__33516));
    LocalMux I__8178 (
            .O(N__33541),
            .I(N__33516));
    Span4Mux_v I__8177 (
            .O(N__33534),
            .I(N__33509));
    LocalMux I__8176 (
            .O(N__33531),
            .I(N__33509));
    LocalMux I__8175 (
            .O(N__33528),
            .I(N__33509));
    InMux I__8174 (
            .O(N__33525),
            .I(N__33506));
    CascadeMux I__8173 (
            .O(N__33524),
            .I(N__33503));
    Span12Mux_h I__8172 (
            .O(N__33521),
            .I(N__33500));
    Span4Mux_v I__8171 (
            .O(N__33516),
            .I(N__33493));
    Span4Mux_v I__8170 (
            .O(N__33509),
            .I(N__33493));
    LocalMux I__8169 (
            .O(N__33506),
            .I(N__33493));
    InMux I__8168 (
            .O(N__33503),
            .I(N__33490));
    Odrv12 I__8167 (
            .O(N__33500),
            .I(M_this_ppu_sprites_addr_6));
    Odrv4 I__8166 (
            .O(N__33493),
            .I(M_this_ppu_sprites_addr_6));
    LocalMux I__8165 (
            .O(N__33490),
            .I(M_this_ppu_sprites_addr_6));
    CEMux I__8164 (
            .O(N__33483),
            .I(N__33479));
    CEMux I__8163 (
            .O(N__33482),
            .I(N__33476));
    LocalMux I__8162 (
            .O(N__33479),
            .I(N__33473));
    LocalMux I__8161 (
            .O(N__33476),
            .I(N__33470));
    Span4Mux_v I__8160 (
            .O(N__33473),
            .I(N__33467));
    Span4Mux_v I__8159 (
            .O(N__33470),
            .I(N__33464));
    Odrv4 I__8158 (
            .O(N__33467),
            .I(\this_sprites_ram.mem_WE_14 ));
    Odrv4 I__8157 (
            .O(N__33464),
            .I(\this_sprites_ram.mem_WE_14 ));
    CEMux I__8156 (
            .O(N__33459),
            .I(N__33455));
    CEMux I__8155 (
            .O(N__33458),
            .I(N__33452));
    LocalMux I__8154 (
            .O(N__33455),
            .I(N__33449));
    LocalMux I__8153 (
            .O(N__33452),
            .I(N__33446));
    Span4Mux_v I__8152 (
            .O(N__33449),
            .I(N__33443));
    Span4Mux_v I__8151 (
            .O(N__33446),
            .I(N__33440));
    Span4Mux_h I__8150 (
            .O(N__33443),
            .I(N__33437));
    Odrv4 I__8149 (
            .O(N__33440),
            .I(\this_sprites_ram.mem_WE_12 ));
    Odrv4 I__8148 (
            .O(N__33437),
            .I(\this_sprites_ram.mem_WE_12 ));
    CEMux I__8147 (
            .O(N__33432),
            .I(N__33429));
    LocalMux I__8146 (
            .O(N__33429),
            .I(N__33425));
    CEMux I__8145 (
            .O(N__33428),
            .I(N__33422));
    Span4Mux_h I__8144 (
            .O(N__33425),
            .I(N__33419));
    LocalMux I__8143 (
            .O(N__33422),
            .I(N__33416));
    Odrv4 I__8142 (
            .O(N__33419),
            .I(\this_sprites_ram.mem_WE_0 ));
    Odrv4 I__8141 (
            .O(N__33416),
            .I(\this_sprites_ram.mem_WE_0 ));
    InMux I__8140 (
            .O(N__33411),
            .I(N__33408));
    LocalMux I__8139 (
            .O(N__33408),
            .I(N__33404));
    InMux I__8138 (
            .O(N__33407),
            .I(N__33401));
    Span4Mux_v I__8137 (
            .O(N__33404),
            .I(N__33395));
    LocalMux I__8136 (
            .O(N__33401),
            .I(N__33395));
    CascadeMux I__8135 (
            .O(N__33400),
            .I(N__33392));
    Span4Mux_v I__8134 (
            .O(N__33395),
            .I(N__33388));
    InMux I__8133 (
            .O(N__33392),
            .I(N__33385));
    CascadeMux I__8132 (
            .O(N__33391),
            .I(N__33382));
    Span4Mux_v I__8131 (
            .O(N__33388),
            .I(N__33379));
    LocalMux I__8130 (
            .O(N__33385),
            .I(N__33376));
    InMux I__8129 (
            .O(N__33382),
            .I(N__33373));
    Span4Mux_v I__8128 (
            .O(N__33379),
            .I(N__33364));
    Span4Mux_h I__8127 (
            .O(N__33376),
            .I(N__33364));
    LocalMux I__8126 (
            .O(N__33373),
            .I(N__33364));
    CascadeMux I__8125 (
            .O(N__33372),
            .I(N__33361));
    InMux I__8124 (
            .O(N__33371),
            .I(N__33356));
    Span4Mux_v I__8123 (
            .O(N__33364),
            .I(N__33351));
    InMux I__8122 (
            .O(N__33361),
            .I(N__33348));
    CascadeMux I__8121 (
            .O(N__33360),
            .I(N__33345));
    InMux I__8120 (
            .O(N__33359),
            .I(N__33342));
    LocalMux I__8119 (
            .O(N__33356),
            .I(N__33339));
    InMux I__8118 (
            .O(N__33355),
            .I(N__33334));
    InMux I__8117 (
            .O(N__33354),
            .I(N__33334));
    Span4Mux_v I__8116 (
            .O(N__33351),
            .I(N__33329));
    LocalMux I__8115 (
            .O(N__33348),
            .I(N__33329));
    InMux I__8114 (
            .O(N__33345),
            .I(N__33326));
    LocalMux I__8113 (
            .O(N__33342),
            .I(N__33323));
    Span4Mux_v I__8112 (
            .O(N__33339),
            .I(N__33320));
    LocalMux I__8111 (
            .O(N__33334),
            .I(N__33317));
    Span4Mux_h I__8110 (
            .O(N__33329),
            .I(N__33312));
    LocalMux I__8109 (
            .O(N__33326),
            .I(N__33312));
    Span12Mux_h I__8108 (
            .O(N__33323),
            .I(N__33308));
    Sp12to4 I__8107 (
            .O(N__33320),
            .I(N__33305));
    Span4Mux_v I__8106 (
            .O(N__33317),
            .I(N__33302));
    Span4Mux_v I__8105 (
            .O(N__33312),
            .I(N__33299));
    InMux I__8104 (
            .O(N__33311),
            .I(N__33296));
    Span12Mux_v I__8103 (
            .O(N__33308),
            .I(N__33293));
    Span12Mux_v I__8102 (
            .O(N__33305),
            .I(N__33286));
    Sp12to4 I__8101 (
            .O(N__33302),
            .I(N__33286));
    Sp12to4 I__8100 (
            .O(N__33299),
            .I(N__33286));
    LocalMux I__8099 (
            .O(N__33296),
            .I(N__33283));
    Span12Mux_v I__8098 (
            .O(N__33293),
            .I(N__33280));
    Span12Mux_h I__8097 (
            .O(N__33286),
            .I(N__33277));
    Span4Mux_v I__8096 (
            .O(N__33283),
            .I(N__33274));
    Odrv12 I__8095 (
            .O(N__33280),
            .I(port_data_c_1));
    Odrv12 I__8094 (
            .O(N__33277),
            .I(port_data_c_1));
    Odrv4 I__8093 (
            .O(N__33274),
            .I(port_data_c_1));
    InMux I__8092 (
            .O(N__33267),
            .I(N__33264));
    LocalMux I__8091 (
            .O(N__33264),
            .I(this_vga_signals_M_this_external_address_q_3_i_0_0_15));
    CascadeMux I__8090 (
            .O(N__33261),
            .I(N__33258));
    InMux I__8089 (
            .O(N__33258),
            .I(N__33252));
    InMux I__8088 (
            .O(N__33257),
            .I(N__33252));
    LocalMux I__8087 (
            .O(N__33252),
            .I(N__33247));
    CascadeMux I__8086 (
            .O(N__33251),
            .I(N__33241));
    InMux I__8085 (
            .O(N__33250),
            .I(N__33236));
    Span4Mux_v I__8084 (
            .O(N__33247),
            .I(N__33233));
    InMux I__8083 (
            .O(N__33246),
            .I(N__33228));
    InMux I__8082 (
            .O(N__33245),
            .I(N__33228));
    InMux I__8081 (
            .O(N__33244),
            .I(N__33224));
    InMux I__8080 (
            .O(N__33241),
            .I(N__33219));
    InMux I__8079 (
            .O(N__33240),
            .I(N__33219));
    InMux I__8078 (
            .O(N__33239),
            .I(N__33216));
    LocalMux I__8077 (
            .O(N__33236),
            .I(N__33211));
    Span4Mux_v I__8076 (
            .O(N__33233),
            .I(N__33211));
    LocalMux I__8075 (
            .O(N__33228),
            .I(N__33208));
    InMux I__8074 (
            .O(N__33227),
            .I(N__33205));
    LocalMux I__8073 (
            .O(N__33224),
            .I(N__33202));
    LocalMux I__8072 (
            .O(N__33219),
            .I(N__33199));
    LocalMux I__8071 (
            .O(N__33216),
            .I(N__33196));
    Span4Mux_v I__8070 (
            .O(N__33211),
            .I(N__33193));
    Span12Mux_v I__8069 (
            .O(N__33208),
            .I(N__33190));
    LocalMux I__8068 (
            .O(N__33205),
            .I(N__33183));
    Span4Mux_v I__8067 (
            .O(N__33202),
            .I(N__33183));
    Span4Mux_v I__8066 (
            .O(N__33199),
            .I(N__33183));
    Odrv12 I__8065 (
            .O(N__33196),
            .I(N_661));
    Odrv4 I__8064 (
            .O(N__33193),
            .I(N_661));
    Odrv12 I__8063 (
            .O(N__33190),
            .I(N_661));
    Odrv4 I__8062 (
            .O(N__33183),
            .I(N_661));
    CEMux I__8061 (
            .O(N__33174),
            .I(N__33171));
    LocalMux I__8060 (
            .O(N__33171),
            .I(N__33167));
    CEMux I__8059 (
            .O(N__33170),
            .I(N__33164));
    Span4Mux_v I__8058 (
            .O(N__33167),
            .I(N__33161));
    LocalMux I__8057 (
            .O(N__33164),
            .I(N__33158));
    Odrv4 I__8056 (
            .O(N__33161),
            .I(\this_sprites_ram.mem_WE_2 ));
    Odrv4 I__8055 (
            .O(N__33158),
            .I(\this_sprites_ram.mem_WE_2 ));
    InMux I__8054 (
            .O(N__33153),
            .I(N__33150));
    LocalMux I__8053 (
            .O(N__33150),
            .I(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ));
    InMux I__8052 (
            .O(N__33147),
            .I(N__33144));
    LocalMux I__8051 (
            .O(N__33144),
            .I(N__33141));
    Odrv12 I__8050 (
            .O(N__33141),
            .I(M_this_oam_ram_read_data_i_9));
    InMux I__8049 (
            .O(N__33138),
            .I(\this_ppu.un2_hscroll_cry_0 ));
    CascadeMux I__8048 (
            .O(N__33135),
            .I(N__33132));
    InMux I__8047 (
            .O(N__33132),
            .I(N__33127));
    InMux I__8046 (
            .O(N__33131),
            .I(N__33124));
    CascadeMux I__8045 (
            .O(N__33130),
            .I(N__33121));
    LocalMux I__8044 (
            .O(N__33127),
            .I(N__33118));
    LocalMux I__8043 (
            .O(N__33124),
            .I(N__33115));
    InMux I__8042 (
            .O(N__33121),
            .I(N__33112));
    Span4Mux_h I__8041 (
            .O(N__33118),
            .I(N__33109));
    Span4Mux_v I__8040 (
            .O(N__33115),
            .I(N__33106));
    LocalMux I__8039 (
            .O(N__33112),
            .I(N__33103));
    Span4Mux_h I__8038 (
            .O(N__33109),
            .I(N__33100));
    Odrv4 I__8037 (
            .O(N__33106),
            .I(M_this_oam_ram_read_data_10));
    Odrv12 I__8036 (
            .O(N__33103),
            .I(M_this_oam_ram_read_data_10));
    Odrv4 I__8035 (
            .O(N__33100),
            .I(M_this_oam_ram_read_data_10));
    InMux I__8034 (
            .O(N__33093),
            .I(\this_ppu.un2_hscroll_cry_1 ));
    InMux I__8033 (
            .O(N__33090),
            .I(N__33087));
    LocalMux I__8032 (
            .O(N__33087),
            .I(N__33084));
    Span4Mux_v I__8031 (
            .O(N__33084),
            .I(N__33081));
    Odrv4 I__8030 (
            .O(N__33081),
            .I(M_this_oam_ram_write_data_26));
    InMux I__8029 (
            .O(N__33078),
            .I(N__33075));
    LocalMux I__8028 (
            .O(N__33075),
            .I(N__33072));
    Span4Mux_h I__8027 (
            .O(N__33072),
            .I(N__33069));
    Odrv4 I__8026 (
            .O(N__33069),
            .I(M_this_oam_ram_write_data_19));
    CascadeMux I__8025 (
            .O(N__33066),
            .I(N__33061));
    CascadeMux I__8024 (
            .O(N__33065),
            .I(N__33057));
    InMux I__8023 (
            .O(N__33064),
            .I(N__33054));
    InMux I__8022 (
            .O(N__33061),
            .I(N__33051));
    InMux I__8021 (
            .O(N__33060),
            .I(N__33048));
    InMux I__8020 (
            .O(N__33057),
            .I(N__33045));
    LocalMux I__8019 (
            .O(N__33054),
            .I(N__33040));
    LocalMux I__8018 (
            .O(N__33051),
            .I(N__33040));
    LocalMux I__8017 (
            .O(N__33048),
            .I(N__33036));
    LocalMux I__8016 (
            .O(N__33045),
            .I(N__33033));
    Span4Mux_v I__8015 (
            .O(N__33040),
            .I(N__33028));
    InMux I__8014 (
            .O(N__33039),
            .I(N__33025));
    Span4Mux_v I__8013 (
            .O(N__33036),
            .I(N__33022));
    Span12Mux_v I__8012 (
            .O(N__33033),
            .I(N__33019));
    InMux I__8011 (
            .O(N__33032),
            .I(N__33016));
    InMux I__8010 (
            .O(N__33031),
            .I(N__33013));
    Span4Mux_h I__8009 (
            .O(N__33028),
            .I(N__33010));
    LocalMux I__8008 (
            .O(N__33025),
            .I(N__33005));
    Span4Mux_v I__8007 (
            .O(N__33022),
            .I(N__33005));
    Odrv12 I__8006 (
            .O(N__33019),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__8005 (
            .O(N__33016),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__8004 (
            .O(N__33013),
            .I(M_this_ppu_vram_addr_1));
    Odrv4 I__8003 (
            .O(N__33010),
            .I(M_this_ppu_vram_addr_1));
    Odrv4 I__8002 (
            .O(N__33005),
            .I(M_this_ppu_vram_addr_1));
    InMux I__8001 (
            .O(N__32994),
            .I(N__32991));
    LocalMux I__8000 (
            .O(N__32991),
            .I(\this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ));
    CascadeMux I__7999 (
            .O(N__32988),
            .I(N__32985));
    InMux I__7998 (
            .O(N__32985),
            .I(N__32978));
    CascadeMux I__7997 (
            .O(N__32984),
            .I(N__32975));
    CascadeMux I__7996 (
            .O(N__32983),
            .I(N__32972));
    CascadeMux I__7995 (
            .O(N__32982),
            .I(N__32968));
    CascadeMux I__7994 (
            .O(N__32981),
            .I(N__32965));
    LocalMux I__7993 (
            .O(N__32978),
            .I(N__32960));
    InMux I__7992 (
            .O(N__32975),
            .I(N__32957));
    InMux I__7991 (
            .O(N__32972),
            .I(N__32954));
    CascadeMux I__7990 (
            .O(N__32971),
            .I(N__32951));
    InMux I__7989 (
            .O(N__32968),
            .I(N__32948));
    InMux I__7988 (
            .O(N__32965),
            .I(N__32945));
    CascadeMux I__7987 (
            .O(N__32964),
            .I(N__32942));
    CascadeMux I__7986 (
            .O(N__32963),
            .I(N__32939));
    Span4Mux_v I__7985 (
            .O(N__32960),
            .I(N__32930));
    LocalMux I__7984 (
            .O(N__32957),
            .I(N__32930));
    LocalMux I__7983 (
            .O(N__32954),
            .I(N__32930));
    InMux I__7982 (
            .O(N__32951),
            .I(N__32927));
    LocalMux I__7981 (
            .O(N__32948),
            .I(N__32922));
    LocalMux I__7980 (
            .O(N__32945),
            .I(N__32922));
    InMux I__7979 (
            .O(N__32942),
            .I(N__32919));
    InMux I__7978 (
            .O(N__32939),
            .I(N__32916));
    CascadeMux I__7977 (
            .O(N__32938),
            .I(N__32913));
    CascadeMux I__7976 (
            .O(N__32937),
            .I(N__32910));
    Span4Mux_v I__7975 (
            .O(N__32930),
            .I(N__32903));
    LocalMux I__7974 (
            .O(N__32927),
            .I(N__32903));
    Span4Mux_v I__7973 (
            .O(N__32922),
            .I(N__32900));
    LocalMux I__7972 (
            .O(N__32919),
            .I(N__32895));
    LocalMux I__7971 (
            .O(N__32916),
            .I(N__32895));
    InMux I__7970 (
            .O(N__32913),
            .I(N__32892));
    InMux I__7969 (
            .O(N__32910),
            .I(N__32889));
    CascadeMux I__7968 (
            .O(N__32909),
            .I(N__32886));
    CascadeMux I__7967 (
            .O(N__32908),
            .I(N__32883));
    Span4Mux_v I__7966 (
            .O(N__32903),
            .I(N__32879));
    Span4Mux_v I__7965 (
            .O(N__32900),
            .I(N__32869));
    Span4Mux_v I__7964 (
            .O(N__32895),
            .I(N__32869));
    LocalMux I__7963 (
            .O(N__32892),
            .I(N__32869));
    LocalMux I__7962 (
            .O(N__32889),
            .I(N__32869));
    InMux I__7961 (
            .O(N__32886),
            .I(N__32866));
    InMux I__7960 (
            .O(N__32883),
            .I(N__32863));
    CascadeMux I__7959 (
            .O(N__32882),
            .I(N__32860));
    Span4Mux_v I__7958 (
            .O(N__32879),
            .I(N__32857));
    CascadeMux I__7957 (
            .O(N__32878),
            .I(N__32854));
    Span4Mux_v I__7956 (
            .O(N__32869),
            .I(N__32847));
    LocalMux I__7955 (
            .O(N__32866),
            .I(N__32847));
    LocalMux I__7954 (
            .O(N__32863),
            .I(N__32847));
    InMux I__7953 (
            .O(N__32860),
            .I(N__32844));
    Sp12to4 I__7952 (
            .O(N__32857),
            .I(N__32839));
    InMux I__7951 (
            .O(N__32854),
            .I(N__32836));
    Span4Mux_v I__7950 (
            .O(N__32847),
            .I(N__32831));
    LocalMux I__7949 (
            .O(N__32844),
            .I(N__32831));
    CascadeMux I__7948 (
            .O(N__32843),
            .I(N__32828));
    CascadeMux I__7947 (
            .O(N__32842),
            .I(N__32825));
    Span12Mux_h I__7946 (
            .O(N__32839),
            .I(N__32822));
    LocalMux I__7945 (
            .O(N__32836),
            .I(N__32819));
    Span4Mux_v I__7944 (
            .O(N__32831),
            .I(N__32816));
    InMux I__7943 (
            .O(N__32828),
            .I(N__32813));
    InMux I__7942 (
            .O(N__32825),
            .I(N__32810));
    Odrv12 I__7941 (
            .O(N__32822),
            .I(M_this_ppu_sprites_addr_1));
    Odrv4 I__7940 (
            .O(N__32819),
            .I(M_this_ppu_sprites_addr_1));
    Odrv4 I__7939 (
            .O(N__32816),
            .I(M_this_ppu_sprites_addr_1));
    LocalMux I__7938 (
            .O(N__32813),
            .I(M_this_ppu_sprites_addr_1));
    LocalMux I__7937 (
            .O(N__32810),
            .I(M_this_ppu_sprites_addr_1));
    InMux I__7936 (
            .O(N__32799),
            .I(N__32795));
    InMux I__7935 (
            .O(N__32798),
            .I(N__32790));
    LocalMux I__7934 (
            .O(N__32795),
            .I(N__32787));
    InMux I__7933 (
            .O(N__32794),
            .I(N__32784));
    InMux I__7932 (
            .O(N__32793),
            .I(N__32781));
    LocalMux I__7931 (
            .O(N__32790),
            .I(N__32778));
    Span4Mux_h I__7930 (
            .O(N__32787),
            .I(N__32775));
    LocalMux I__7929 (
            .O(N__32784),
            .I(N__32770));
    LocalMux I__7928 (
            .O(N__32781),
            .I(N__32770));
    Span4Mux_h I__7927 (
            .O(N__32778),
            .I(N__32767));
    Span4Mux_h I__7926 (
            .O(N__32775),
            .I(N__32764));
    Span4Mux_v I__7925 (
            .O(N__32770),
            .I(N__32761));
    Odrv4 I__7924 (
            .O(N__32767),
            .I(M_this_oam_ram_read_data_8));
    Odrv4 I__7923 (
            .O(N__32764),
            .I(M_this_oam_ram_read_data_8));
    Odrv4 I__7922 (
            .O(N__32761),
            .I(M_this_oam_ram_read_data_8));
    CascadeMux I__7921 (
            .O(N__32754),
            .I(N__32751));
    InMux I__7920 (
            .O(N__32751),
            .I(N__32748));
    LocalMux I__7919 (
            .O(N__32748),
            .I(N__32744));
    CascadeMux I__7918 (
            .O(N__32747),
            .I(N__32740));
    Span4Mux_v I__7917 (
            .O(N__32744),
            .I(N__32734));
    InMux I__7916 (
            .O(N__32743),
            .I(N__32731));
    InMux I__7915 (
            .O(N__32740),
            .I(N__32728));
    InMux I__7914 (
            .O(N__32739),
            .I(N__32725));
    CascadeMux I__7913 (
            .O(N__32738),
            .I(N__32722));
    CascadeMux I__7912 (
            .O(N__32737),
            .I(N__32717));
    Span4Mux_h I__7911 (
            .O(N__32734),
            .I(N__32714));
    LocalMux I__7910 (
            .O(N__32731),
            .I(N__32711));
    LocalMux I__7909 (
            .O(N__32728),
            .I(N__32706));
    LocalMux I__7908 (
            .O(N__32725),
            .I(N__32706));
    InMux I__7907 (
            .O(N__32722),
            .I(N__32701));
    InMux I__7906 (
            .O(N__32721),
            .I(N__32701));
    InMux I__7905 (
            .O(N__32720),
            .I(N__32698));
    InMux I__7904 (
            .O(N__32717),
            .I(N__32695));
    Span4Mux_h I__7903 (
            .O(N__32714),
            .I(N__32692));
    Span4Mux_v I__7902 (
            .O(N__32711),
            .I(N__32689));
    Span12Mux_v I__7901 (
            .O(N__32706),
            .I(N__32686));
    LocalMux I__7900 (
            .O(N__32701),
            .I(N__32681));
    LocalMux I__7899 (
            .O(N__32698),
            .I(N__32681));
    LocalMux I__7898 (
            .O(N__32695),
            .I(M_this_ppu_vram_addr_2));
    Odrv4 I__7897 (
            .O(N__32692),
            .I(M_this_ppu_vram_addr_2));
    Odrv4 I__7896 (
            .O(N__32689),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__7895 (
            .O(N__32686),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__7894 (
            .O(N__32681),
            .I(M_this_ppu_vram_addr_2));
    InMux I__7893 (
            .O(N__32670),
            .I(N__32667));
    LocalMux I__7892 (
            .O(N__32667),
            .I(N__32664));
    Odrv4 I__7891 (
            .O(N__32664),
            .I(\this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ));
    CascadeMux I__7890 (
            .O(N__32661),
            .I(N__32657));
    CascadeMux I__7889 (
            .O(N__32660),
            .I(N__32654));
    InMux I__7888 (
            .O(N__32657),
            .I(N__32645));
    InMux I__7887 (
            .O(N__32654),
            .I(N__32642));
    CascadeMux I__7886 (
            .O(N__32653),
            .I(N__32639));
    CascadeMux I__7885 (
            .O(N__32652),
            .I(N__32636));
    CascadeMux I__7884 (
            .O(N__32651),
            .I(N__32631));
    CascadeMux I__7883 (
            .O(N__32650),
            .I(N__32628));
    CascadeMux I__7882 (
            .O(N__32649),
            .I(N__32625));
    CascadeMux I__7881 (
            .O(N__32648),
            .I(N__32622));
    LocalMux I__7880 (
            .O(N__32645),
            .I(N__32616));
    LocalMux I__7879 (
            .O(N__32642),
            .I(N__32616));
    InMux I__7878 (
            .O(N__32639),
            .I(N__32613));
    InMux I__7877 (
            .O(N__32636),
            .I(N__32610));
    CascadeMux I__7876 (
            .O(N__32635),
            .I(N__32607));
    CascadeMux I__7875 (
            .O(N__32634),
            .I(N__32604));
    InMux I__7874 (
            .O(N__32631),
            .I(N__32599));
    InMux I__7873 (
            .O(N__32628),
            .I(N__32596));
    InMux I__7872 (
            .O(N__32625),
            .I(N__32593));
    InMux I__7871 (
            .O(N__32622),
            .I(N__32590));
    CascadeMux I__7870 (
            .O(N__32621),
            .I(N__32587));
    Span4Mux_v I__7869 (
            .O(N__32616),
            .I(N__32580));
    LocalMux I__7868 (
            .O(N__32613),
            .I(N__32580));
    LocalMux I__7867 (
            .O(N__32610),
            .I(N__32580));
    InMux I__7866 (
            .O(N__32607),
            .I(N__32577));
    InMux I__7865 (
            .O(N__32604),
            .I(N__32574));
    CascadeMux I__7864 (
            .O(N__32603),
            .I(N__32571));
    CascadeMux I__7863 (
            .O(N__32602),
            .I(N__32568));
    LocalMux I__7862 (
            .O(N__32599),
            .I(N__32557));
    LocalMux I__7861 (
            .O(N__32596),
            .I(N__32557));
    LocalMux I__7860 (
            .O(N__32593),
            .I(N__32557));
    LocalMux I__7859 (
            .O(N__32590),
            .I(N__32557));
    InMux I__7858 (
            .O(N__32587),
            .I(N__32554));
    Span4Mux_v I__7857 (
            .O(N__32580),
            .I(N__32547));
    LocalMux I__7856 (
            .O(N__32577),
            .I(N__32547));
    LocalMux I__7855 (
            .O(N__32574),
            .I(N__32547));
    InMux I__7854 (
            .O(N__32571),
            .I(N__32544));
    InMux I__7853 (
            .O(N__32568),
            .I(N__32541));
    CascadeMux I__7852 (
            .O(N__32567),
            .I(N__32538));
    CascadeMux I__7851 (
            .O(N__32566),
            .I(N__32535));
    Span12Mux_v I__7850 (
            .O(N__32557),
            .I(N__32531));
    LocalMux I__7849 (
            .O(N__32554),
            .I(N__32528));
    Span4Mux_v I__7848 (
            .O(N__32547),
            .I(N__32521));
    LocalMux I__7847 (
            .O(N__32544),
            .I(N__32521));
    LocalMux I__7846 (
            .O(N__32541),
            .I(N__32521));
    InMux I__7845 (
            .O(N__32538),
            .I(N__32518));
    InMux I__7844 (
            .O(N__32535),
            .I(N__32515));
    CascadeMux I__7843 (
            .O(N__32534),
            .I(N__32512));
    Span12Mux_h I__7842 (
            .O(N__32531),
            .I(N__32509));
    Span4Mux_v I__7841 (
            .O(N__32528),
            .I(N__32502));
    Span4Mux_v I__7840 (
            .O(N__32521),
            .I(N__32502));
    LocalMux I__7839 (
            .O(N__32518),
            .I(N__32502));
    LocalMux I__7838 (
            .O(N__32515),
            .I(N__32499));
    InMux I__7837 (
            .O(N__32512),
            .I(N__32496));
    Odrv12 I__7836 (
            .O(N__32509),
            .I(M_this_ppu_sprites_addr_2));
    Odrv4 I__7835 (
            .O(N__32502),
            .I(M_this_ppu_sprites_addr_2));
    Odrv4 I__7834 (
            .O(N__32499),
            .I(M_this_ppu_sprites_addr_2));
    LocalMux I__7833 (
            .O(N__32496),
            .I(M_this_ppu_sprites_addr_2));
    InMux I__7832 (
            .O(N__32487),
            .I(N__32484));
    LocalMux I__7831 (
            .O(N__32484),
            .I(N__32481));
    Span4Mux_v I__7830 (
            .O(N__32481),
            .I(N__32478));
    Odrv4 I__7829 (
            .O(N__32478),
            .I(M_this_data_tmp_qZ0Z_22));
    InMux I__7828 (
            .O(N__32475),
            .I(N__32472));
    LocalMux I__7827 (
            .O(N__32472),
            .I(N__32469));
    Odrv4 I__7826 (
            .O(N__32469),
            .I(M_this_oam_ram_write_data_22));
    InMux I__7825 (
            .O(N__32466),
            .I(N__32463));
    LocalMux I__7824 (
            .O(N__32463),
            .I(M_this_oam_ram_write_data_31));
    InMux I__7823 (
            .O(N__32460),
            .I(N__32457));
    LocalMux I__7822 (
            .O(N__32457),
            .I(M_this_data_tmp_qZ0Z_18));
    InMux I__7821 (
            .O(N__32454),
            .I(N__32451));
    LocalMux I__7820 (
            .O(N__32451),
            .I(M_this_data_tmp_qZ0Z_20));
    InMux I__7819 (
            .O(N__32448),
            .I(N__32445));
    LocalMux I__7818 (
            .O(N__32445),
            .I(N__32438));
    InMux I__7817 (
            .O(N__32444),
            .I(N__32435));
    InMux I__7816 (
            .O(N__32443),
            .I(N__32430));
    InMux I__7815 (
            .O(N__32442),
            .I(N__32430));
    CascadeMux I__7814 (
            .O(N__32441),
            .I(N__32427));
    Span4Mux_v I__7813 (
            .O(N__32438),
            .I(N__32421));
    LocalMux I__7812 (
            .O(N__32435),
            .I(N__32421));
    LocalMux I__7811 (
            .O(N__32430),
            .I(N__32418));
    InMux I__7810 (
            .O(N__32427),
            .I(N__32414));
    CascadeMux I__7809 (
            .O(N__32426),
            .I(N__32410));
    Span4Mux_v I__7808 (
            .O(N__32421),
            .I(N__32407));
    Span4Mux_v I__7807 (
            .O(N__32418),
            .I(N__32402));
    InMux I__7806 (
            .O(N__32417),
            .I(N__32399));
    LocalMux I__7805 (
            .O(N__32414),
            .I(N__32396));
    CascadeMux I__7804 (
            .O(N__32413),
            .I(N__32393));
    InMux I__7803 (
            .O(N__32410),
            .I(N__32390));
    Span4Mux_v I__7802 (
            .O(N__32407),
            .I(N__32387));
    InMux I__7801 (
            .O(N__32406),
            .I(N__32384));
    CascadeMux I__7800 (
            .O(N__32405),
            .I(N__32380));
    Span4Mux_v I__7799 (
            .O(N__32402),
            .I(N__32377));
    LocalMux I__7798 (
            .O(N__32399),
            .I(N__32374));
    Span4Mux_v I__7797 (
            .O(N__32396),
            .I(N__32371));
    InMux I__7796 (
            .O(N__32393),
            .I(N__32368));
    LocalMux I__7795 (
            .O(N__32390),
            .I(N__32365));
    Span4Mux_v I__7794 (
            .O(N__32387),
            .I(N__32360));
    LocalMux I__7793 (
            .O(N__32384),
            .I(N__32360));
    InMux I__7792 (
            .O(N__32383),
            .I(N__32357));
    InMux I__7791 (
            .O(N__32380),
            .I(N__32354));
    Sp12to4 I__7790 (
            .O(N__32377),
            .I(N__32351));
    Span4Mux_v I__7789 (
            .O(N__32374),
            .I(N__32348));
    Span4Mux_h I__7788 (
            .O(N__32371),
            .I(N__32343));
    LocalMux I__7787 (
            .O(N__32368),
            .I(N__32343));
    Span4Mux_v I__7786 (
            .O(N__32365),
            .I(N__32340));
    Span4Mux_v I__7785 (
            .O(N__32360),
            .I(N__32337));
    LocalMux I__7784 (
            .O(N__32357),
            .I(N__32332));
    LocalMux I__7783 (
            .O(N__32354),
            .I(N__32332));
    Span12Mux_h I__7782 (
            .O(N__32351),
            .I(N__32329));
    Sp12to4 I__7781 (
            .O(N__32348),
            .I(N__32326));
    Sp12to4 I__7780 (
            .O(N__32343),
            .I(N__32323));
    Span4Mux_h I__7779 (
            .O(N__32340),
            .I(N__32318));
    Span4Mux_v I__7778 (
            .O(N__32337),
            .I(N__32318));
    Span4Mux_v I__7777 (
            .O(N__32332),
            .I(N__32315));
    Span12Mux_v I__7776 (
            .O(N__32329),
            .I(N__32312));
    Span12Mux_h I__7775 (
            .O(N__32326),
            .I(N__32303));
    Span12Mux_v I__7774 (
            .O(N__32323),
            .I(N__32303));
    Sp12to4 I__7773 (
            .O(N__32318),
            .I(N__32303));
    Sp12to4 I__7772 (
            .O(N__32315),
            .I(N__32303));
    Odrv12 I__7771 (
            .O(N__32312),
            .I(port_data_c_4));
    Odrv12 I__7770 (
            .O(N__32303),
            .I(port_data_c_4));
    InMux I__7769 (
            .O(N__32298),
            .I(N__32295));
    LocalMux I__7768 (
            .O(N__32295),
            .I(N__32292));
    Odrv4 I__7767 (
            .O(N__32292),
            .I(M_this_oam_ram_write_data_28));
    InMux I__7766 (
            .O(N__32289),
            .I(N__32286));
    LocalMux I__7765 (
            .O(N__32286),
            .I(N__32283));
    Odrv4 I__7764 (
            .O(N__32283),
            .I(M_this_data_tmp_qZ0Z_21));
    InMux I__7763 (
            .O(N__32280),
            .I(N__32277));
    LocalMux I__7762 (
            .O(N__32277),
            .I(M_this_oam_ram_write_data_21));
    CascadeMux I__7761 (
            .O(N__32274),
            .I(N__32271));
    CascadeBuf I__7760 (
            .O(N__32271),
            .I(N__32268));
    CascadeMux I__7759 (
            .O(N__32268),
            .I(N__32263));
    InMux I__7758 (
            .O(N__32267),
            .I(N__32258));
    InMux I__7757 (
            .O(N__32266),
            .I(N__32258));
    InMux I__7756 (
            .O(N__32263),
            .I(N__32255));
    LocalMux I__7755 (
            .O(N__32258),
            .I(M_this_oam_address_qZ0Z_6));
    LocalMux I__7754 (
            .O(N__32255),
            .I(M_this_oam_address_qZ0Z_6));
    InMux I__7753 (
            .O(N__32250),
            .I(N__32244));
    InMux I__7752 (
            .O(N__32249),
            .I(N__32244));
    LocalMux I__7751 (
            .O(N__32244),
            .I(un1_M_this_oam_address_q_c6));
    CascadeMux I__7750 (
            .O(N__32241),
            .I(N__32238));
    CascadeBuf I__7749 (
            .O(N__32238),
            .I(N__32234));
    CascadeMux I__7748 (
            .O(N__32237),
            .I(N__32231));
    CascadeMux I__7747 (
            .O(N__32234),
            .I(N__32228));
    InMux I__7746 (
            .O(N__32231),
            .I(N__32225));
    InMux I__7745 (
            .O(N__32228),
            .I(N__32222));
    LocalMux I__7744 (
            .O(N__32225),
            .I(M_this_oam_address_qZ0Z_7));
    LocalMux I__7743 (
            .O(N__32222),
            .I(M_this_oam_address_qZ0Z_7));
    SRMux I__7742 (
            .O(N__32217),
            .I(N__32172));
    SRMux I__7741 (
            .O(N__32216),
            .I(N__32172));
    SRMux I__7740 (
            .O(N__32215),
            .I(N__32172));
    SRMux I__7739 (
            .O(N__32214),
            .I(N__32172));
    SRMux I__7738 (
            .O(N__32213),
            .I(N__32172));
    SRMux I__7737 (
            .O(N__32212),
            .I(N__32172));
    SRMux I__7736 (
            .O(N__32211),
            .I(N__32172));
    SRMux I__7735 (
            .O(N__32210),
            .I(N__32172));
    SRMux I__7734 (
            .O(N__32209),
            .I(N__32172));
    SRMux I__7733 (
            .O(N__32208),
            .I(N__32172));
    SRMux I__7732 (
            .O(N__32207),
            .I(N__32172));
    SRMux I__7731 (
            .O(N__32206),
            .I(N__32172));
    SRMux I__7730 (
            .O(N__32205),
            .I(N__32172));
    SRMux I__7729 (
            .O(N__32204),
            .I(N__32172));
    SRMux I__7728 (
            .O(N__32203),
            .I(N__32172));
    GlobalMux I__7727 (
            .O(N__32172),
            .I(N__32169));
    gio2CtrlBuf I__7726 (
            .O(N__32169),
            .I(N_404_g));
    InMux I__7725 (
            .O(N__32166),
            .I(N__32163));
    LocalMux I__7724 (
            .O(N__32163),
            .I(N__32160));
    Odrv12 I__7723 (
            .O(N__32160),
            .I(M_this_data_tmp_qZ0Z_9));
    InMux I__7722 (
            .O(N__32157),
            .I(N__32154));
    LocalMux I__7721 (
            .O(N__32154),
            .I(N__32151));
    Odrv4 I__7720 (
            .O(N__32151),
            .I(M_this_data_tmp_qZ0Z_12));
    InMux I__7719 (
            .O(N__32148),
            .I(N__32145));
    LocalMux I__7718 (
            .O(N__32145),
            .I(M_this_oam_ram_write_data_12));
    CascadeMux I__7717 (
            .O(N__32142),
            .I(N__32139));
    InMux I__7716 (
            .O(N__32139),
            .I(N__32134));
    InMux I__7715 (
            .O(N__32138),
            .I(N__32129));
    InMux I__7714 (
            .O(N__32137),
            .I(N__32129));
    LocalMux I__7713 (
            .O(N__32134),
            .I(N__32125));
    LocalMux I__7712 (
            .O(N__32129),
            .I(N__32122));
    InMux I__7711 (
            .O(N__32128),
            .I(N__32119));
    Span12Mux_h I__7710 (
            .O(N__32125),
            .I(N__32116));
    Span4Mux_h I__7709 (
            .O(N__32122),
            .I(N__32113));
    LocalMux I__7708 (
            .O(N__32119),
            .I(N__32110));
    Odrv12 I__7707 (
            .O(N__32116),
            .I(M_this_oam_ram_read_data_21));
    Odrv4 I__7706 (
            .O(N__32113),
            .I(M_this_oam_ram_read_data_21));
    Odrv4 I__7705 (
            .O(N__32110),
            .I(M_this_oam_ram_read_data_21));
    InMux I__7704 (
            .O(N__32103),
            .I(N__32100));
    LocalMux I__7703 (
            .O(N__32100),
            .I(N__32094));
    InMux I__7702 (
            .O(N__32099),
            .I(N__32089));
    InMux I__7701 (
            .O(N__32098),
            .I(N__32089));
    InMux I__7700 (
            .O(N__32097),
            .I(N__32086));
    Span4Mux_v I__7699 (
            .O(N__32094),
            .I(N__32081));
    LocalMux I__7698 (
            .O(N__32089),
            .I(N__32081));
    LocalMux I__7697 (
            .O(N__32086),
            .I(N__32078));
    Span4Mux_h I__7696 (
            .O(N__32081),
            .I(N__32075));
    Odrv4 I__7695 (
            .O(N__32078),
            .I(M_this_oam_ram_read_data_20));
    Odrv4 I__7694 (
            .O(N__32075),
            .I(M_this_oam_ram_read_data_20));
    InMux I__7693 (
            .O(N__32070),
            .I(N__32067));
    LocalMux I__7692 (
            .O(N__32067),
            .I(N__32060));
    InMux I__7691 (
            .O(N__32066),
            .I(N__32057));
    InMux I__7690 (
            .O(N__32065),
            .I(N__32052));
    InMux I__7689 (
            .O(N__32064),
            .I(N__32052));
    InMux I__7688 (
            .O(N__32063),
            .I(N__32049));
    Span4Mux_v I__7687 (
            .O(N__32060),
            .I(N__32042));
    LocalMux I__7686 (
            .O(N__32057),
            .I(N__32042));
    LocalMux I__7685 (
            .O(N__32052),
            .I(N__32042));
    LocalMux I__7684 (
            .O(N__32049),
            .I(N__32039));
    Span4Mux_h I__7683 (
            .O(N__32042),
            .I(N__32036));
    Odrv4 I__7682 (
            .O(N__32039),
            .I(M_this_oam_ram_read_data_19));
    Odrv4 I__7681 (
            .O(N__32036),
            .I(M_this_oam_ram_read_data_19));
    InMux I__7680 (
            .O(N__32031),
            .I(N__32028));
    LocalMux I__7679 (
            .O(N__32028),
            .I(N__32025));
    Odrv4 I__7678 (
            .O(N__32025),
            .I(\this_ppu.un1_M_vaddress_q_3_5 ));
    InMux I__7677 (
            .O(N__32022),
            .I(N__32019));
    LocalMux I__7676 (
            .O(N__32019),
            .I(N__32016));
    Span4Mux_h I__7675 (
            .O(N__32016),
            .I(N__32013));
    Span4Mux_h I__7674 (
            .O(N__32013),
            .I(N__32010));
    Odrv4 I__7673 (
            .O(N__32010),
            .I(M_this_data_tmp_qZ0Z_5));
    InMux I__7672 (
            .O(N__32007),
            .I(N__32004));
    LocalMux I__7671 (
            .O(N__32004),
            .I(M_this_oam_ram_write_data_5));
    InMux I__7670 (
            .O(N__32001),
            .I(N__31997));
    CascadeMux I__7669 (
            .O(N__32000),
            .I(N__31994));
    LocalMux I__7668 (
            .O(N__31997),
            .I(N__31991));
    InMux I__7667 (
            .O(N__31994),
            .I(N__31988));
    Span4Mux_h I__7666 (
            .O(N__31991),
            .I(N__31985));
    LocalMux I__7665 (
            .O(N__31988),
            .I(N__31981));
    Span4Mux_h I__7664 (
            .O(N__31985),
            .I(N__31978));
    InMux I__7663 (
            .O(N__31984),
            .I(N__31975));
    Odrv12 I__7662 (
            .O(N__31981),
            .I(M_this_oam_ram_read_data_9));
    Odrv4 I__7661 (
            .O(N__31978),
            .I(M_this_oam_ram_read_data_9));
    LocalMux I__7660 (
            .O(N__31975),
            .I(M_this_oam_ram_read_data_9));
    InMux I__7659 (
            .O(N__31968),
            .I(N__31965));
    LocalMux I__7658 (
            .O(N__31965),
            .I(M_this_oam_ram_write_data_9));
    InMux I__7657 (
            .O(N__31962),
            .I(N__31959));
    LocalMux I__7656 (
            .O(N__31959),
            .I(M_this_oam_ram_write_data_18));
    InMux I__7655 (
            .O(N__31956),
            .I(N__31953));
    LocalMux I__7654 (
            .O(N__31953),
            .I(M_this_oam_ram_write_data_20));
    InMux I__7653 (
            .O(N__31950),
            .I(N__31947));
    LocalMux I__7652 (
            .O(N__31947),
            .I(M_this_oam_ram_write_data_29));
    InMux I__7651 (
            .O(N__31944),
            .I(N__31941));
    LocalMux I__7650 (
            .O(N__31941),
            .I(M_this_oam_ram_write_data_30));
    InMux I__7649 (
            .O(N__31938),
            .I(N__31935));
    LocalMux I__7648 (
            .O(N__31935),
            .I(N__31932));
    Odrv4 I__7647 (
            .O(N__31932),
            .I(M_this_external_address_q_3_0_12));
    CEMux I__7646 (
            .O(N__31929),
            .I(N__31926));
    LocalMux I__7645 (
            .O(N__31926),
            .I(N__31922));
    CEMux I__7644 (
            .O(N__31925),
            .I(N__31919));
    Span4Mux_h I__7643 (
            .O(N__31922),
            .I(N__31916));
    LocalMux I__7642 (
            .O(N__31919),
            .I(N__31913));
    Span4Mux_h I__7641 (
            .O(N__31916),
            .I(N__31910));
    Span4Mux_h I__7640 (
            .O(N__31913),
            .I(N__31907));
    Odrv4 I__7639 (
            .O(N__31910),
            .I(\this_sprites_ram.mem_WE_4 ));
    Odrv4 I__7638 (
            .O(N__31907),
            .I(\this_sprites_ram.mem_WE_4 ));
    InMux I__7637 (
            .O(N__31902),
            .I(N__31899));
    LocalMux I__7636 (
            .O(N__31899),
            .I(N__31896));
    Span4Mux_h I__7635 (
            .O(N__31896),
            .I(N__31893));
    Span4Mux_h I__7634 (
            .O(N__31893),
            .I(N__31890));
    Odrv4 I__7633 (
            .O(N__31890),
            .I(\this_ppu.un1_M_haddress_q_2_5 ));
    InMux I__7632 (
            .O(N__31887),
            .I(N__31884));
    LocalMux I__7631 (
            .O(N__31884),
            .I(M_this_oam_ram_write_data_13));
    InMux I__7630 (
            .O(N__31881),
            .I(N__31878));
    LocalMux I__7629 (
            .O(N__31878),
            .I(M_this_oam_ram_write_data_15));
    InMux I__7628 (
            .O(N__31875),
            .I(N__31872));
    LocalMux I__7627 (
            .O(N__31872),
            .I(N__31868));
    CascadeMux I__7626 (
            .O(N__31871),
            .I(N__31865));
    Span4Mux_h I__7625 (
            .O(N__31868),
            .I(N__31862));
    InMux I__7624 (
            .O(N__31865),
            .I(N__31859));
    Odrv4 I__7623 (
            .O(N__31862),
            .I(M_this_oam_ram_read_data_15));
    LocalMux I__7622 (
            .O(N__31859),
            .I(M_this_oam_ram_read_data_15));
    InMux I__7621 (
            .O(N__31854),
            .I(N__31851));
    LocalMux I__7620 (
            .O(N__31851),
            .I(N__31848));
    Span4Mux_h I__7619 (
            .O(N__31848),
            .I(N__31845));
    Span4Mux_h I__7618 (
            .O(N__31845),
            .I(N__31842));
    Odrv4 I__7617 (
            .O(N__31842),
            .I(\this_ppu.un1_M_haddress_q_2_7 ));
    InMux I__7616 (
            .O(N__31839),
            .I(N__31835));
    InMux I__7615 (
            .O(N__31838),
            .I(N__31832));
    LocalMux I__7614 (
            .O(N__31835),
            .I(N__31825));
    LocalMux I__7613 (
            .O(N__31832),
            .I(N__31825));
    InMux I__7612 (
            .O(N__31831),
            .I(N__31820));
    InMux I__7611 (
            .O(N__31830),
            .I(N__31820));
    Odrv12 I__7610 (
            .O(N__31825),
            .I(M_this_oam_ram_read_data_12));
    LocalMux I__7609 (
            .O(N__31820),
            .I(M_this_oam_ram_read_data_12));
    InMux I__7608 (
            .O(N__31815),
            .I(N__31812));
    LocalMux I__7607 (
            .O(N__31812),
            .I(N__31807));
    InMux I__7606 (
            .O(N__31811),
            .I(N__31804));
    InMux I__7605 (
            .O(N__31810),
            .I(N__31801));
    Span4Mux_h I__7604 (
            .O(N__31807),
            .I(N__31798));
    LocalMux I__7603 (
            .O(N__31804),
            .I(N__31791));
    LocalMux I__7602 (
            .O(N__31801),
            .I(N__31791));
    Span4Mux_h I__7601 (
            .O(N__31798),
            .I(N__31788));
    InMux I__7600 (
            .O(N__31797),
            .I(N__31783));
    InMux I__7599 (
            .O(N__31796),
            .I(N__31783));
    Odrv12 I__7598 (
            .O(N__31791),
            .I(M_this_oam_ram_read_data_11));
    Odrv4 I__7597 (
            .O(N__31788),
            .I(M_this_oam_ram_read_data_11));
    LocalMux I__7596 (
            .O(N__31783),
            .I(M_this_oam_ram_read_data_11));
    InMux I__7595 (
            .O(N__31776),
            .I(N__31773));
    LocalMux I__7594 (
            .O(N__31773),
            .I(\this_ppu.un1_oam_data_1_c2 ));
    InMux I__7593 (
            .O(N__31770),
            .I(N__31767));
    LocalMux I__7592 (
            .O(N__31767),
            .I(N__31764));
    Span4Mux_h I__7591 (
            .O(N__31764),
            .I(N__31759));
    InMux I__7590 (
            .O(N__31763),
            .I(N__31756));
    InMux I__7589 (
            .O(N__31762),
            .I(N__31753));
    Odrv4 I__7588 (
            .O(N__31759),
            .I(M_this_oam_ram_read_data_14));
    LocalMux I__7587 (
            .O(N__31756),
            .I(M_this_oam_ram_read_data_14));
    LocalMux I__7586 (
            .O(N__31753),
            .I(M_this_oam_ram_read_data_14));
    CascadeMux I__7585 (
            .O(N__31746),
            .I(\this_ppu.un1_oam_data_1_c2_cascade_ ));
    InMux I__7584 (
            .O(N__31743),
            .I(N__31740));
    LocalMux I__7583 (
            .O(N__31740),
            .I(N__31734));
    InMux I__7582 (
            .O(N__31739),
            .I(N__31727));
    InMux I__7581 (
            .O(N__31738),
            .I(N__31727));
    InMux I__7580 (
            .O(N__31737),
            .I(N__31727));
    Odrv12 I__7579 (
            .O(N__31734),
            .I(M_this_oam_ram_read_data_13));
    LocalMux I__7578 (
            .O(N__31727),
            .I(M_this_oam_ram_read_data_13));
    InMux I__7577 (
            .O(N__31722),
            .I(N__31719));
    LocalMux I__7576 (
            .O(N__31719),
            .I(N__31716));
    Span4Mux_h I__7575 (
            .O(N__31716),
            .I(N__31713));
    Span4Mux_h I__7574 (
            .O(N__31713),
            .I(N__31710));
    Odrv4 I__7573 (
            .O(N__31710),
            .I(\this_ppu.un1_M_haddress_q_2_6 ));
    InMux I__7572 (
            .O(N__31707),
            .I(N__31703));
    InMux I__7571 (
            .O(N__31706),
            .I(N__31699));
    LocalMux I__7570 (
            .O(N__31703),
            .I(N__31696));
    InMux I__7569 (
            .O(N__31702),
            .I(N__31693));
    LocalMux I__7568 (
            .O(N__31699),
            .I(N__31690));
    Span4Mux_v I__7567 (
            .O(N__31696),
            .I(N__31685));
    LocalMux I__7566 (
            .O(N__31693),
            .I(N__31685));
    Span4Mux_v I__7565 (
            .O(N__31690),
            .I(N__31680));
    Span4Mux_h I__7564 (
            .O(N__31685),
            .I(N__31680));
    Odrv4 I__7563 (
            .O(N__31680),
            .I(\this_vga_signals.N_746 ));
    InMux I__7562 (
            .O(N__31677),
            .I(N__31674));
    LocalMux I__7561 (
            .O(N__31674),
            .I(\this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12 ));
    InMux I__7560 (
            .O(N__31671),
            .I(N__31667));
    InMux I__7559 (
            .O(N__31670),
            .I(N__31664));
    LocalMux I__7558 (
            .O(N__31667),
            .I(N__31661));
    LocalMux I__7557 (
            .O(N__31664),
            .I(M_this_oam_address_q_0_i_o3_0_a2_5));
    Odrv4 I__7556 (
            .O(N__31661),
            .I(M_this_oam_address_q_0_i_o3_0_a2_5));
    CascadeMux I__7555 (
            .O(N__31656),
            .I(\this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12_cascade_ ));
    IoInMux I__7554 (
            .O(N__31653),
            .I(N__31650));
    LocalMux I__7553 (
            .O(N__31650),
            .I(N__31647));
    IoSpan4Mux I__7552 (
            .O(N__31647),
            .I(N__31643));
    InMux I__7551 (
            .O(N__31646),
            .I(N__31640));
    Span4Mux_s2_h I__7550 (
            .O(N__31643),
            .I(N__31635));
    LocalMux I__7549 (
            .O(N__31640),
            .I(N__31632));
    InMux I__7548 (
            .O(N__31639),
            .I(N__31629));
    InMux I__7547 (
            .O(N__31638),
            .I(N__31626));
    Sp12to4 I__7546 (
            .O(N__31635),
            .I(N__31621));
    Span4Mux_h I__7545 (
            .O(N__31632),
            .I(N__31618));
    LocalMux I__7544 (
            .O(N__31629),
            .I(N__31615));
    LocalMux I__7543 (
            .O(N__31626),
            .I(N__31612));
    InMux I__7542 (
            .O(N__31625),
            .I(N__31609));
    InMux I__7541 (
            .O(N__31624),
            .I(N__31606));
    Span12Mux_s11_h I__7540 (
            .O(N__31621),
            .I(N__31603));
    Span4Mux_v I__7539 (
            .O(N__31618),
            .I(N__31598));
    Span4Mux_h I__7538 (
            .O(N__31615),
            .I(N__31598));
    Span4Mux_v I__7537 (
            .O(N__31612),
            .I(N__31595));
    LocalMux I__7536 (
            .O(N__31609),
            .I(N__31590));
    LocalMux I__7535 (
            .O(N__31606),
            .I(N__31590));
    Span12Mux_v I__7534 (
            .O(N__31603),
            .I(N__31586));
    Span4Mux_h I__7533 (
            .O(N__31598),
            .I(N__31583));
    Span4Mux_h I__7532 (
            .O(N__31595),
            .I(N__31578));
    Span4Mux_v I__7531 (
            .O(N__31590),
            .I(N__31578));
    InMux I__7530 (
            .O(N__31589),
            .I(N__31575));
    Odrv12 I__7529 (
            .O(N__31586),
            .I(led_c_1));
    Odrv4 I__7528 (
            .O(N__31583),
            .I(led_c_1));
    Odrv4 I__7527 (
            .O(N__31578),
            .I(led_c_1));
    LocalMux I__7526 (
            .O(N__31575),
            .I(led_c_1));
    InMux I__7525 (
            .O(N__31566),
            .I(N__31563));
    LocalMux I__7524 (
            .O(N__31563),
            .I(N__31559));
    InMux I__7523 (
            .O(N__31562),
            .I(N__31556));
    Span4Mux_v I__7522 (
            .O(N__31559),
            .I(N__31550));
    LocalMux I__7521 (
            .O(N__31556),
            .I(N__31550));
    InMux I__7520 (
            .O(N__31555),
            .I(N__31547));
    Span4Mux_h I__7519 (
            .O(N__31550),
            .I(N__31544));
    LocalMux I__7518 (
            .O(N__31547),
            .I(M_this_substate_qZ0));
    Odrv4 I__7517 (
            .O(N__31544),
            .I(M_this_substate_qZ0));
    InMux I__7516 (
            .O(N__31539),
            .I(N__31535));
    InMux I__7515 (
            .O(N__31538),
            .I(N__31532));
    LocalMux I__7514 (
            .O(N__31535),
            .I(N__31528));
    LocalMux I__7513 (
            .O(N__31532),
            .I(N__31525));
    InMux I__7512 (
            .O(N__31531),
            .I(N__31522));
    Span4Mux_v I__7511 (
            .O(N__31528),
            .I(N__31519));
    Span4Mux_v I__7510 (
            .O(N__31525),
            .I(N__31516));
    LocalMux I__7509 (
            .O(N__31522),
            .I(N__31513));
    Odrv4 I__7508 (
            .O(N__31519),
            .I(\this_vga_signals.N_419_0 ));
    Odrv4 I__7507 (
            .O(N__31516),
            .I(\this_vga_signals.N_419_0 ));
    Odrv12 I__7506 (
            .O(N__31513),
            .I(\this_vga_signals.N_419_0 ));
    InMux I__7505 (
            .O(N__31506),
            .I(N__31503));
    LocalMux I__7504 (
            .O(N__31503),
            .I(N__31500));
    Span4Mux_h I__7503 (
            .O(N__31500),
            .I(N__31497));
    Odrv4 I__7502 (
            .O(N__31497),
            .I(M_this_data_count_q_cry_6_THRU_CO));
    InMux I__7501 (
            .O(N__31494),
            .I(N__31476));
    InMux I__7500 (
            .O(N__31493),
            .I(N__31465));
    InMux I__7499 (
            .O(N__31492),
            .I(N__31465));
    InMux I__7498 (
            .O(N__31491),
            .I(N__31465));
    InMux I__7497 (
            .O(N__31490),
            .I(N__31465));
    InMux I__7496 (
            .O(N__31489),
            .I(N__31465));
    InMux I__7495 (
            .O(N__31488),
            .I(N__31458));
    InMux I__7494 (
            .O(N__31487),
            .I(N__31458));
    InMux I__7493 (
            .O(N__31486),
            .I(N__31458));
    InMux I__7492 (
            .O(N__31485),
            .I(N__31451));
    InMux I__7491 (
            .O(N__31484),
            .I(N__31451));
    InMux I__7490 (
            .O(N__31483),
            .I(N__31451));
    InMux I__7489 (
            .O(N__31482),
            .I(N__31442));
    InMux I__7488 (
            .O(N__31481),
            .I(N__31442));
    InMux I__7487 (
            .O(N__31480),
            .I(N__31442));
    InMux I__7486 (
            .O(N__31479),
            .I(N__31442));
    LocalMux I__7485 (
            .O(N__31476),
            .I(N_716_i));
    LocalMux I__7484 (
            .O(N__31465),
            .I(N_716_i));
    LocalMux I__7483 (
            .O(N__31458),
            .I(N_716_i));
    LocalMux I__7482 (
            .O(N__31451),
            .I(N_716_i));
    LocalMux I__7481 (
            .O(N__31442),
            .I(N_716_i));
    CascadeMux I__7480 (
            .O(N__31431),
            .I(N__31428));
    InMux I__7479 (
            .O(N__31428),
            .I(N__31424));
    CascadeMux I__7478 (
            .O(N__31427),
            .I(N__31421));
    LocalMux I__7477 (
            .O(N__31424),
            .I(N__31417));
    InMux I__7476 (
            .O(N__31421),
            .I(N__31414));
    InMux I__7475 (
            .O(N__31420),
            .I(N__31411));
    Span4Mux_v I__7474 (
            .O(N__31417),
            .I(N__31406));
    LocalMux I__7473 (
            .O(N__31414),
            .I(N__31406));
    LocalMux I__7472 (
            .O(N__31411),
            .I(M_this_data_count_qZ0Z_7));
    Odrv4 I__7471 (
            .O(N__31406),
            .I(M_this_data_count_qZ0Z_7));
    CEMux I__7470 (
            .O(N__31401),
            .I(N__31397));
    CEMux I__7469 (
            .O(N__31400),
            .I(N__31394));
    LocalMux I__7468 (
            .O(N__31397),
            .I(N__31389));
    LocalMux I__7467 (
            .O(N__31394),
            .I(N__31386));
    CEMux I__7466 (
            .O(N__31393),
            .I(N__31383));
    CEMux I__7465 (
            .O(N__31392),
            .I(N__31380));
    Span4Mux_v I__7464 (
            .O(N__31389),
            .I(N__31377));
    Span4Mux_v I__7463 (
            .O(N__31386),
            .I(N__31374));
    LocalMux I__7462 (
            .O(N__31383),
            .I(N__31369));
    LocalMux I__7461 (
            .O(N__31380),
            .I(N__31369));
    Odrv4 I__7460 (
            .O(N__31377),
            .I(N_364));
    Odrv4 I__7459 (
            .O(N__31374),
            .I(N_364));
    Odrv4 I__7458 (
            .O(N__31369),
            .I(N_364));
    CascadeMux I__7457 (
            .O(N__31362),
            .I(N__31357));
    InMux I__7456 (
            .O(N__31361),
            .I(N__31352));
    CascadeMux I__7455 (
            .O(N__31360),
            .I(N__31347));
    InMux I__7454 (
            .O(N__31357),
            .I(N__31344));
    InMux I__7453 (
            .O(N__31356),
            .I(N__31341));
    CascadeMux I__7452 (
            .O(N__31355),
            .I(N__31338));
    LocalMux I__7451 (
            .O(N__31352),
            .I(N__31334));
    InMux I__7450 (
            .O(N__31351),
            .I(N__31331));
    InMux I__7449 (
            .O(N__31350),
            .I(N__31328));
    InMux I__7448 (
            .O(N__31347),
            .I(N__31325));
    LocalMux I__7447 (
            .O(N__31344),
            .I(N__31321));
    LocalMux I__7446 (
            .O(N__31341),
            .I(N__31318));
    InMux I__7445 (
            .O(N__31338),
            .I(N__31315));
    CascadeMux I__7444 (
            .O(N__31337),
            .I(N__31312));
    Span4Mux_v I__7443 (
            .O(N__31334),
            .I(N__31307));
    LocalMux I__7442 (
            .O(N__31331),
            .I(N__31307));
    LocalMux I__7441 (
            .O(N__31328),
            .I(N__31304));
    LocalMux I__7440 (
            .O(N__31325),
            .I(N__31300));
    InMux I__7439 (
            .O(N__31324),
            .I(N__31297));
    Span4Mux_v I__7438 (
            .O(N__31321),
            .I(N__31292));
    Span4Mux_v I__7437 (
            .O(N__31318),
            .I(N__31292));
    LocalMux I__7436 (
            .O(N__31315),
            .I(N__31289));
    InMux I__7435 (
            .O(N__31312),
            .I(N__31286));
    Span4Mux_v I__7434 (
            .O(N__31307),
            .I(N__31283));
    Span4Mux_v I__7433 (
            .O(N__31304),
            .I(N__31280));
    InMux I__7432 (
            .O(N__31303),
            .I(N__31277));
    Span4Mux_v I__7431 (
            .O(N__31300),
            .I(N__31274));
    LocalMux I__7430 (
            .O(N__31297),
            .I(N__31271));
    Span4Mux_h I__7429 (
            .O(N__31292),
            .I(N__31264));
    Span4Mux_v I__7428 (
            .O(N__31289),
            .I(N__31264));
    LocalMux I__7427 (
            .O(N__31286),
            .I(N__31264));
    Sp12to4 I__7426 (
            .O(N__31283),
            .I(N__31256));
    Sp12to4 I__7425 (
            .O(N__31280),
            .I(N__31256));
    LocalMux I__7424 (
            .O(N__31277),
            .I(N__31256));
    Span4Mux_v I__7423 (
            .O(N__31274),
            .I(N__31253));
    Span4Mux_v I__7422 (
            .O(N__31271),
            .I(N__31250));
    Span4Mux_h I__7421 (
            .O(N__31264),
            .I(N__31247));
    InMux I__7420 (
            .O(N__31263),
            .I(N__31244));
    Span12Mux_h I__7419 (
            .O(N__31256),
            .I(N__31241));
    Sp12to4 I__7418 (
            .O(N__31253),
            .I(N__31236));
    Sp12to4 I__7417 (
            .O(N__31250),
            .I(N__31236));
    Span4Mux_v I__7416 (
            .O(N__31247),
            .I(N__31231));
    LocalMux I__7415 (
            .O(N__31244),
            .I(N__31231));
    Span12Mux_v I__7414 (
            .O(N__31241),
            .I(N__31228));
    Span12Mux_h I__7413 (
            .O(N__31236),
            .I(N__31225));
    Span4Mux_v I__7412 (
            .O(N__31231),
            .I(N__31222));
    Odrv12 I__7411 (
            .O(N__31228),
            .I(port_data_c_0));
    Odrv12 I__7410 (
            .O(N__31225),
            .I(port_data_c_0));
    Odrv4 I__7409 (
            .O(N__31222),
            .I(port_data_c_0));
    CascadeMux I__7408 (
            .O(N__31215),
            .I(N__31210));
    InMux I__7407 (
            .O(N__31214),
            .I(N__31206));
    InMux I__7406 (
            .O(N__31213),
            .I(N__31202));
    InMux I__7405 (
            .O(N__31210),
            .I(N__31197));
    InMux I__7404 (
            .O(N__31209),
            .I(N__31197));
    LocalMux I__7403 (
            .O(N__31206),
            .I(N__31194));
    InMux I__7402 (
            .O(N__31205),
            .I(N__31191));
    LocalMux I__7401 (
            .O(N__31202),
            .I(N__31188));
    LocalMux I__7400 (
            .O(N__31197),
            .I(N__31185));
    Span4Mux_v I__7399 (
            .O(N__31194),
            .I(N__31179));
    LocalMux I__7398 (
            .O(N__31191),
            .I(N__31179));
    Span4Mux_v I__7397 (
            .O(N__31188),
            .I(N__31173));
    Span4Mux_v I__7396 (
            .O(N__31185),
            .I(N__31173));
    InMux I__7395 (
            .O(N__31184),
            .I(N__31170));
    Span4Mux_h I__7394 (
            .O(N__31179),
            .I(N__31167));
    InMux I__7393 (
            .O(N__31178),
            .I(N__31164));
    Sp12to4 I__7392 (
            .O(N__31173),
            .I(N__31159));
    LocalMux I__7391 (
            .O(N__31170),
            .I(N__31159));
    Span4Mux_v I__7390 (
            .O(N__31167),
            .I(N__31156));
    LocalMux I__7389 (
            .O(N__31164),
            .I(M_this_state_qZ0Z_4));
    Odrv12 I__7388 (
            .O(N__31159),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__7387 (
            .O(N__31156),
            .I(M_this_state_qZ0Z_4));
    InMux I__7386 (
            .O(N__31149),
            .I(N__31137));
    InMux I__7385 (
            .O(N__31148),
            .I(N__31137));
    InMux I__7384 (
            .O(N__31147),
            .I(N__31134));
    InMux I__7383 (
            .O(N__31146),
            .I(N__31131));
    CascadeMux I__7382 (
            .O(N__31145),
            .I(N__31128));
    InMux I__7381 (
            .O(N__31144),
            .I(N__31112));
    CascadeMux I__7380 (
            .O(N__31143),
            .I(N__31108));
    CascadeMux I__7379 (
            .O(N__31142),
            .I(N__31098));
    LocalMux I__7378 (
            .O(N__31137),
            .I(N__31090));
    LocalMux I__7377 (
            .O(N__31134),
            .I(N__31090));
    LocalMux I__7376 (
            .O(N__31131),
            .I(N__31090));
    InMux I__7375 (
            .O(N__31128),
            .I(N__31085));
    InMux I__7374 (
            .O(N__31127),
            .I(N__31085));
    InMux I__7373 (
            .O(N__31126),
            .I(N__31077));
    InMux I__7372 (
            .O(N__31125),
            .I(N__31077));
    InMux I__7371 (
            .O(N__31124),
            .I(N__31073));
    InMux I__7370 (
            .O(N__31123),
            .I(N__31068));
    InMux I__7369 (
            .O(N__31122),
            .I(N__31068));
    InMux I__7368 (
            .O(N__31121),
            .I(N__31063));
    InMux I__7367 (
            .O(N__31120),
            .I(N__31063));
    InMux I__7366 (
            .O(N__31119),
            .I(N__31060));
    InMux I__7365 (
            .O(N__31118),
            .I(N__31057));
    InMux I__7364 (
            .O(N__31117),
            .I(N__31054));
    InMux I__7363 (
            .O(N__31116),
            .I(N__31049));
    InMux I__7362 (
            .O(N__31115),
            .I(N__31049));
    LocalMux I__7361 (
            .O(N__31112),
            .I(N__31046));
    InMux I__7360 (
            .O(N__31111),
            .I(N__31041));
    InMux I__7359 (
            .O(N__31108),
            .I(N__31041));
    InMux I__7358 (
            .O(N__31107),
            .I(N__31038));
    InMux I__7357 (
            .O(N__31106),
            .I(N__31035));
    InMux I__7356 (
            .O(N__31105),
            .I(N__31030));
    InMux I__7355 (
            .O(N__31104),
            .I(N__31030));
    InMux I__7354 (
            .O(N__31103),
            .I(N__31027));
    InMux I__7353 (
            .O(N__31102),
            .I(N__31024));
    InMux I__7352 (
            .O(N__31101),
            .I(N__31017));
    InMux I__7351 (
            .O(N__31098),
            .I(N__31017));
    InMux I__7350 (
            .O(N__31097),
            .I(N__31017));
    Span4Mux_v I__7349 (
            .O(N__31090),
            .I(N__31014));
    LocalMux I__7348 (
            .O(N__31085),
            .I(N__31011));
    InMux I__7347 (
            .O(N__31084),
            .I(N__31004));
    InMux I__7346 (
            .O(N__31083),
            .I(N__31004));
    InMux I__7345 (
            .O(N__31082),
            .I(N__31004));
    LocalMux I__7344 (
            .O(N__31077),
            .I(N__30997));
    InMux I__7343 (
            .O(N__31076),
            .I(N__30994));
    LocalMux I__7342 (
            .O(N__31073),
            .I(N__30987));
    LocalMux I__7341 (
            .O(N__31068),
            .I(N__30987));
    LocalMux I__7340 (
            .O(N__31063),
            .I(N__30987));
    LocalMux I__7339 (
            .O(N__31060),
            .I(N__30982));
    LocalMux I__7338 (
            .O(N__31057),
            .I(N__30982));
    LocalMux I__7337 (
            .O(N__31054),
            .I(N__30973));
    LocalMux I__7336 (
            .O(N__31049),
            .I(N__30973));
    Span4Mux_v I__7335 (
            .O(N__31046),
            .I(N__30973));
    LocalMux I__7334 (
            .O(N__31041),
            .I(N__30973));
    LocalMux I__7333 (
            .O(N__31038),
            .I(N__30970));
    LocalMux I__7332 (
            .O(N__31035),
            .I(N__30967));
    LocalMux I__7331 (
            .O(N__31030),
            .I(N__30963));
    LocalMux I__7330 (
            .O(N__31027),
            .I(N__30960));
    LocalMux I__7329 (
            .O(N__31024),
            .I(N__30949));
    LocalMux I__7328 (
            .O(N__31017),
            .I(N__30949));
    Span4Mux_h I__7327 (
            .O(N__31014),
            .I(N__30949));
    Span4Mux_h I__7326 (
            .O(N__31011),
            .I(N__30949));
    LocalMux I__7325 (
            .O(N__31004),
            .I(N__30949));
    InMux I__7324 (
            .O(N__31003),
            .I(N__30940));
    InMux I__7323 (
            .O(N__31002),
            .I(N__30935));
    InMux I__7322 (
            .O(N__31001),
            .I(N__30935));
    InMux I__7321 (
            .O(N__31000),
            .I(N__30932));
    Span4Mux_h I__7320 (
            .O(N__30997),
            .I(N__30923));
    LocalMux I__7319 (
            .O(N__30994),
            .I(N__30923));
    Span4Mux_v I__7318 (
            .O(N__30987),
            .I(N__30923));
    Span4Mux_v I__7317 (
            .O(N__30982),
            .I(N__30923));
    Span4Mux_h I__7316 (
            .O(N__30973),
            .I(N__30918));
    Span4Mux_h I__7315 (
            .O(N__30970),
            .I(N__30918));
    Span4Mux_h I__7314 (
            .O(N__30967),
            .I(N__30915));
    InMux I__7313 (
            .O(N__30966),
            .I(N__30912));
    Span4Mux_v I__7312 (
            .O(N__30963),
            .I(N__30905));
    Span4Mux_h I__7311 (
            .O(N__30960),
            .I(N__30905));
    Span4Mux_v I__7310 (
            .O(N__30949),
            .I(N__30905));
    InMux I__7309 (
            .O(N__30948),
            .I(N__30898));
    InMux I__7308 (
            .O(N__30947),
            .I(N__30898));
    InMux I__7307 (
            .O(N__30946),
            .I(N__30898));
    InMux I__7306 (
            .O(N__30945),
            .I(N__30891));
    InMux I__7305 (
            .O(N__30944),
            .I(N__30891));
    InMux I__7304 (
            .O(N__30943),
            .I(N__30891));
    LocalMux I__7303 (
            .O(N__30940),
            .I(N_888_0));
    LocalMux I__7302 (
            .O(N__30935),
            .I(N_888_0));
    LocalMux I__7301 (
            .O(N__30932),
            .I(N_888_0));
    Odrv4 I__7300 (
            .O(N__30923),
            .I(N_888_0));
    Odrv4 I__7299 (
            .O(N__30918),
            .I(N_888_0));
    Odrv4 I__7298 (
            .O(N__30915),
            .I(N_888_0));
    LocalMux I__7297 (
            .O(N__30912),
            .I(N_888_0));
    Odrv4 I__7296 (
            .O(N__30905),
            .I(N_888_0));
    LocalMux I__7295 (
            .O(N__30898),
            .I(N_888_0));
    LocalMux I__7294 (
            .O(N__30891),
            .I(N_888_0));
    CascadeMux I__7293 (
            .O(N__30870),
            .I(N_760_cascade_));
    InMux I__7292 (
            .O(N__30867),
            .I(N__30864));
    LocalMux I__7291 (
            .O(N__30864),
            .I(N__30861));
    Span4Mux_v I__7290 (
            .O(N__30861),
            .I(N__30858));
    Odrv4 I__7289 (
            .O(N__30858),
            .I(M_this_data_tmp_qZ0Z_8));
    CascadeMux I__7288 (
            .O(N__30855),
            .I(N__30849));
    CascadeMux I__7287 (
            .O(N__30854),
            .I(N__30846));
    CascadeMux I__7286 (
            .O(N__30853),
            .I(N__30841));
    CascadeMux I__7285 (
            .O(N__30852),
            .I(N__30838));
    InMux I__7284 (
            .O(N__30849),
            .I(N__30835));
    InMux I__7283 (
            .O(N__30846),
            .I(N__30832));
    CascadeMux I__7282 (
            .O(N__30845),
            .I(N__30829));
    InMux I__7281 (
            .O(N__30844),
            .I(N__30826));
    InMux I__7280 (
            .O(N__30841),
            .I(N__30823));
    InMux I__7279 (
            .O(N__30838),
            .I(N__30820));
    LocalMux I__7278 (
            .O(N__30835),
            .I(N__30815));
    LocalMux I__7277 (
            .O(N__30832),
            .I(N__30815));
    InMux I__7276 (
            .O(N__30829),
            .I(N__30812));
    LocalMux I__7275 (
            .O(N__30826),
            .I(N__30808));
    LocalMux I__7274 (
            .O(N__30823),
            .I(N__30805));
    LocalMux I__7273 (
            .O(N__30820),
            .I(N__30802));
    Span4Mux_v I__7272 (
            .O(N__30815),
            .I(N__30797));
    LocalMux I__7271 (
            .O(N__30812),
            .I(N__30797));
    InMux I__7270 (
            .O(N__30811),
            .I(N__30794));
    Span4Mux_v I__7269 (
            .O(N__30808),
            .I(N__30787));
    Span4Mux_v I__7268 (
            .O(N__30805),
            .I(N__30787));
    Span4Mux_h I__7267 (
            .O(N__30802),
            .I(N__30787));
    Sp12to4 I__7266 (
            .O(N__30797),
            .I(N__30782));
    LocalMux I__7265 (
            .O(N__30794),
            .I(N__30782));
    Span4Mux_v I__7264 (
            .O(N__30787),
            .I(N__30779));
    Span12Mux_v I__7263 (
            .O(N__30782),
            .I(N__30776));
    Odrv4 I__7262 (
            .O(N__30779),
            .I(N_413_0));
    Odrv12 I__7261 (
            .O(N__30776),
            .I(N_413_0));
    InMux I__7260 (
            .O(N__30771),
            .I(N__30765));
    InMux I__7259 (
            .O(N__30770),
            .I(N__30765));
    LocalMux I__7258 (
            .O(N__30765),
            .I(N__30761));
    InMux I__7257 (
            .O(N__30764),
            .I(N__30758));
    Span4Mux_v I__7256 (
            .O(N__30761),
            .I(N__30755));
    LocalMux I__7255 (
            .O(N__30758),
            .I(N__30752));
    Odrv4 I__7254 (
            .O(N__30755),
            .I(un1_M_this_oam_address_q_c4));
    Odrv12 I__7253 (
            .O(N__30752),
            .I(un1_M_this_oam_address_q_c4));
    CascadeMux I__7252 (
            .O(N__30747),
            .I(N__30744));
    CascadeBuf I__7251 (
            .O(N__30744),
            .I(N__30741));
    CascadeMux I__7250 (
            .O(N__30741),
            .I(N__30738));
    InMux I__7249 (
            .O(N__30738),
            .I(N__30735));
    LocalMux I__7248 (
            .O(N__30735),
            .I(N__30732));
    Span4Mux_h I__7247 (
            .O(N__30732),
            .I(N__30729));
    Span4Mux_v I__7246 (
            .O(N__30729),
            .I(N__30724));
    InMux I__7245 (
            .O(N__30728),
            .I(N__30721));
    InMux I__7244 (
            .O(N__30727),
            .I(N__30718));
    Span4Mux_h I__7243 (
            .O(N__30724),
            .I(N__30715));
    LocalMux I__7242 (
            .O(N__30721),
            .I(M_this_oam_address_qZ0Z_3));
    LocalMux I__7241 (
            .O(N__30718),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv4 I__7240 (
            .O(N__30715),
            .I(M_this_oam_address_qZ0Z_3));
    CascadeMux I__7239 (
            .O(N__30708),
            .I(N__30705));
    CascadeBuf I__7238 (
            .O(N__30705),
            .I(N__30702));
    CascadeMux I__7237 (
            .O(N__30702),
            .I(N__30699));
    InMux I__7236 (
            .O(N__30699),
            .I(N__30696));
    LocalMux I__7235 (
            .O(N__30696),
            .I(N__30693));
    Span4Mux_h I__7234 (
            .O(N__30693),
            .I(N__30687));
    InMux I__7233 (
            .O(N__30692),
            .I(N__30682));
    InMux I__7232 (
            .O(N__30691),
            .I(N__30682));
    InMux I__7231 (
            .O(N__30690),
            .I(N__30679));
    Span4Mux_v I__7230 (
            .O(N__30687),
            .I(N__30676));
    LocalMux I__7229 (
            .O(N__30682),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__7228 (
            .O(N__30679),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv4 I__7227 (
            .O(N__30676),
            .I(M_this_oam_address_qZ0Z_2));
    InMux I__7226 (
            .O(N__30669),
            .I(N__30662));
    InMux I__7225 (
            .O(N__30668),
            .I(N__30659));
    InMux I__7224 (
            .O(N__30667),
            .I(N__30655));
    InMux I__7223 (
            .O(N__30666),
            .I(N__30652));
    InMux I__7222 (
            .O(N__30665),
            .I(N__30649));
    LocalMux I__7221 (
            .O(N__30662),
            .I(N__30645));
    LocalMux I__7220 (
            .O(N__30659),
            .I(N__30642));
    InMux I__7219 (
            .O(N__30658),
            .I(N__30639));
    LocalMux I__7218 (
            .O(N__30655),
            .I(N__30636));
    LocalMux I__7217 (
            .O(N__30652),
            .I(N__30631));
    LocalMux I__7216 (
            .O(N__30649),
            .I(N__30631));
    InMux I__7215 (
            .O(N__30648),
            .I(N__30628));
    Span4Mux_h I__7214 (
            .O(N__30645),
            .I(N__30625));
    Span4Mux_h I__7213 (
            .O(N__30642),
            .I(N__30620));
    LocalMux I__7212 (
            .O(N__30639),
            .I(N__30620));
    Span4Mux_h I__7211 (
            .O(N__30636),
            .I(N__30615));
    Span4Mux_h I__7210 (
            .O(N__30631),
            .I(N__30615));
    LocalMux I__7209 (
            .O(N__30628),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__7208 (
            .O(N__30625),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__7207 (
            .O(N__30620),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__7206 (
            .O(N__30615),
            .I(M_this_oam_address_qZ0Z_0));
    InMux I__7205 (
            .O(N__30606),
            .I(N__30601));
    CascadeMux I__7204 (
            .O(N__30605),
            .I(N__30598));
    InMux I__7203 (
            .O(N__30604),
            .I(N__30594));
    LocalMux I__7202 (
            .O(N__30601),
            .I(N__30590));
    InMux I__7201 (
            .O(N__30598),
            .I(N__30587));
    InMux I__7200 (
            .O(N__30597),
            .I(N__30583));
    LocalMux I__7199 (
            .O(N__30594),
            .I(N__30580));
    InMux I__7198 (
            .O(N__30593),
            .I(N__30577));
    Span4Mux_h I__7197 (
            .O(N__30590),
            .I(N__30572));
    LocalMux I__7196 (
            .O(N__30587),
            .I(N__30572));
    InMux I__7195 (
            .O(N__30586),
            .I(N__30569));
    LocalMux I__7194 (
            .O(N__30583),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__7193 (
            .O(N__30580),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__7192 (
            .O(N__30577),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__7191 (
            .O(N__30572),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__7190 (
            .O(N__30569),
            .I(M_this_state_qZ0Z_13));
    InMux I__7189 (
            .O(N__30558),
            .I(N__30553));
    InMux I__7188 (
            .O(N__30557),
            .I(N__30549));
    InMux I__7187 (
            .O(N__30556),
            .I(N__30544));
    LocalMux I__7186 (
            .O(N__30553),
            .I(N__30541));
    InMux I__7185 (
            .O(N__30552),
            .I(N__30538));
    LocalMux I__7184 (
            .O(N__30549),
            .I(N__30535));
    CascadeMux I__7183 (
            .O(N__30548),
            .I(N__30532));
    InMux I__7182 (
            .O(N__30547),
            .I(N__30529));
    LocalMux I__7181 (
            .O(N__30544),
            .I(N__30526));
    Span4Mux_v I__7180 (
            .O(N__30541),
            .I(N__30519));
    LocalMux I__7179 (
            .O(N__30538),
            .I(N__30519));
    Span4Mux_h I__7178 (
            .O(N__30535),
            .I(N__30519));
    InMux I__7177 (
            .O(N__30532),
            .I(N__30516));
    LocalMux I__7176 (
            .O(N__30529),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv12 I__7175 (
            .O(N__30526),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__7174 (
            .O(N__30519),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__7173 (
            .O(N__30516),
            .I(M_this_oam_address_qZ0Z_1));
    InMux I__7172 (
            .O(N__30507),
            .I(N__30500));
    InMux I__7171 (
            .O(N__30506),
            .I(N__30500));
    InMux I__7170 (
            .O(N__30505),
            .I(N__30497));
    LocalMux I__7169 (
            .O(N__30500),
            .I(N__30492));
    LocalMux I__7168 (
            .O(N__30497),
            .I(N__30492));
    Odrv4 I__7167 (
            .O(N__30492),
            .I(un1_M_this_oam_address_q_c2));
    InMux I__7166 (
            .O(N__30489),
            .I(N__30485));
    InMux I__7165 (
            .O(N__30488),
            .I(N__30482));
    LocalMux I__7164 (
            .O(N__30485),
            .I(N__30477));
    LocalMux I__7163 (
            .O(N__30482),
            .I(N__30474));
    InMux I__7162 (
            .O(N__30481),
            .I(N__30471));
    InMux I__7161 (
            .O(N__30480),
            .I(N__30468));
    Odrv4 I__7160 (
            .O(N__30477),
            .I(\this_vga_signals.N_461_0 ));
    Odrv4 I__7159 (
            .O(N__30474),
            .I(\this_vga_signals.N_461_0 ));
    LocalMux I__7158 (
            .O(N__30471),
            .I(\this_vga_signals.N_461_0 ));
    LocalMux I__7157 (
            .O(N__30468),
            .I(\this_vga_signals.N_461_0 ));
    CascadeMux I__7156 (
            .O(N__30459),
            .I(N__30456));
    InMux I__7155 (
            .O(N__30456),
            .I(N__30453));
    LocalMux I__7154 (
            .O(N__30453),
            .I(N__30450));
    Span4Mux_h I__7153 (
            .O(N__30450),
            .I(N__30447));
    Odrv4 I__7152 (
            .O(N__30447),
            .I(\this_vga_signals.N_747 ));
    InMux I__7151 (
            .O(N__30444),
            .I(N__30439));
    InMux I__7150 (
            .O(N__30443),
            .I(N__30435));
    CascadeMux I__7149 (
            .O(N__30442),
            .I(N__30432));
    LocalMux I__7148 (
            .O(N__30439),
            .I(N__30428));
    InMux I__7147 (
            .O(N__30438),
            .I(N__30425));
    LocalMux I__7146 (
            .O(N__30435),
            .I(N__30422));
    InMux I__7145 (
            .O(N__30432),
            .I(N__30417));
    InMux I__7144 (
            .O(N__30431),
            .I(N__30417));
    Span4Mux_v I__7143 (
            .O(N__30428),
            .I(N__30411));
    LocalMux I__7142 (
            .O(N__30425),
            .I(N__30411));
    Span4Mux_v I__7141 (
            .O(N__30422),
            .I(N__30408));
    LocalMux I__7140 (
            .O(N__30417),
            .I(N__30405));
    CascadeMux I__7139 (
            .O(N__30416),
            .I(N__30401));
    Span4Mux_h I__7138 (
            .O(N__30411),
            .I(N__30398));
    Span4Mux_h I__7137 (
            .O(N__30408),
            .I(N__30393));
    Span4Mux_v I__7136 (
            .O(N__30405),
            .I(N__30393));
    InMux I__7135 (
            .O(N__30404),
            .I(N__30390));
    InMux I__7134 (
            .O(N__30401),
            .I(N__30387));
    Odrv4 I__7133 (
            .O(N__30398),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__7132 (
            .O(N__30393),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__7131 (
            .O(N__30390),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__7130 (
            .O(N__30387),
            .I(M_this_state_qZ0Z_9));
    InMux I__7129 (
            .O(N__30378),
            .I(N__30371));
    InMux I__7128 (
            .O(N__30377),
            .I(N__30368));
    InMux I__7127 (
            .O(N__30376),
            .I(N__30365));
    InMux I__7126 (
            .O(N__30375),
            .I(N__30362));
    InMux I__7125 (
            .O(N__30374),
            .I(N__30358));
    LocalMux I__7124 (
            .O(N__30371),
            .I(N__30355));
    LocalMux I__7123 (
            .O(N__30368),
            .I(N__30352));
    LocalMux I__7122 (
            .O(N__30365),
            .I(N__30347));
    LocalMux I__7121 (
            .O(N__30362),
            .I(N__30347));
    InMux I__7120 (
            .O(N__30361),
            .I(N__30344));
    LocalMux I__7119 (
            .O(N__30358),
            .I(N__30339));
    Span4Mux_v I__7118 (
            .O(N__30355),
            .I(N__30339));
    Span4Mux_v I__7117 (
            .O(N__30352),
            .I(N__30332));
    Span4Mux_v I__7116 (
            .O(N__30347),
            .I(N__30332));
    LocalMux I__7115 (
            .O(N__30344),
            .I(N__30332));
    Odrv4 I__7114 (
            .O(N__30339),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__7113 (
            .O(N__30332),
            .I(M_this_state_qZ0Z_7));
    InMux I__7112 (
            .O(N__30327),
            .I(N__30324));
    LocalMux I__7111 (
            .O(N__30324),
            .I(N__30320));
    InMux I__7110 (
            .O(N__30323),
            .I(N__30317));
    Odrv4 I__7109 (
            .O(N__30320),
            .I(\this_vga_signals.N_433_0 ));
    LocalMux I__7108 (
            .O(N__30317),
            .I(\this_vga_signals.N_433_0 ));
    InMux I__7107 (
            .O(N__30312),
            .I(N__30309));
    LocalMux I__7106 (
            .O(N__30309),
            .I(N__30306));
    Span4Mux_v I__7105 (
            .O(N__30306),
            .I(N__30303));
    Odrv4 I__7104 (
            .O(N__30303),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_i_1Z0Z_0 ));
    CascadeMux I__7103 (
            .O(N__30300),
            .I(N__30297));
    InMux I__7102 (
            .O(N__30297),
            .I(N__30294));
    LocalMux I__7101 (
            .O(N__30294),
            .I(N__30291));
    Span4Mux_v I__7100 (
            .O(N__30291),
            .I(N__30288));
    Odrv4 I__7099 (
            .O(N__30288),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_i_a4_4Z0Z_0 ));
    InMux I__7098 (
            .O(N__30285),
            .I(N__30281));
    InMux I__7097 (
            .O(N__30284),
            .I(N__30276));
    LocalMux I__7096 (
            .O(N__30281),
            .I(N__30273));
    InMux I__7095 (
            .O(N__30280),
            .I(N__30270));
    InMux I__7094 (
            .O(N__30279),
            .I(N__30267));
    LocalMux I__7093 (
            .O(N__30276),
            .I(N__30264));
    Span4Mux_h I__7092 (
            .O(N__30273),
            .I(N__30261));
    LocalMux I__7091 (
            .O(N__30270),
            .I(N__30256));
    LocalMux I__7090 (
            .O(N__30267),
            .I(N__30256));
    Odrv4 I__7089 (
            .O(N__30264),
            .I(M_this_state_d62));
    Odrv4 I__7088 (
            .O(N__30261),
            .I(M_this_state_d62));
    Odrv4 I__7087 (
            .O(N__30256),
            .I(M_this_state_d62));
    InMux I__7086 (
            .O(N__30249),
            .I(N__30246));
    LocalMux I__7085 (
            .O(N__30246),
            .I(M_this_data_tmp_qZ0Z_4));
    InMux I__7084 (
            .O(N__30243),
            .I(N__30240));
    LocalMux I__7083 (
            .O(N__30240),
            .I(M_this_data_tmp_qZ0Z_0));
    CEMux I__7082 (
            .O(N__30237),
            .I(N__30234));
    LocalMux I__7081 (
            .O(N__30234),
            .I(N__30231));
    Span4Mux_v I__7080 (
            .O(N__30231),
            .I(N__30225));
    CEMux I__7079 (
            .O(N__30230),
            .I(N__30222));
    CEMux I__7078 (
            .O(N__30229),
            .I(N__30219));
    CEMux I__7077 (
            .O(N__30228),
            .I(N__30216));
    Span4Mux_v I__7076 (
            .O(N__30225),
            .I(N__30212));
    LocalMux I__7075 (
            .O(N__30222),
            .I(N__30209));
    LocalMux I__7074 (
            .O(N__30219),
            .I(N__30206));
    LocalMux I__7073 (
            .O(N__30216),
            .I(N__30203));
    CEMux I__7072 (
            .O(N__30215),
            .I(N__30200));
    Span4Mux_h I__7071 (
            .O(N__30212),
            .I(N__30197));
    Span4Mux_v I__7070 (
            .O(N__30209),
            .I(N__30194));
    Span4Mux_h I__7069 (
            .O(N__30206),
            .I(N__30191));
    Span4Mux_h I__7068 (
            .O(N__30203),
            .I(N__30188));
    LocalMux I__7067 (
            .O(N__30200),
            .I(N__30185));
    Odrv4 I__7066 (
            .O(N__30197),
            .I(N_1412_0));
    Odrv4 I__7065 (
            .O(N__30194),
            .I(N_1412_0));
    Odrv4 I__7064 (
            .O(N__30191),
            .I(N_1412_0));
    Odrv4 I__7063 (
            .O(N__30188),
            .I(N_1412_0));
    Odrv12 I__7062 (
            .O(N__30185),
            .I(N_1412_0));
    InMux I__7061 (
            .O(N__30174),
            .I(N__30171));
    LocalMux I__7060 (
            .O(N__30171),
            .I(N__30168));
    Span4Mux_h I__7059 (
            .O(N__30168),
            .I(N__30165));
    Odrv4 I__7058 (
            .O(N__30165),
            .I(M_this_data_tmp_qZ0Z_3));
    InMux I__7057 (
            .O(N__30162),
            .I(N__30159));
    LocalMux I__7056 (
            .O(N__30159),
            .I(N__30156));
    Span4Mux_h I__7055 (
            .O(N__30156),
            .I(N__30153));
    Odrv4 I__7054 (
            .O(N__30153),
            .I(M_this_oam_ram_write_data_3));
    InMux I__7053 (
            .O(N__30150),
            .I(N__30147));
    LocalMux I__7052 (
            .O(N__30147),
            .I(N__30144));
    Span4Mux_h I__7051 (
            .O(N__30144),
            .I(N__30141));
    Odrv4 I__7050 (
            .O(N__30141),
            .I(M_this_oam_ram_write_data_10));
    InMux I__7049 (
            .O(N__30138),
            .I(N__30135));
    LocalMux I__7048 (
            .O(N__30135),
            .I(M_this_data_tmp_qZ0Z_10));
    InMux I__7047 (
            .O(N__30132),
            .I(N__30129));
    LocalMux I__7046 (
            .O(N__30129),
            .I(N__30126));
    Span4Mux_h I__7045 (
            .O(N__30126),
            .I(N__30123));
    Odrv4 I__7044 (
            .O(N__30123),
            .I(M_this_oam_ram_write_data_11));
    CascadeMux I__7043 (
            .O(N__30120),
            .I(N__30117));
    CascadeBuf I__7042 (
            .O(N__30117),
            .I(N__30114));
    CascadeMux I__7041 (
            .O(N__30114),
            .I(N__30111));
    InMux I__7040 (
            .O(N__30111),
            .I(N__30107));
    InMux I__7039 (
            .O(N__30110),
            .I(N__30103));
    LocalMux I__7038 (
            .O(N__30107),
            .I(N__30100));
    InMux I__7037 (
            .O(N__30106),
            .I(N__30097));
    LocalMux I__7036 (
            .O(N__30103),
            .I(N__30094));
    Span4Mux_v I__7035 (
            .O(N__30100),
            .I(N__30091));
    LocalMux I__7034 (
            .O(N__30097),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv4 I__7033 (
            .O(N__30094),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv4 I__7032 (
            .O(N__30091),
            .I(M_this_oam_address_qZ0Z_5));
    CascadeMux I__7031 (
            .O(N__30084),
            .I(N__30081));
    CascadeBuf I__7030 (
            .O(N__30081),
            .I(N__30078));
    CascadeMux I__7029 (
            .O(N__30078),
            .I(N__30074));
    InMux I__7028 (
            .O(N__30077),
            .I(N__30071));
    InMux I__7027 (
            .O(N__30074),
            .I(N__30068));
    LocalMux I__7026 (
            .O(N__30071),
            .I(N__30063));
    LocalMux I__7025 (
            .O(N__30068),
            .I(N__30060));
    InMux I__7024 (
            .O(N__30067),
            .I(N__30055));
    InMux I__7023 (
            .O(N__30066),
            .I(N__30055));
    Span4Mux_h I__7022 (
            .O(N__30063),
            .I(N__30052));
    Span4Mux_v I__7021 (
            .O(N__30060),
            .I(N__30049));
    LocalMux I__7020 (
            .O(N__30055),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv4 I__7019 (
            .O(N__30052),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv4 I__7018 (
            .O(N__30049),
            .I(M_this_oam_address_qZ0Z_4));
    InMux I__7017 (
            .O(N__30042),
            .I(N__30039));
    LocalMux I__7016 (
            .O(N__30039),
            .I(M_this_data_tmp_qZ0Z_11));
    InMux I__7015 (
            .O(N__30036),
            .I(N__30033));
    LocalMux I__7014 (
            .O(N__30033),
            .I(M_this_data_count_q_cry_0_THRU_CO));
    CascadeMux I__7013 (
            .O(N__30030),
            .I(N__30026));
    InMux I__7012 (
            .O(N__30029),
            .I(N__30022));
    InMux I__7011 (
            .O(N__30026),
            .I(N__30019));
    InMux I__7010 (
            .O(N__30025),
            .I(N__30016));
    LocalMux I__7009 (
            .O(N__30022),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__7008 (
            .O(N__30019),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__7007 (
            .O(N__30016),
            .I(M_this_data_count_qZ0Z_1));
    CascadeMux I__7006 (
            .O(N__30009),
            .I(N__30006));
    InMux I__7005 (
            .O(N__30006),
            .I(N__30003));
    LocalMux I__7004 (
            .O(N__30003),
            .I(M_this_data_count_q_cry_2_THRU_CO));
    CascadeMux I__7003 (
            .O(N__30000),
            .I(N__29995));
    CascadeMux I__7002 (
            .O(N__29999),
            .I(N__29992));
    InMux I__7001 (
            .O(N__29998),
            .I(N__29989));
    InMux I__7000 (
            .O(N__29995),
            .I(N__29986));
    InMux I__6999 (
            .O(N__29992),
            .I(N__29983));
    LocalMux I__6998 (
            .O(N__29989),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__6997 (
            .O(N__29986),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__6996 (
            .O(N__29983),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__6995 (
            .O(N__29976),
            .I(N__29973));
    LocalMux I__6994 (
            .O(N__29973),
            .I(M_this_data_count_q_cry_3_THRU_CO));
    InMux I__6993 (
            .O(N__29970),
            .I(N__29965));
    InMux I__6992 (
            .O(N__29969),
            .I(N__29962));
    InMux I__6991 (
            .O(N__29968),
            .I(N__29959));
    LocalMux I__6990 (
            .O(N__29965),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__6989 (
            .O(N__29962),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__6988 (
            .O(N__29959),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__6987 (
            .O(N__29952),
            .I(N__29949));
    LocalMux I__6986 (
            .O(N__29949),
            .I(M_this_data_count_q_cry_4_THRU_CO));
    CascadeMux I__6985 (
            .O(N__29946),
            .I(N__29942));
    InMux I__6984 (
            .O(N__29945),
            .I(N__29938));
    InMux I__6983 (
            .O(N__29942),
            .I(N__29935));
    InMux I__6982 (
            .O(N__29941),
            .I(N__29932));
    LocalMux I__6981 (
            .O(N__29938),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__6980 (
            .O(N__29935),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__6979 (
            .O(N__29932),
            .I(M_this_data_count_qZ0Z_5));
    InMux I__6978 (
            .O(N__29925),
            .I(N__29922));
    LocalMux I__6977 (
            .O(N__29922),
            .I(M_this_data_count_q_cry_5_THRU_CO));
    InMux I__6976 (
            .O(N__29919),
            .I(N__29914));
    InMux I__6975 (
            .O(N__29918),
            .I(N__29911));
    InMux I__6974 (
            .O(N__29917),
            .I(N__29908));
    LocalMux I__6973 (
            .O(N__29914),
            .I(N__29905));
    LocalMux I__6972 (
            .O(N__29911),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__6971 (
            .O(N__29908),
            .I(M_this_data_count_qZ0Z_6));
    Odrv4 I__6970 (
            .O(N__29905),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__6969 (
            .O(N__29898),
            .I(N__29895));
    LocalMux I__6968 (
            .O(N__29895),
            .I(N__29892));
    Span4Mux_h I__6967 (
            .O(N__29892),
            .I(N__29889));
    Odrv4 I__6966 (
            .O(N__29889),
            .I(M_this_oam_ram_write_data_4));
    InMux I__6965 (
            .O(N__29886),
            .I(N__29883));
    LocalMux I__6964 (
            .O(N__29883),
            .I(N__29880));
    Span4Mux_h I__6963 (
            .O(N__29880),
            .I(N__29877));
    Span4Mux_v I__6962 (
            .O(N__29877),
            .I(N__29874));
    Odrv4 I__6961 (
            .O(N__29874),
            .I(M_this_data_tmp_qZ0Z_7));
    InMux I__6960 (
            .O(N__29871),
            .I(N__29868));
    LocalMux I__6959 (
            .O(N__29868),
            .I(N__29865));
    Span4Mux_h I__6958 (
            .O(N__29865),
            .I(N__29862));
    Odrv4 I__6957 (
            .O(N__29862),
            .I(M_this_oam_ram_write_data_7));
    InMux I__6956 (
            .O(N__29859),
            .I(N__29856));
    LocalMux I__6955 (
            .O(N__29856),
            .I(N__29853));
    Odrv12 I__6954 (
            .O(N__29853),
            .I(M_this_oam_ram_write_data_8));
    InMux I__6953 (
            .O(N__29850),
            .I(N__29847));
    LocalMux I__6952 (
            .O(N__29847),
            .I(N__29844));
    Span4Mux_h I__6951 (
            .O(N__29844),
            .I(N__29841));
    Odrv4 I__6950 (
            .O(N__29841),
            .I(M_this_oam_ram_write_data_0));
    CascadeMux I__6949 (
            .O(N__29838),
            .I(N__29835));
    InMux I__6948 (
            .O(N__29835),
            .I(N__29832));
    LocalMux I__6947 (
            .O(N__29832),
            .I(N__29828));
    InMux I__6946 (
            .O(N__29831),
            .I(N__29825));
    Odrv4 I__6945 (
            .O(N__29828),
            .I(M_this_data_count_qZ0Z_14));
    LocalMux I__6944 (
            .O(N__29825),
            .I(M_this_data_count_qZ0Z_14));
    InMux I__6943 (
            .O(N__29820),
            .I(N__29816));
    InMux I__6942 (
            .O(N__29819),
            .I(N__29812));
    LocalMux I__6941 (
            .O(N__29816),
            .I(N__29809));
    InMux I__6940 (
            .O(N__29815),
            .I(N__29806));
    LocalMux I__6939 (
            .O(N__29812),
            .I(M_this_data_count_qZ0Z_13));
    Odrv4 I__6938 (
            .O(N__29809),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__6937 (
            .O(N__29806),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__6936 (
            .O(N__29799),
            .I(N__29795));
    CascadeMux I__6935 (
            .O(N__29798),
            .I(N__29792));
    LocalMux I__6934 (
            .O(N__29795),
            .I(N__29789));
    InMux I__6933 (
            .O(N__29792),
            .I(N__29786));
    Odrv4 I__6932 (
            .O(N__29789),
            .I(M_this_data_count_qZ0Z_15));
    LocalMux I__6931 (
            .O(N__29786),
            .I(M_this_data_count_qZ0Z_15));
    CascadeMux I__6930 (
            .O(N__29781),
            .I(N__29778));
    InMux I__6929 (
            .O(N__29778),
            .I(N__29775));
    LocalMux I__6928 (
            .O(N__29775),
            .I(N__29771));
    InMux I__6927 (
            .O(N__29774),
            .I(N__29768));
    Odrv12 I__6926 (
            .O(N__29771),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__6925 (
            .O(N__29768),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__6924 (
            .O(N__29763),
            .I(N__29758));
    InMux I__6923 (
            .O(N__29762),
            .I(N__29755));
    InMux I__6922 (
            .O(N__29761),
            .I(N__29752));
    LocalMux I__6921 (
            .O(N__29758),
            .I(N__29747));
    LocalMux I__6920 (
            .O(N__29755),
            .I(N__29744));
    LocalMux I__6919 (
            .O(N__29752),
            .I(N__29741));
    InMux I__6918 (
            .O(N__29751),
            .I(N__29736));
    InMux I__6917 (
            .O(N__29750),
            .I(N__29736));
    Odrv4 I__6916 (
            .O(N__29747),
            .I(\this_vga_signals.N_745 ));
    Odrv4 I__6915 (
            .O(N__29744),
            .I(\this_vga_signals.N_745 ));
    Odrv4 I__6914 (
            .O(N__29741),
            .I(\this_vga_signals.N_745 ));
    LocalMux I__6913 (
            .O(N__29736),
            .I(\this_vga_signals.N_745 ));
    InMux I__6912 (
            .O(N__29727),
            .I(N__29724));
    LocalMux I__6911 (
            .O(N__29724),
            .I(\this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2 ));
    InMux I__6910 (
            .O(N__29721),
            .I(N__29718));
    LocalMux I__6909 (
            .O(N__29718),
            .I(\this_vga_signals.N_442_0 ));
    InMux I__6908 (
            .O(N__29715),
            .I(N__29712));
    LocalMux I__6907 (
            .O(N__29712),
            .I(N__29707));
    InMux I__6906 (
            .O(N__29711),
            .I(N__29704));
    InMux I__6905 (
            .O(N__29710),
            .I(N__29701));
    Span4Mux_v I__6904 (
            .O(N__29707),
            .I(N__29692));
    LocalMux I__6903 (
            .O(N__29704),
            .I(N__29692));
    LocalMux I__6902 (
            .O(N__29701),
            .I(N__29689));
    InMux I__6901 (
            .O(N__29700),
            .I(N__29686));
    CascadeMux I__6900 (
            .O(N__29699),
            .I(N__29681));
    IoInMux I__6899 (
            .O(N__29698),
            .I(N__29675));
    InMux I__6898 (
            .O(N__29697),
            .I(N__29672));
    Span4Mux_h I__6897 (
            .O(N__29692),
            .I(N__29669));
    Span4Mux_h I__6896 (
            .O(N__29689),
            .I(N__29666));
    LocalMux I__6895 (
            .O(N__29686),
            .I(N__29663));
    InMux I__6894 (
            .O(N__29685),
            .I(N__29657));
    InMux I__6893 (
            .O(N__29684),
            .I(N__29657));
    InMux I__6892 (
            .O(N__29681),
            .I(N__29652));
    InMux I__6891 (
            .O(N__29680),
            .I(N__29652));
    InMux I__6890 (
            .O(N__29679),
            .I(N__29649));
    InMux I__6889 (
            .O(N__29678),
            .I(N__29646));
    LocalMux I__6888 (
            .O(N__29675),
            .I(N__29643));
    LocalMux I__6887 (
            .O(N__29672),
            .I(N__29640));
    Span4Mux_h I__6886 (
            .O(N__29669),
            .I(N__29633));
    Span4Mux_h I__6885 (
            .O(N__29666),
            .I(N__29633));
    Span4Mux_h I__6884 (
            .O(N__29663),
            .I(N__29633));
    InMux I__6883 (
            .O(N__29662),
            .I(N__29630));
    LocalMux I__6882 (
            .O(N__29657),
            .I(N__29619));
    LocalMux I__6881 (
            .O(N__29652),
            .I(N__29619));
    LocalMux I__6880 (
            .O(N__29649),
            .I(N__29619));
    LocalMux I__6879 (
            .O(N__29646),
            .I(N__29619));
    Span12Mux_s9_h I__6878 (
            .O(N__29643),
            .I(N__29619));
    Odrv4 I__6877 (
            .O(N__29640),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__6876 (
            .O(N__29633),
            .I(M_this_reset_cond_out_0));
    LocalMux I__6875 (
            .O(N__29630),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__6874 (
            .O(N__29619),
            .I(M_this_reset_cond_out_0));
    CascadeMux I__6873 (
            .O(N__29610),
            .I(\this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2_cascade_ ));
    InMux I__6872 (
            .O(N__29607),
            .I(N__29604));
    LocalMux I__6871 (
            .O(N__29604),
            .I(\this_vga_signals.M_this_data_count_qlde_iZ0Z_1 ));
    InMux I__6870 (
            .O(N__29601),
            .I(N__29598));
    LocalMux I__6869 (
            .O(N__29598),
            .I(N__29594));
    InMux I__6868 (
            .O(N__29597),
            .I(N__29591));
    Odrv4 I__6867 (
            .O(N__29594),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__6866 (
            .O(N__29591),
            .I(M_this_data_count_qZ0Z_2));
    InMux I__6865 (
            .O(N__29586),
            .I(N__29581));
    InMux I__6864 (
            .O(N__29585),
            .I(N__29578));
    InMux I__6863 (
            .O(N__29584),
            .I(N__29575));
    LocalMux I__6862 (
            .O(N__29581),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__6861 (
            .O(N__29578),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__6860 (
            .O(N__29575),
            .I(M_this_data_count_qZ0Z_0));
    InMux I__6859 (
            .O(N__29568),
            .I(N__29565));
    LocalMux I__6858 (
            .O(N__29565),
            .I(N__29562));
    Odrv4 I__6857 (
            .O(N__29562),
            .I(M_this_state_d62_11));
    CascadeMux I__6856 (
            .O(N__29559),
            .I(M_this_state_d62_8_cascade_));
    InMux I__6855 (
            .O(N__29556),
            .I(N__29553));
    LocalMux I__6854 (
            .O(N__29553),
            .I(N__29549));
    InMux I__6853 (
            .O(N__29552),
            .I(N__29545));
    Span4Mux_h I__6852 (
            .O(N__29549),
            .I(N__29542));
    InMux I__6851 (
            .O(N__29548),
            .I(N__29539));
    LocalMux I__6850 (
            .O(N__29545),
            .I(N__29536));
    Odrv4 I__6849 (
            .O(N__29542),
            .I(un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2));
    LocalMux I__6848 (
            .O(N__29539),
            .I(un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2));
    Odrv12 I__6847 (
            .O(N__29536),
            .I(un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2));
    CascadeMux I__6846 (
            .O(N__29529),
            .I(M_this_state_d62_cascade_));
    CascadeMux I__6845 (
            .O(N__29526),
            .I(N__29523));
    InMux I__6844 (
            .O(N__29523),
            .I(N__29520));
    LocalMux I__6843 (
            .O(N__29520),
            .I(N__29515));
    InMux I__6842 (
            .O(N__29519),
            .I(N__29512));
    InMux I__6841 (
            .O(N__29518),
            .I(N__29509));
    Span4Mux_v I__6840 (
            .O(N__29515),
            .I(N__29506));
    LocalMux I__6839 (
            .O(N__29512),
            .I(N__29503));
    LocalMux I__6838 (
            .O(N__29509),
            .I(M_this_data_count_qZ0Z_10));
    Odrv4 I__6837 (
            .O(N__29506),
            .I(M_this_data_count_qZ0Z_10));
    Odrv4 I__6836 (
            .O(N__29503),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__6835 (
            .O(N__29496),
            .I(N__29493));
    LocalMux I__6834 (
            .O(N__29493),
            .I(N__29489));
    InMux I__6833 (
            .O(N__29492),
            .I(N__29486));
    Odrv4 I__6832 (
            .O(N__29489),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__6831 (
            .O(N__29486),
            .I(M_this_data_count_qZ0Z_9));
    CascadeMux I__6830 (
            .O(N__29481),
            .I(N__29477));
    InMux I__6829 (
            .O(N__29480),
            .I(N__29474));
    InMux I__6828 (
            .O(N__29477),
            .I(N__29471));
    LocalMux I__6827 (
            .O(N__29474),
            .I(N__29468));
    LocalMux I__6826 (
            .O(N__29471),
            .I(N__29465));
    Odrv4 I__6825 (
            .O(N__29468),
            .I(M_this_data_count_qZ0Z_11));
    Odrv4 I__6824 (
            .O(N__29465),
            .I(M_this_data_count_qZ0Z_11));
    CascadeMux I__6823 (
            .O(N__29460),
            .I(N__29457));
    InMux I__6822 (
            .O(N__29457),
            .I(N__29454));
    LocalMux I__6821 (
            .O(N__29454),
            .I(N__29450));
    InMux I__6820 (
            .O(N__29453),
            .I(N__29447));
    Odrv4 I__6819 (
            .O(N__29450),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__6818 (
            .O(N__29447),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__6817 (
            .O(N__29442),
            .I(N__29439));
    LocalMux I__6816 (
            .O(N__29439),
            .I(M_this_state_d62_10));
    InMux I__6815 (
            .O(N__29436),
            .I(N__29433));
    LocalMux I__6814 (
            .O(N__29433),
            .I(M_this_state_d62_9));
    InMux I__6813 (
            .O(N__29430),
            .I(N__29427));
    LocalMux I__6812 (
            .O(N__29427),
            .I(N__29424));
    Span4Mux_h I__6811 (
            .O(N__29424),
            .I(N__29421));
    Odrv4 I__6810 (
            .O(N__29421),
            .I(M_this_oam_ram_write_data_24));
    InMux I__6809 (
            .O(N__29418),
            .I(N__29413));
    InMux I__6808 (
            .O(N__29417),
            .I(N__29410));
    InMux I__6807 (
            .O(N__29416),
            .I(N__29407));
    LocalMux I__6806 (
            .O(N__29413),
            .I(N__29403));
    LocalMux I__6805 (
            .O(N__29410),
            .I(N__29397));
    LocalMux I__6804 (
            .O(N__29407),
            .I(N__29397));
    InMux I__6803 (
            .O(N__29406),
            .I(N__29394));
    Span4Mux_h I__6802 (
            .O(N__29403),
            .I(N__29391));
    InMux I__6801 (
            .O(N__29402),
            .I(N__29388));
    Span4Mux_h I__6800 (
            .O(N__29397),
            .I(N__29385));
    LocalMux I__6799 (
            .O(N__29394),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__6798 (
            .O(N__29391),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__6797 (
            .O(N__29388),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__6796 (
            .O(N__29385),
            .I(M_this_state_qZ0Z_12));
    CascadeMux I__6795 (
            .O(N__29376),
            .I(N__29370));
    InMux I__6794 (
            .O(N__29375),
            .I(N__29367));
    CascadeMux I__6793 (
            .O(N__29374),
            .I(N__29364));
    InMux I__6792 (
            .O(N__29373),
            .I(N__29360));
    InMux I__6791 (
            .O(N__29370),
            .I(N__29357));
    LocalMux I__6790 (
            .O(N__29367),
            .I(N__29354));
    InMux I__6789 (
            .O(N__29364),
            .I(N__29349));
    InMux I__6788 (
            .O(N__29363),
            .I(N__29349));
    LocalMux I__6787 (
            .O(N__29360),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__6786 (
            .O(N__29357),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__6785 (
            .O(N__29354),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__6784 (
            .O(N__29349),
            .I(M_this_state_qZ0Z_11));
    CascadeMux I__6783 (
            .O(N__29340),
            .I(\this_vga_signals.N_469_0_cascade_ ));
    CascadeMux I__6782 (
            .O(N__29337),
            .I(\this_vga_signals.N_506_cascade_ ));
    InMux I__6781 (
            .O(N__29334),
            .I(N__29331));
    LocalMux I__6780 (
            .O(N__29331),
            .I(N__29326));
    InMux I__6779 (
            .O(N__29330),
            .I(N__29323));
    InMux I__6778 (
            .O(N__29329),
            .I(N__29320));
    Span4Mux_h I__6777 (
            .O(N__29326),
            .I(N__29312));
    LocalMux I__6776 (
            .O(N__29323),
            .I(N__29307));
    LocalMux I__6775 (
            .O(N__29320),
            .I(N__29307));
    InMux I__6774 (
            .O(N__29319),
            .I(N__29300));
    InMux I__6773 (
            .O(N__29318),
            .I(N__29300));
    InMux I__6772 (
            .O(N__29317),
            .I(N__29300));
    InMux I__6771 (
            .O(N__29316),
            .I(N__29292));
    InMux I__6770 (
            .O(N__29315),
            .I(N__29292));
    Span4Mux_v I__6769 (
            .O(N__29312),
            .I(N__29289));
    Span4Mux_v I__6768 (
            .O(N__29307),
            .I(N__29284));
    LocalMux I__6767 (
            .O(N__29300),
            .I(N__29284));
    InMux I__6766 (
            .O(N__29299),
            .I(N__29277));
    InMux I__6765 (
            .O(N__29298),
            .I(N__29277));
    InMux I__6764 (
            .O(N__29297),
            .I(N__29277));
    LocalMux I__6763 (
            .O(N__29292),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__6762 (
            .O(N__29289),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__6761 (
            .O(N__29284),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__6760 (
            .O(N__29277),
            .I(M_this_state_qZ0Z_6));
    CascadeMux I__6759 (
            .O(N__29268),
            .I(\this_ppu.un1_oam_data_c2_cascade_ ));
    InMux I__6758 (
            .O(N__29265),
            .I(N__29262));
    LocalMux I__6757 (
            .O(N__29262),
            .I(\this_ppu.un1_M_vaddress_q_3_6 ));
    InMux I__6756 (
            .O(N__29259),
            .I(N__29256));
    LocalMux I__6755 (
            .O(N__29256),
            .I(M_this_data_tmp_qZ0Z_23));
    InMux I__6754 (
            .O(N__29253),
            .I(N__29250));
    LocalMux I__6753 (
            .O(N__29250),
            .I(N__29247));
    Span4Mux_h I__6752 (
            .O(N__29247),
            .I(N__29244));
    Odrv4 I__6751 (
            .O(N__29244),
            .I(M_this_oam_ram_write_data_23));
    InMux I__6750 (
            .O(N__29241),
            .I(N__29236));
    InMux I__6749 (
            .O(N__29240),
            .I(N__29231));
    InMux I__6748 (
            .O(N__29239),
            .I(N__29231));
    LocalMux I__6747 (
            .O(N__29236),
            .I(N__29228));
    LocalMux I__6746 (
            .O(N__29231),
            .I(N__29225));
    Span12Mux_s7_v I__6745 (
            .O(N__29228),
            .I(N__29222));
    Span4Mux_v I__6744 (
            .O(N__29225),
            .I(N__29219));
    Odrv12 I__6743 (
            .O(N__29222),
            .I(M_this_oam_ram_read_data_22));
    Odrv4 I__6742 (
            .O(N__29219),
            .I(M_this_oam_ram_read_data_22));
    InMux I__6741 (
            .O(N__29214),
            .I(N__29210));
    CascadeMux I__6740 (
            .O(N__29213),
            .I(N__29207));
    LocalMux I__6739 (
            .O(N__29210),
            .I(N__29204));
    InMux I__6738 (
            .O(N__29207),
            .I(N__29201));
    Span4Mux_h I__6737 (
            .O(N__29204),
            .I(N__29198));
    LocalMux I__6736 (
            .O(N__29201),
            .I(N__29195));
    Span4Mux_h I__6735 (
            .O(N__29198),
            .I(N__29192));
    Span4Mux_v I__6734 (
            .O(N__29195),
            .I(N__29189));
    Odrv4 I__6733 (
            .O(N__29192),
            .I(M_this_oam_ram_read_data_23));
    Odrv4 I__6732 (
            .O(N__29189),
            .I(M_this_oam_ram_read_data_23));
    InMux I__6731 (
            .O(N__29184),
            .I(N__29181));
    LocalMux I__6730 (
            .O(N__29181),
            .I(\this_ppu.un1_oam_data_c2 ));
    InMux I__6729 (
            .O(N__29178),
            .I(N__29175));
    LocalMux I__6728 (
            .O(N__29175),
            .I(\this_ppu.un1_M_vaddress_q_3_7 ));
    InMux I__6727 (
            .O(N__29172),
            .I(N__29169));
    LocalMux I__6726 (
            .O(N__29169),
            .I(N__29166));
    Odrv4 I__6725 (
            .O(N__29166),
            .I(M_this_oam_ram_write_data_25));
    CascadeMux I__6724 (
            .O(N__29163),
            .I(N__29160));
    InMux I__6723 (
            .O(N__29160),
            .I(N__29157));
    LocalMux I__6722 (
            .O(N__29157),
            .I(M_this_data_tmp_qZ0Z_17));
    InMux I__6721 (
            .O(N__29154),
            .I(N__29151));
    LocalMux I__6720 (
            .O(N__29151),
            .I(N__29148));
    Span4Mux_h I__6719 (
            .O(N__29148),
            .I(N__29145));
    Odrv4 I__6718 (
            .O(N__29145),
            .I(M_this_oam_ram_write_data_17));
    InMux I__6717 (
            .O(N__29142),
            .I(N__29139));
    LocalMux I__6716 (
            .O(N__29139),
            .I(\this_ppu.un1_M_vaddress_q_3_4 ));
    InMux I__6715 (
            .O(N__29136),
            .I(N__29133));
    LocalMux I__6714 (
            .O(N__29133),
            .I(N__29130));
    Odrv4 I__6713 (
            .O(N__29130),
            .I(M_this_data_count_q_cry_12_THRU_CO));
    InMux I__6712 (
            .O(N__29127),
            .I(M_this_data_count_q_cry_12));
    IoInMux I__6711 (
            .O(N__29124),
            .I(N__29118));
    SRMux I__6710 (
            .O(N__29123),
            .I(N__29114));
    SRMux I__6709 (
            .O(N__29122),
            .I(N__29111));
    SRMux I__6708 (
            .O(N__29121),
            .I(N__29108));
    LocalMux I__6707 (
            .O(N__29118),
            .I(N__29103));
    SRMux I__6706 (
            .O(N__29117),
            .I(N__29099));
    LocalMux I__6705 (
            .O(N__29114),
            .I(N__29093));
    LocalMux I__6704 (
            .O(N__29111),
            .I(N__29093));
    LocalMux I__6703 (
            .O(N__29108),
            .I(N__29090));
    SRMux I__6702 (
            .O(N__29107),
            .I(N__29087));
    SRMux I__6701 (
            .O(N__29106),
            .I(N__29084));
    IoSpan4Mux I__6700 (
            .O(N__29103),
            .I(N__29078));
    SRMux I__6699 (
            .O(N__29102),
            .I(N__29075));
    LocalMux I__6698 (
            .O(N__29099),
            .I(N__29072));
    SRMux I__6697 (
            .O(N__29098),
            .I(N__29069));
    Span4Mux_s3_v I__6696 (
            .O(N__29093),
            .I(N__29052));
    Span4Mux_h I__6695 (
            .O(N__29090),
            .I(N__29052));
    LocalMux I__6694 (
            .O(N__29087),
            .I(N__29052));
    LocalMux I__6693 (
            .O(N__29084),
            .I(N__29052));
    SRMux I__6692 (
            .O(N__29083),
            .I(N__29049));
    SRMux I__6691 (
            .O(N__29082),
            .I(N__29043));
    SRMux I__6690 (
            .O(N__29081),
            .I(N__29039));
    Span4Mux_s2_h I__6689 (
            .O(N__29078),
            .I(N__29036));
    LocalMux I__6688 (
            .O(N__29075),
            .I(N__29029));
    Span4Mux_h I__6687 (
            .O(N__29072),
            .I(N__29029));
    LocalMux I__6686 (
            .O(N__29069),
            .I(N__29029));
    SRMux I__6685 (
            .O(N__29068),
            .I(N__29026));
    SRMux I__6684 (
            .O(N__29067),
            .I(N__29020));
    SRMux I__6683 (
            .O(N__29066),
            .I(N__29017));
    SRMux I__6682 (
            .O(N__29065),
            .I(N__29012));
    CascadeMux I__6681 (
            .O(N__29064),
            .I(N__29007));
    CascadeMux I__6680 (
            .O(N__29063),
            .I(N__29004));
    CascadeMux I__6679 (
            .O(N__29062),
            .I(N__28998));
    SRMux I__6678 (
            .O(N__29061),
            .I(N__28995));
    Span4Mux_v I__6677 (
            .O(N__29052),
            .I(N__28990));
    LocalMux I__6676 (
            .O(N__29049),
            .I(N__28990));
    CascadeMux I__6675 (
            .O(N__29048),
            .I(N__28986));
    CascadeMux I__6674 (
            .O(N__29047),
            .I(N__28982));
    CascadeMux I__6673 (
            .O(N__29046),
            .I(N__28977));
    LocalMux I__6672 (
            .O(N__29043),
            .I(N__28974));
    SRMux I__6671 (
            .O(N__29042),
            .I(N__28971));
    LocalMux I__6670 (
            .O(N__29039),
            .I(N__28968));
    Span4Mux_h I__6669 (
            .O(N__29036),
            .I(N__28961));
    Span4Mux_v I__6668 (
            .O(N__29029),
            .I(N__28961));
    LocalMux I__6667 (
            .O(N__29026),
            .I(N__28961));
    SRMux I__6666 (
            .O(N__29025),
            .I(N__28958));
    SRMux I__6665 (
            .O(N__29024),
            .I(N__28955));
    SRMux I__6664 (
            .O(N__29023),
            .I(N__28952));
    LocalMux I__6663 (
            .O(N__29020),
            .I(N__28949));
    LocalMux I__6662 (
            .O(N__29017),
            .I(N__28946));
    SRMux I__6661 (
            .O(N__29016),
            .I(N__28943));
    SRMux I__6660 (
            .O(N__29015),
            .I(N__28940));
    LocalMux I__6659 (
            .O(N__29012),
            .I(N__28931));
    SRMux I__6658 (
            .O(N__29011),
            .I(N__28928));
    InMux I__6657 (
            .O(N__29010),
            .I(N__28913));
    InMux I__6656 (
            .O(N__29007),
            .I(N__28913));
    InMux I__6655 (
            .O(N__29004),
            .I(N__28913));
    InMux I__6654 (
            .O(N__29003),
            .I(N__28913));
    InMux I__6653 (
            .O(N__29002),
            .I(N__28913));
    InMux I__6652 (
            .O(N__29001),
            .I(N__28913));
    InMux I__6651 (
            .O(N__28998),
            .I(N__28913));
    LocalMux I__6650 (
            .O(N__28995),
            .I(N__28910));
    Span4Mux_v I__6649 (
            .O(N__28990),
            .I(N__28907));
    InMux I__6648 (
            .O(N__28989),
            .I(N__28892));
    InMux I__6647 (
            .O(N__28986),
            .I(N__28892));
    InMux I__6646 (
            .O(N__28985),
            .I(N__28892));
    InMux I__6645 (
            .O(N__28982),
            .I(N__28892));
    InMux I__6644 (
            .O(N__28981),
            .I(N__28892));
    InMux I__6643 (
            .O(N__28980),
            .I(N__28892));
    InMux I__6642 (
            .O(N__28977),
            .I(N__28892));
    Span4Mux_v I__6641 (
            .O(N__28974),
            .I(N__28887));
    LocalMux I__6640 (
            .O(N__28971),
            .I(N__28887));
    Span4Mux_v I__6639 (
            .O(N__28968),
            .I(N__28878));
    Span4Mux_h I__6638 (
            .O(N__28961),
            .I(N__28878));
    LocalMux I__6637 (
            .O(N__28958),
            .I(N__28878));
    LocalMux I__6636 (
            .O(N__28955),
            .I(N__28878));
    LocalMux I__6635 (
            .O(N__28952),
            .I(N__28875));
    Span4Mux_v I__6634 (
            .O(N__28949),
            .I(N__28866));
    Span4Mux_h I__6633 (
            .O(N__28946),
            .I(N__28866));
    LocalMux I__6632 (
            .O(N__28943),
            .I(N__28866));
    LocalMux I__6631 (
            .O(N__28940),
            .I(N__28866));
    SRMux I__6630 (
            .O(N__28939),
            .I(N__28863));
    SRMux I__6629 (
            .O(N__28938),
            .I(N__28860));
    SRMux I__6628 (
            .O(N__28937),
            .I(N__28857));
    SRMux I__6627 (
            .O(N__28936),
            .I(N__28854));
    SRMux I__6626 (
            .O(N__28935),
            .I(N__28847));
    SRMux I__6625 (
            .O(N__28934),
            .I(N__28844));
    Span4Mux_v I__6624 (
            .O(N__28931),
            .I(N__28839));
    LocalMux I__6623 (
            .O(N__28928),
            .I(N__28836));
    LocalMux I__6622 (
            .O(N__28913),
            .I(N__28833));
    Span4Mux_h I__6621 (
            .O(N__28910),
            .I(N__28826));
    Span4Mux_h I__6620 (
            .O(N__28907),
            .I(N__28826));
    LocalMux I__6619 (
            .O(N__28892),
            .I(N__28826));
    Span4Mux_v I__6618 (
            .O(N__28887),
            .I(N__28813));
    Span4Mux_v I__6617 (
            .O(N__28878),
            .I(N__28813));
    Span4Mux_v I__6616 (
            .O(N__28875),
            .I(N__28813));
    Span4Mux_v I__6615 (
            .O(N__28866),
            .I(N__28813));
    LocalMux I__6614 (
            .O(N__28863),
            .I(N__28813));
    LocalMux I__6613 (
            .O(N__28860),
            .I(N__28813));
    LocalMux I__6612 (
            .O(N__28857),
            .I(N__28810));
    LocalMux I__6611 (
            .O(N__28854),
            .I(N__28804));
    SRMux I__6610 (
            .O(N__28853),
            .I(N__28801));
    SRMux I__6609 (
            .O(N__28852),
            .I(N__28798));
    SRMux I__6608 (
            .O(N__28851),
            .I(N__28795));
    SRMux I__6607 (
            .O(N__28850),
            .I(N__28792));
    LocalMux I__6606 (
            .O(N__28847),
            .I(N__28789));
    LocalMux I__6605 (
            .O(N__28844),
            .I(N__28786));
    SRMux I__6604 (
            .O(N__28843),
            .I(N__28783));
    SRMux I__6603 (
            .O(N__28842),
            .I(N__28780));
    Span4Mux_h I__6602 (
            .O(N__28839),
            .I(N__28772));
    Span4Mux_h I__6601 (
            .O(N__28836),
            .I(N__28772));
    Span4Mux_v I__6600 (
            .O(N__28833),
            .I(N__28767));
    Span4Mux_v I__6599 (
            .O(N__28826),
            .I(N__28767));
    Span4Mux_v I__6598 (
            .O(N__28813),
            .I(N__28764));
    Span4Mux_v I__6597 (
            .O(N__28810),
            .I(N__28761));
    CascadeMux I__6596 (
            .O(N__28809),
            .I(N__28758));
    CascadeMux I__6595 (
            .O(N__28808),
            .I(N__28754));
    CascadeMux I__6594 (
            .O(N__28807),
            .I(N__28750));
    Span4Mux_h I__6593 (
            .O(N__28804),
            .I(N__28746));
    LocalMux I__6592 (
            .O(N__28801),
            .I(N__28743));
    LocalMux I__6591 (
            .O(N__28798),
            .I(N__28738));
    LocalMux I__6590 (
            .O(N__28795),
            .I(N__28738));
    LocalMux I__6589 (
            .O(N__28792),
            .I(N__28733));
    Span4Mux_v I__6588 (
            .O(N__28789),
            .I(N__28724));
    Span4Mux_h I__6587 (
            .O(N__28786),
            .I(N__28724));
    LocalMux I__6586 (
            .O(N__28783),
            .I(N__28724));
    LocalMux I__6585 (
            .O(N__28780),
            .I(N__28724));
    SRMux I__6584 (
            .O(N__28779),
            .I(N__28721));
    SRMux I__6583 (
            .O(N__28778),
            .I(N__28718));
    IoInMux I__6582 (
            .O(N__28777),
            .I(N__28714));
    Span4Mux_h I__6581 (
            .O(N__28772),
            .I(N__28711));
    Span4Mux_v I__6580 (
            .O(N__28767),
            .I(N__28704));
    Span4Mux_h I__6579 (
            .O(N__28764),
            .I(N__28704));
    Span4Mux_h I__6578 (
            .O(N__28761),
            .I(N__28704));
    InMux I__6577 (
            .O(N__28758),
            .I(N__28691));
    InMux I__6576 (
            .O(N__28757),
            .I(N__28691));
    InMux I__6575 (
            .O(N__28754),
            .I(N__28691));
    InMux I__6574 (
            .O(N__28753),
            .I(N__28691));
    InMux I__6573 (
            .O(N__28750),
            .I(N__28691));
    InMux I__6572 (
            .O(N__28749),
            .I(N__28691));
    Span4Mux_v I__6571 (
            .O(N__28746),
            .I(N__28686));
    Span4Mux_h I__6570 (
            .O(N__28743),
            .I(N__28686));
    Span4Mux_v I__6569 (
            .O(N__28738),
            .I(N__28683));
    SRMux I__6568 (
            .O(N__28737),
            .I(N__28680));
    SRMux I__6567 (
            .O(N__28736),
            .I(N__28677));
    Span4Mux_v I__6566 (
            .O(N__28733),
            .I(N__28670));
    Span4Mux_v I__6565 (
            .O(N__28724),
            .I(N__28670));
    LocalMux I__6564 (
            .O(N__28721),
            .I(N__28670));
    LocalMux I__6563 (
            .O(N__28718),
            .I(N__28667));
    SRMux I__6562 (
            .O(N__28717),
            .I(N__28664));
    LocalMux I__6561 (
            .O(N__28714),
            .I(N__28661));
    Span4Mux_v I__6560 (
            .O(N__28711),
            .I(N__28653));
    Span4Mux_h I__6559 (
            .O(N__28704),
            .I(N__28653));
    LocalMux I__6558 (
            .O(N__28691),
            .I(N__28653));
    Sp12to4 I__6557 (
            .O(N__28686),
            .I(N__28649));
    Span4Mux_v I__6556 (
            .O(N__28683),
            .I(N__28642));
    LocalMux I__6555 (
            .O(N__28680),
            .I(N__28642));
    LocalMux I__6554 (
            .O(N__28677),
            .I(N__28642));
    Span4Mux_v I__6553 (
            .O(N__28670),
            .I(N__28635));
    Span4Mux_v I__6552 (
            .O(N__28667),
            .I(N__28635));
    LocalMux I__6551 (
            .O(N__28664),
            .I(N__28635));
    IoSpan4Mux I__6550 (
            .O(N__28661),
            .I(N__28632));
    SRMux I__6549 (
            .O(N__28660),
            .I(N__28629));
    Span4Mux_h I__6548 (
            .O(N__28653),
            .I(N__28626));
    SRMux I__6547 (
            .O(N__28652),
            .I(N__28623));
    Span12Mux_h I__6546 (
            .O(N__28649),
            .I(N__28620));
    Span4Mux_v I__6545 (
            .O(N__28642),
            .I(N__28617));
    Span4Mux_h I__6544 (
            .O(N__28635),
            .I(N__28614));
    Span4Mux_s3_h I__6543 (
            .O(N__28632),
            .I(N__28611));
    LocalMux I__6542 (
            .O(N__28629),
            .I(N__28608));
    Span4Mux_h I__6541 (
            .O(N__28626),
            .I(N__28603));
    LocalMux I__6540 (
            .O(N__28623),
            .I(N__28603));
    Span12Mux_v I__6539 (
            .O(N__28620),
            .I(N__28600));
    Span4Mux_v I__6538 (
            .O(N__28617),
            .I(N__28595));
    Span4Mux_v I__6537 (
            .O(N__28614),
            .I(N__28595));
    Span4Mux_v I__6536 (
            .O(N__28611),
            .I(N__28590));
    Span4Mux_v I__6535 (
            .O(N__28608),
            .I(N__28590));
    Span4Mux_h I__6534 (
            .O(N__28603),
            .I(N__28587));
    Odrv12 I__6533 (
            .O(N__28600),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6532 (
            .O(N__28595),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6531 (
            .O(N__28590),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6530 (
            .O(N__28587),
            .I(CONSTANT_ONE_NET));
    InMux I__6529 (
            .O(N__28578),
            .I(N__28575));
    LocalMux I__6528 (
            .O(N__28575),
            .I(N__28572));
    Odrv12 I__6527 (
            .O(N__28572),
            .I(M_this_data_count_q_s_14));
    InMux I__6526 (
            .O(N__28569),
            .I(M_this_data_count_q_cry_13));
    InMux I__6525 (
            .O(N__28566),
            .I(M_this_data_count_q_cry_14));
    InMux I__6524 (
            .O(N__28563),
            .I(N__28560));
    LocalMux I__6523 (
            .O(N__28560),
            .I(N__28557));
    Span4Mux_h I__6522 (
            .O(N__28557),
            .I(N__28554));
    Odrv4 I__6521 (
            .O(N__28554),
            .I(M_this_data_count_q_s_15));
    InMux I__6520 (
            .O(N__28551),
            .I(N__28548));
    LocalMux I__6519 (
            .O(N__28548),
            .I(N__28542));
    InMux I__6518 (
            .O(N__28547),
            .I(N__28537));
    InMux I__6517 (
            .O(N__28546),
            .I(N__28537));
    InMux I__6516 (
            .O(N__28545),
            .I(N__28534));
    Odrv4 I__6515 (
            .O(N__28542),
            .I(\this_vga_signals.N_431_0 ));
    LocalMux I__6514 (
            .O(N__28537),
            .I(\this_vga_signals.N_431_0 ));
    LocalMux I__6513 (
            .O(N__28534),
            .I(\this_vga_signals.N_431_0 ));
    InMux I__6512 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__6511 (
            .O(N__28524),
            .I(N__28518));
    InMux I__6510 (
            .O(N__28523),
            .I(N__28511));
    InMux I__6509 (
            .O(N__28522),
            .I(N__28511));
    InMux I__6508 (
            .O(N__28521),
            .I(N__28511));
    Span4Mux_v I__6507 (
            .O(N__28518),
            .I(N__28507));
    LocalMux I__6506 (
            .O(N__28511),
            .I(N__28504));
    InMux I__6505 (
            .O(N__28510),
            .I(N__28501));
    Odrv4 I__6504 (
            .O(N__28507),
            .I(\this_vga_signals.N_428_0 ));
    Odrv12 I__6503 (
            .O(N__28504),
            .I(\this_vga_signals.N_428_0 ));
    LocalMux I__6502 (
            .O(N__28501),
            .I(\this_vga_signals.N_428_0 ));
    InMux I__6501 (
            .O(N__28494),
            .I(N__28490));
    InMux I__6500 (
            .O(N__28493),
            .I(N__28486));
    LocalMux I__6499 (
            .O(N__28490),
            .I(N__28482));
    InMux I__6498 (
            .O(N__28489),
            .I(N__28479));
    LocalMux I__6497 (
            .O(N__28486),
            .I(N__28476));
    InMux I__6496 (
            .O(N__28485),
            .I(N__28473));
    Span4Mux_h I__6495 (
            .O(N__28482),
            .I(N__28470));
    LocalMux I__6494 (
            .O(N__28479),
            .I(N__28467));
    Span4Mux_v I__6493 (
            .O(N__28476),
            .I(N__28462));
    LocalMux I__6492 (
            .O(N__28473),
            .I(N__28462));
    Span4Mux_v I__6491 (
            .O(N__28470),
            .I(N__28455));
    Span4Mux_h I__6490 (
            .O(N__28467),
            .I(N__28455));
    Span4Mux_v I__6489 (
            .O(N__28462),
            .I(N__28452));
    InMux I__6488 (
            .O(N__28461),
            .I(N__28449));
    InMux I__6487 (
            .O(N__28460),
            .I(N__28446));
    Span4Mux_h I__6486 (
            .O(N__28455),
            .I(N__28441));
    Span4Mux_v I__6485 (
            .O(N__28452),
            .I(N__28436));
    LocalMux I__6484 (
            .O(N__28449),
            .I(N__28436));
    LocalMux I__6483 (
            .O(N__28446),
            .I(N__28433));
    InMux I__6482 (
            .O(N__28445),
            .I(N__28430));
    InMux I__6481 (
            .O(N__28444),
            .I(N__28427));
    Span4Mux_h I__6480 (
            .O(N__28441),
            .I(N__28424));
    Span4Mux_h I__6479 (
            .O(N__28436),
            .I(N__28421));
    Span4Mux_v I__6478 (
            .O(N__28433),
            .I(N__28416));
    LocalMux I__6477 (
            .O(N__28430),
            .I(N__28416));
    LocalMux I__6476 (
            .O(N__28427),
            .I(N__28413));
    Span4Mux_h I__6475 (
            .O(N__28424),
            .I(N__28404));
    Span4Mux_v I__6474 (
            .O(N__28421),
            .I(N__28404));
    Span4Mux_h I__6473 (
            .O(N__28416),
            .I(N__28404));
    Span4Mux_h I__6472 (
            .O(N__28413),
            .I(N__28404));
    Odrv4 I__6471 (
            .O(N__28404),
            .I(N_226));
    InMux I__6470 (
            .O(N__28401),
            .I(N__28398));
    LocalMux I__6469 (
            .O(N__28398),
            .I(M_this_data_tmp_qZ0Z_6));
    InMux I__6468 (
            .O(N__28395),
            .I(N__28392));
    LocalMux I__6467 (
            .O(N__28392),
            .I(N__28389));
    Span4Mux_h I__6466 (
            .O(N__28389),
            .I(N__28386));
    Odrv4 I__6465 (
            .O(N__28386),
            .I(M_this_oam_ram_write_data_6));
    InMux I__6464 (
            .O(N__28383),
            .I(N__28380));
    LocalMux I__6463 (
            .O(N__28380),
            .I(N__28377));
    Span12Mux_s8_v I__6462 (
            .O(N__28377),
            .I(N__28374));
    Odrv12 I__6461 (
            .O(N__28374),
            .I(M_this_data_tmp_qZ0Z_2));
    InMux I__6460 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__6459 (
            .O(N__28368),
            .I(N__28365));
    Span4Mux_v I__6458 (
            .O(N__28365),
            .I(N__28362));
    Odrv4 I__6457 (
            .O(N__28362),
            .I(M_this_oam_ram_write_data_2));
    InMux I__6456 (
            .O(N__28359),
            .I(N__28356));
    LocalMux I__6455 (
            .O(N__28356),
            .I(M_this_data_tmp_qZ0Z_1));
    InMux I__6454 (
            .O(N__28353),
            .I(N__28350));
    LocalMux I__6453 (
            .O(N__28350),
            .I(N__28347));
    Span4Mux_h I__6452 (
            .O(N__28347),
            .I(N__28344));
    Odrv4 I__6451 (
            .O(N__28344),
            .I(M_this_oam_ram_write_data_1));
    InMux I__6450 (
            .O(N__28341),
            .I(M_this_data_count_q_cry_3));
    InMux I__6449 (
            .O(N__28338),
            .I(M_this_data_count_q_cry_4));
    InMux I__6448 (
            .O(N__28335),
            .I(M_this_data_count_q_cry_5));
    InMux I__6447 (
            .O(N__28332),
            .I(M_this_data_count_q_cry_6));
    InMux I__6446 (
            .O(N__28329),
            .I(N__28326));
    LocalMux I__6445 (
            .O(N__28326),
            .I(N__28323));
    Odrv4 I__6444 (
            .O(N__28323),
            .I(M_this_data_count_q_s_8));
    InMux I__6443 (
            .O(N__28320),
            .I(bfn_21_23_0_));
    InMux I__6442 (
            .O(N__28317),
            .I(N__28314));
    LocalMux I__6441 (
            .O(N__28314),
            .I(N__28311));
    Span4Mux_v I__6440 (
            .O(N__28311),
            .I(N__28308));
    Odrv4 I__6439 (
            .O(N__28308),
            .I(M_this_data_count_q_s_9));
    InMux I__6438 (
            .O(N__28305),
            .I(M_this_data_count_q_cry_8));
    InMux I__6437 (
            .O(N__28302),
            .I(N__28299));
    LocalMux I__6436 (
            .O(N__28299),
            .I(N__28296));
    Odrv12 I__6435 (
            .O(N__28296),
            .I(M_this_data_count_q_cry_9_THRU_CO));
    InMux I__6434 (
            .O(N__28293),
            .I(M_this_data_count_q_cry_9));
    InMux I__6433 (
            .O(N__28290),
            .I(N__28287));
    LocalMux I__6432 (
            .O(N__28287),
            .I(N__28284));
    Odrv4 I__6431 (
            .O(N__28284),
            .I(M_this_data_count_q_s_11));
    InMux I__6430 (
            .O(N__28281),
            .I(M_this_data_count_q_cry_10));
    InMux I__6429 (
            .O(N__28278),
            .I(N__28275));
    LocalMux I__6428 (
            .O(N__28275),
            .I(N__28272));
    Odrv4 I__6427 (
            .O(N__28272),
            .I(M_this_data_count_q_s_12));
    InMux I__6426 (
            .O(N__28269),
            .I(M_this_data_count_q_cry_11));
    InMux I__6425 (
            .O(N__28266),
            .I(N__28246));
    InMux I__6424 (
            .O(N__28265),
            .I(N__28246));
    InMux I__6423 (
            .O(N__28264),
            .I(N__28246));
    InMux I__6422 (
            .O(N__28263),
            .I(N__28246));
    InMux I__6421 (
            .O(N__28262),
            .I(N__28246));
    InMux I__6420 (
            .O(N__28261),
            .I(N__28246));
    InMux I__6419 (
            .O(N__28260),
            .I(N__28241));
    InMux I__6418 (
            .O(N__28259),
            .I(N__28241));
    LocalMux I__6417 (
            .O(N__28246),
            .I(N_755));
    LocalMux I__6416 (
            .O(N__28241),
            .I(N_755));
    InMux I__6415 (
            .O(N__28236),
            .I(M_this_data_count_q_cry_0));
    CascadeMux I__6414 (
            .O(N__28233),
            .I(N__28230));
    InMux I__6413 (
            .O(N__28230),
            .I(N__28227));
    LocalMux I__6412 (
            .O(N__28227),
            .I(N__28224));
    Odrv4 I__6411 (
            .O(N__28224),
            .I(M_this_data_count_q_s_2));
    InMux I__6410 (
            .O(N__28221),
            .I(M_this_data_count_q_cry_1));
    InMux I__6409 (
            .O(N__28218),
            .I(M_this_data_count_q_cry_2));
    InMux I__6408 (
            .O(N__28215),
            .I(N__28212));
    LocalMux I__6407 (
            .O(N__28212),
            .I(this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2));
    CascadeMux I__6406 (
            .O(N__28209),
            .I(this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2_cascade_));
    CascadeMux I__6405 (
            .O(N__28206),
            .I(N_307_0_cascade_));
    InMux I__6404 (
            .O(N__28203),
            .I(N__28199));
    InMux I__6403 (
            .O(N__28202),
            .I(N__28196));
    LocalMux I__6402 (
            .O(N__28199),
            .I(N__28188));
    LocalMux I__6401 (
            .O(N__28196),
            .I(N__28185));
    InMux I__6400 (
            .O(N__28195),
            .I(N__28180));
    InMux I__6399 (
            .O(N__28194),
            .I(N__28180));
    InMux I__6398 (
            .O(N__28193),
            .I(N__28177));
    InMux I__6397 (
            .O(N__28192),
            .I(N__28174));
    InMux I__6396 (
            .O(N__28191),
            .I(N__28171));
    Span4Mux_h I__6395 (
            .O(N__28188),
            .I(N__28168));
    Span4Mux_v I__6394 (
            .O(N__28185),
            .I(N__28165));
    LocalMux I__6393 (
            .O(N__28180),
            .I(N__28160));
    LocalMux I__6392 (
            .O(N__28177),
            .I(N__28160));
    LocalMux I__6391 (
            .O(N__28174),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__6390 (
            .O(N__28171),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__6389 (
            .O(N__28168),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__6388 (
            .O(N__28165),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__6387 (
            .O(N__28160),
            .I(M_this_state_qZ0Z_5));
    CascadeMux I__6386 (
            .O(N__28149),
            .I(\this_vga_signals.N_665_1_cascade_ ));
    CascadeMux I__6385 (
            .O(N__28146),
            .I(M_this_data_count_q_3_0_13_cascade_));
    InMux I__6384 (
            .O(N__28143),
            .I(N__28140));
    LocalMux I__6383 (
            .O(N__28140),
            .I(this_vga_signals_un20_i_a2_0_a3_0_a4_2_2));
    InMux I__6382 (
            .O(N__28137),
            .I(N__28134));
    LocalMux I__6381 (
            .O(N__28134),
            .I(N__28131));
    Span4Mux_h I__6380 (
            .O(N__28131),
            .I(N__28128));
    Sp12to4 I__6379 (
            .O(N__28128),
            .I(N__28125));
    Odrv12 I__6378 (
            .O(N__28125),
            .I(\this_sprites_ram.mem_out_bus5_0 ));
    InMux I__6377 (
            .O(N__28122),
            .I(N__28119));
    LocalMux I__6376 (
            .O(N__28119),
            .I(N__28116));
    Span4Mux_v I__6375 (
            .O(N__28116),
            .I(N__28113));
    Odrv4 I__6374 (
            .O(N__28113),
            .I(\this_sprites_ram.mem_out_bus1_0 ));
    InMux I__6373 (
            .O(N__28110),
            .I(N__28105));
    InMux I__6372 (
            .O(N__28109),
            .I(N__28102));
    InMux I__6371 (
            .O(N__28108),
            .I(N__28099));
    LocalMux I__6370 (
            .O(N__28105),
            .I(N__28091));
    LocalMux I__6369 (
            .O(N__28102),
            .I(N__28083));
    LocalMux I__6368 (
            .O(N__28099),
            .I(N__28080));
    InMux I__6367 (
            .O(N__28098),
            .I(N__28071));
    InMux I__6366 (
            .O(N__28097),
            .I(N__28071));
    InMux I__6365 (
            .O(N__28096),
            .I(N__28071));
    InMux I__6364 (
            .O(N__28095),
            .I(N__28071));
    InMux I__6363 (
            .O(N__28094),
            .I(N__28065));
    Span4Mux_h I__6362 (
            .O(N__28091),
            .I(N__28062));
    InMux I__6361 (
            .O(N__28090),
            .I(N__28053));
    InMux I__6360 (
            .O(N__28089),
            .I(N__28053));
    InMux I__6359 (
            .O(N__28088),
            .I(N__28053));
    InMux I__6358 (
            .O(N__28087),
            .I(N__28053));
    InMux I__6357 (
            .O(N__28086),
            .I(N__28050));
    Span4Mux_h I__6356 (
            .O(N__28083),
            .I(N__28043));
    Span4Mux_v I__6355 (
            .O(N__28080),
            .I(N__28043));
    LocalMux I__6354 (
            .O(N__28071),
            .I(N__28043));
    InMux I__6353 (
            .O(N__28070),
            .I(N__28036));
    InMux I__6352 (
            .O(N__28069),
            .I(N__28036));
    InMux I__6351 (
            .O(N__28068),
            .I(N__28036));
    LocalMux I__6350 (
            .O(N__28065),
            .I(N__28033));
    Odrv4 I__6349 (
            .O(N__28062),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__6348 (
            .O(N__28053),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__6347 (
            .O(N__28050),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__6346 (
            .O(N__28043),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    LocalMux I__6345 (
            .O(N__28036),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    Odrv4 I__6344 (
            .O(N__28033),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    InMux I__6343 (
            .O(N__28020),
            .I(N__28017));
    LocalMux I__6342 (
            .O(N__28017),
            .I(N__28014));
    Odrv4 I__6341 (
            .O(N__28014),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ));
    InMux I__6340 (
            .O(N__28011),
            .I(N__28002));
    InMux I__6339 (
            .O(N__28010),
            .I(N__28002));
    InMux I__6338 (
            .O(N__28009),
            .I(N__27997));
    InMux I__6337 (
            .O(N__28008),
            .I(N__27997));
    InMux I__6336 (
            .O(N__28007),
            .I(N__27994));
    LocalMux I__6335 (
            .O(N__28002),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__6334 (
            .O(N__27997),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__6333 (
            .O(N__27994),
            .I(M_this_state_qZ0Z_10));
    CascadeMux I__6332 (
            .O(N__27987),
            .I(\this_vga_signals.N_433_0_cascade_ ));
    CascadeMux I__6331 (
            .O(N__27984),
            .I(\this_vga_signals.N_442_0_cascade_ ));
    CascadeMux I__6330 (
            .O(N__27981),
            .I(\this_vga_signals.N_719_cascade_ ));
    CascadeMux I__6329 (
            .O(N__27978),
            .I(N__27975));
    CascadeBuf I__6328 (
            .O(N__27975),
            .I(N__27972));
    CascadeMux I__6327 (
            .O(N__27972),
            .I(N__27969));
    InMux I__6326 (
            .O(N__27969),
            .I(N__27965));
    InMux I__6325 (
            .O(N__27968),
            .I(N__27962));
    LocalMux I__6324 (
            .O(N__27965),
            .I(N__27959));
    LocalMux I__6323 (
            .O(N__27962),
            .I(N__27955));
    Span4Mux_v I__6322 (
            .O(N__27959),
            .I(N__27952));
    CascadeMux I__6321 (
            .O(N__27958),
            .I(N__27949));
    Span4Mux_h I__6320 (
            .O(N__27955),
            .I(N__27946));
    Sp12to4 I__6319 (
            .O(N__27952),
            .I(N__27943));
    InMux I__6318 (
            .O(N__27949),
            .I(N__27940));
    Sp12to4 I__6317 (
            .O(N__27946),
            .I(N__27937));
    Span12Mux_h I__6316 (
            .O(N__27943),
            .I(N__27934));
    LocalMux I__6315 (
            .O(N__27940),
            .I(M_this_ppu_map_addr_9));
    Odrv12 I__6314 (
            .O(N__27937),
            .I(M_this_ppu_map_addr_9));
    Odrv12 I__6313 (
            .O(N__27934),
            .I(M_this_ppu_map_addr_9));
    CascadeMux I__6312 (
            .O(N__27927),
            .I(N__27924));
    InMux I__6311 (
            .O(N__27924),
            .I(N__27920));
    CascadeMux I__6310 (
            .O(N__27923),
            .I(N__27917));
    LocalMux I__6309 (
            .O(N__27920),
            .I(N__27914));
    InMux I__6308 (
            .O(N__27917),
            .I(N__27911));
    Odrv4 I__6307 (
            .O(N__27914),
            .I(\this_ppu.M_this_ppu_map_addr_i_9 ));
    LocalMux I__6306 (
            .O(N__27911),
            .I(\this_ppu.M_this_ppu_map_addr_i_9 ));
    InMux I__6305 (
            .O(N__27906),
            .I(bfn_21_7_0_));
    InMux I__6304 (
            .O(N__27903),
            .I(N__27900));
    LocalMux I__6303 (
            .O(N__27900),
            .I(N__27897));
    Odrv4 I__6302 (
            .O(N__27897),
            .I(\this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ));
    InMux I__6301 (
            .O(N__27894),
            .I(N__27891));
    LocalMux I__6300 (
            .O(N__27891),
            .I(N__27888));
    Span4Mux_h I__6299 (
            .O(N__27888),
            .I(N__27885));
    Odrv4 I__6298 (
            .O(N__27885),
            .I(M_this_oam_ram_write_data_16));
    InMux I__6297 (
            .O(N__27882),
            .I(N__27879));
    LocalMux I__6296 (
            .O(N__27879),
            .I(M_this_oam_ram_read_data_i_19));
    InMux I__6295 (
            .O(N__27876),
            .I(N__27873));
    LocalMux I__6294 (
            .O(N__27873),
            .I(M_this_data_tmp_qZ0Z_16));
    InMux I__6293 (
            .O(N__27870),
            .I(N__27865));
    InMux I__6292 (
            .O(N__27869),
            .I(N__27861));
    InMux I__6291 (
            .O(N__27868),
            .I(N__27858));
    LocalMux I__6290 (
            .O(N__27865),
            .I(N__27855));
    InMux I__6289 (
            .O(N__27864),
            .I(N__27852));
    LocalMux I__6288 (
            .O(N__27861),
            .I(N__27849));
    LocalMux I__6287 (
            .O(N__27858),
            .I(N__27846));
    Span4Mux_h I__6286 (
            .O(N__27855),
            .I(N__27841));
    LocalMux I__6285 (
            .O(N__27852),
            .I(N__27841));
    Span4Mux_v I__6284 (
            .O(N__27849),
            .I(N__27836));
    Span4Mux_h I__6283 (
            .O(N__27846),
            .I(N__27836));
    Span4Mux_h I__6282 (
            .O(N__27841),
            .I(N__27833));
    Span4Mux_h I__6281 (
            .O(N__27836),
            .I(N__27830));
    Odrv4 I__6280 (
            .O(N__27833),
            .I(M_this_oam_ram_read_data_16));
    Odrv4 I__6279 (
            .O(N__27830),
            .I(M_this_oam_ram_read_data_16));
    InMux I__6278 (
            .O(N__27825),
            .I(N__27820));
    CascadeMux I__6277 (
            .O(N__27824),
            .I(N__27817));
    CascadeMux I__6276 (
            .O(N__27823),
            .I(N__27812));
    LocalMux I__6275 (
            .O(N__27820),
            .I(N__27809));
    InMux I__6274 (
            .O(N__27817),
            .I(N__27806));
    InMux I__6273 (
            .O(N__27816),
            .I(N__27803));
    InMux I__6272 (
            .O(N__27815),
            .I(N__27799));
    InMux I__6271 (
            .O(N__27812),
            .I(N__27796));
    Span4Mux_h I__6270 (
            .O(N__27809),
            .I(N__27793));
    LocalMux I__6269 (
            .O(N__27806),
            .I(N__27790));
    LocalMux I__6268 (
            .O(N__27803),
            .I(N__27784));
    InMux I__6267 (
            .O(N__27802),
            .I(N__27781));
    LocalMux I__6266 (
            .O(N__27799),
            .I(N__27778));
    LocalMux I__6265 (
            .O(N__27796),
            .I(N__27773));
    Span4Mux_v I__6264 (
            .O(N__27793),
            .I(N__27773));
    Span12Mux_v I__6263 (
            .O(N__27790),
            .I(N__27770));
    InMux I__6262 (
            .O(N__27789),
            .I(N__27767));
    InMux I__6261 (
            .O(N__27788),
            .I(N__27762));
    InMux I__6260 (
            .O(N__27787),
            .I(N__27762));
    Span4Mux_h I__6259 (
            .O(N__27784),
            .I(N__27759));
    LocalMux I__6258 (
            .O(N__27781),
            .I(N__27756));
    Span4Mux_h I__6257 (
            .O(N__27778),
            .I(N__27751));
    Span4Mux_v I__6256 (
            .O(N__27773),
            .I(N__27751));
    Odrv12 I__6255 (
            .O(N__27770),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__6254 (
            .O(N__27767),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__6253 (
            .O(N__27762),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__6252 (
            .O(N__27759),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__6251 (
            .O(N__27756),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__6250 (
            .O(N__27751),
            .I(M_this_ppu_vram_addr_7));
    CascadeMux I__6249 (
            .O(N__27738),
            .I(N__27734));
    CascadeMux I__6248 (
            .O(N__27737),
            .I(N__27731));
    InMux I__6247 (
            .O(N__27734),
            .I(N__27728));
    InMux I__6246 (
            .O(N__27731),
            .I(N__27725));
    LocalMux I__6245 (
            .O(N__27728),
            .I(\this_ppu.M_this_ppu_vram_addr_i_7 ));
    LocalMux I__6244 (
            .O(N__27725),
            .I(\this_ppu.M_this_ppu_vram_addr_i_7 ));
    CascadeMux I__6243 (
            .O(N__27720),
            .I(N__27717));
    InMux I__6242 (
            .O(N__27717),
            .I(N__27710));
    InMux I__6241 (
            .O(N__27716),
            .I(N__27707));
    CascadeMux I__6240 (
            .O(N__27715),
            .I(N__27704));
    InMux I__6239 (
            .O(N__27714),
            .I(N__27700));
    InMux I__6238 (
            .O(N__27713),
            .I(N__27697));
    LocalMux I__6237 (
            .O(N__27710),
            .I(N__27694));
    LocalMux I__6236 (
            .O(N__27707),
            .I(N__27691));
    InMux I__6235 (
            .O(N__27704),
            .I(N__27688));
    InMux I__6234 (
            .O(N__27703),
            .I(N__27685));
    LocalMux I__6233 (
            .O(N__27700),
            .I(N__27682));
    LocalMux I__6232 (
            .O(N__27697),
            .I(N__27679));
    Span4Mux_v I__6231 (
            .O(N__27694),
            .I(N__27676));
    Span12Mux_h I__6230 (
            .O(N__27691),
            .I(N__27673));
    LocalMux I__6229 (
            .O(N__27688),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    LocalMux I__6228 (
            .O(N__27685),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv4 I__6227 (
            .O(N__27682),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv4 I__6226 (
            .O(N__27679),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv4 I__6225 (
            .O(N__27676),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv12 I__6224 (
            .O(N__27673),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    InMux I__6223 (
            .O(N__27660),
            .I(N__27656));
    InMux I__6222 (
            .O(N__27659),
            .I(N__27652));
    LocalMux I__6221 (
            .O(N__27656),
            .I(N__27649));
    InMux I__6220 (
            .O(N__27655),
            .I(N__27646));
    LocalMux I__6219 (
            .O(N__27652),
            .I(N__27643));
    Span4Mux_h I__6218 (
            .O(N__27649),
            .I(N__27638));
    LocalMux I__6217 (
            .O(N__27646),
            .I(N__27638));
    Span4Mux_h I__6216 (
            .O(N__27643),
            .I(N__27635));
    Span4Mux_h I__6215 (
            .O(N__27638),
            .I(N__27632));
    Span4Mux_h I__6214 (
            .O(N__27635),
            .I(N__27629));
    Odrv4 I__6213 (
            .O(N__27632),
            .I(M_this_oam_ram_read_data_17));
    Odrv4 I__6212 (
            .O(N__27629),
            .I(M_this_oam_ram_read_data_17));
    CascadeMux I__6211 (
            .O(N__27624),
            .I(N__27620));
    CascadeMux I__6210 (
            .O(N__27623),
            .I(N__27617));
    InMux I__6209 (
            .O(N__27620),
            .I(N__27614));
    InMux I__6208 (
            .O(N__27617),
            .I(N__27611));
    LocalMux I__6207 (
            .O(N__27614),
            .I(\this_ppu.M_vaddress_q_i_1 ));
    LocalMux I__6206 (
            .O(N__27611),
            .I(\this_ppu.M_vaddress_q_i_1 ));
    CascadeMux I__6205 (
            .O(N__27606),
            .I(N__27598));
    InMux I__6204 (
            .O(N__27605),
            .I(N__27595));
    InMux I__6203 (
            .O(N__27604),
            .I(N__27592));
    InMux I__6202 (
            .O(N__27603),
            .I(N__27589));
    CascadeMux I__6201 (
            .O(N__27602),
            .I(N__27586));
    InMux I__6200 (
            .O(N__27601),
            .I(N__27580));
    InMux I__6199 (
            .O(N__27598),
            .I(N__27580));
    LocalMux I__6198 (
            .O(N__27595),
            .I(N__27577));
    LocalMux I__6197 (
            .O(N__27592),
            .I(N__27574));
    LocalMux I__6196 (
            .O(N__27589),
            .I(N__27571));
    InMux I__6195 (
            .O(N__27586),
            .I(N__27568));
    InMux I__6194 (
            .O(N__27585),
            .I(N__27565));
    LocalMux I__6193 (
            .O(N__27580),
            .I(N__27562));
    Span4Mux_h I__6192 (
            .O(N__27577),
            .I(N__27557));
    Span4Mux_h I__6191 (
            .O(N__27574),
            .I(N__27557));
    Span12Mux_v I__6190 (
            .O(N__27571),
            .I(N__27554));
    LocalMux I__6189 (
            .O(N__27568),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__6188 (
            .O(N__27565),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    Odrv4 I__6187 (
            .O(N__27562),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    Odrv4 I__6186 (
            .O(N__27557),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    Odrv12 I__6185 (
            .O(N__27554),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    CascadeMux I__6184 (
            .O(N__27543),
            .I(N__27540));
    InMux I__6183 (
            .O(N__27540),
            .I(N__27535));
    InMux I__6182 (
            .O(N__27539),
            .I(N__27532));
    CascadeMux I__6181 (
            .O(N__27538),
            .I(N__27529));
    LocalMux I__6180 (
            .O(N__27535),
            .I(N__27526));
    LocalMux I__6179 (
            .O(N__27532),
            .I(N__27523));
    InMux I__6178 (
            .O(N__27529),
            .I(N__27520));
    Span4Mux_v I__6177 (
            .O(N__27526),
            .I(N__27517));
    Span4Mux_v I__6176 (
            .O(N__27523),
            .I(N__27514));
    LocalMux I__6175 (
            .O(N__27520),
            .I(N__27511));
    Span4Mux_h I__6174 (
            .O(N__27517),
            .I(N__27508));
    Span4Mux_h I__6173 (
            .O(N__27514),
            .I(N__27503));
    Span4Mux_v I__6172 (
            .O(N__27511),
            .I(N__27503));
    Odrv4 I__6171 (
            .O(N__27508),
            .I(M_this_oam_ram_read_data_18));
    Odrv4 I__6170 (
            .O(N__27503),
            .I(M_this_oam_ram_read_data_18));
    InMux I__6169 (
            .O(N__27498),
            .I(N__27494));
    InMux I__6168 (
            .O(N__27497),
            .I(N__27491));
    LocalMux I__6167 (
            .O(N__27494),
            .I(\this_ppu.M_vaddress_q_i_2 ));
    LocalMux I__6166 (
            .O(N__27491),
            .I(\this_ppu.M_vaddress_q_i_2 ));
    CascadeMux I__6165 (
            .O(N__27486),
            .I(N__27483));
    CascadeBuf I__6164 (
            .O(N__27483),
            .I(N__27480));
    CascadeMux I__6163 (
            .O(N__27480),
            .I(N__27477));
    InMux I__6162 (
            .O(N__27477),
            .I(N__27473));
    InMux I__6161 (
            .O(N__27476),
            .I(N__27469));
    LocalMux I__6160 (
            .O(N__27473),
            .I(N__27466));
    InMux I__6159 (
            .O(N__27472),
            .I(N__27463));
    LocalMux I__6158 (
            .O(N__27469),
            .I(N__27458));
    Sp12to4 I__6157 (
            .O(N__27466),
            .I(N__27455));
    LocalMux I__6156 (
            .O(N__27463),
            .I(N__27452));
    InMux I__6155 (
            .O(N__27462),
            .I(N__27447));
    InMux I__6154 (
            .O(N__27461),
            .I(N__27447));
    Span12Mux_v I__6153 (
            .O(N__27458),
            .I(N__27442));
    Span12Mux_v I__6152 (
            .O(N__27455),
            .I(N__27442));
    Odrv4 I__6151 (
            .O(N__27452),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__6150 (
            .O(N__27447),
            .I(M_this_ppu_map_addr_5));
    Odrv12 I__6149 (
            .O(N__27442),
            .I(M_this_ppu_map_addr_5));
    CascadeMux I__6148 (
            .O(N__27435),
            .I(N__27431));
    CascadeMux I__6147 (
            .O(N__27434),
            .I(N__27428));
    InMux I__6146 (
            .O(N__27431),
            .I(N__27425));
    InMux I__6145 (
            .O(N__27428),
            .I(N__27422));
    LocalMux I__6144 (
            .O(N__27425),
            .I(\this_ppu.M_this_ppu_map_addr_i_5 ));
    LocalMux I__6143 (
            .O(N__27422),
            .I(\this_ppu.M_this_ppu_map_addr_i_5 ));
    CascadeMux I__6142 (
            .O(N__27417),
            .I(N__27414));
    CascadeBuf I__6141 (
            .O(N__27414),
            .I(N__27411));
    CascadeMux I__6140 (
            .O(N__27411),
            .I(N__27408));
    InMux I__6139 (
            .O(N__27408),
            .I(N__27405));
    LocalMux I__6138 (
            .O(N__27405),
            .I(N__27401));
    InMux I__6137 (
            .O(N__27404),
            .I(N__27396));
    Span4Mux_v I__6136 (
            .O(N__27401),
            .I(N__27393));
    CascadeMux I__6135 (
            .O(N__27400),
            .I(N__27390));
    InMux I__6134 (
            .O(N__27399),
            .I(N__27387));
    LocalMux I__6133 (
            .O(N__27396),
            .I(N__27384));
    Sp12to4 I__6132 (
            .O(N__27393),
            .I(N__27381));
    InMux I__6131 (
            .O(N__27390),
            .I(N__27378));
    LocalMux I__6130 (
            .O(N__27387),
            .I(N__27375));
    Span12Mux_v I__6129 (
            .O(N__27384),
            .I(N__27370));
    Span12Mux_v I__6128 (
            .O(N__27381),
            .I(N__27370));
    LocalMux I__6127 (
            .O(N__27378),
            .I(M_this_ppu_map_addr_6));
    Odrv4 I__6126 (
            .O(N__27375),
            .I(M_this_ppu_map_addr_6));
    Odrv12 I__6125 (
            .O(N__27370),
            .I(M_this_ppu_map_addr_6));
    CascadeMux I__6124 (
            .O(N__27363),
            .I(N__27359));
    CascadeMux I__6123 (
            .O(N__27362),
            .I(N__27356));
    InMux I__6122 (
            .O(N__27359),
            .I(N__27353));
    InMux I__6121 (
            .O(N__27356),
            .I(N__27350));
    LocalMux I__6120 (
            .O(N__27353),
            .I(N__27347));
    LocalMux I__6119 (
            .O(N__27350),
            .I(\this_ppu.M_this_ppu_map_addr_i_6 ));
    Odrv4 I__6118 (
            .O(N__27347),
            .I(\this_ppu.M_this_ppu_map_addr_i_6 ));
    CascadeMux I__6117 (
            .O(N__27342),
            .I(N__27339));
    CascadeBuf I__6116 (
            .O(N__27339),
            .I(N__27336));
    CascadeMux I__6115 (
            .O(N__27336),
            .I(N__27332));
    InMux I__6114 (
            .O(N__27335),
            .I(N__27329));
    InMux I__6113 (
            .O(N__27332),
            .I(N__27326));
    LocalMux I__6112 (
            .O(N__27329),
            .I(N__27323));
    LocalMux I__6111 (
            .O(N__27326),
            .I(N__27320));
    Span4Mux_h I__6110 (
            .O(N__27323),
            .I(N__27314));
    Span12Mux_h I__6109 (
            .O(N__27320),
            .I(N__27311));
    InMux I__6108 (
            .O(N__27319),
            .I(N__27308));
    InMux I__6107 (
            .O(N__27318),
            .I(N__27303));
    InMux I__6106 (
            .O(N__27317),
            .I(N__27303));
    Sp12to4 I__6105 (
            .O(N__27314),
            .I(N__27298));
    Span12Mux_v I__6104 (
            .O(N__27311),
            .I(N__27298));
    LocalMux I__6103 (
            .O(N__27308),
            .I(M_this_ppu_map_addr_7));
    LocalMux I__6102 (
            .O(N__27303),
            .I(M_this_ppu_map_addr_7));
    Odrv12 I__6101 (
            .O(N__27298),
            .I(M_this_ppu_map_addr_7));
    CascadeMux I__6100 (
            .O(N__27291),
            .I(N__27287));
    InMux I__6099 (
            .O(N__27290),
            .I(N__27284));
    InMux I__6098 (
            .O(N__27287),
            .I(N__27281));
    LocalMux I__6097 (
            .O(N__27284),
            .I(\this_ppu.M_this_ppu_map_addr_i_7 ));
    LocalMux I__6096 (
            .O(N__27281),
            .I(\this_ppu.M_this_ppu_map_addr_i_7 ));
    CascadeMux I__6095 (
            .O(N__27276),
            .I(N__27273));
    CascadeBuf I__6094 (
            .O(N__27273),
            .I(N__27269));
    InMux I__6093 (
            .O(N__27272),
            .I(N__27266));
    CascadeMux I__6092 (
            .O(N__27269),
            .I(N__27263));
    LocalMux I__6091 (
            .O(N__27266),
            .I(N__27260));
    InMux I__6090 (
            .O(N__27263),
            .I(N__27257));
    Span4Mux_h I__6089 (
            .O(N__27260),
            .I(N__27254));
    LocalMux I__6088 (
            .O(N__27257),
            .I(N__27251));
    Span4Mux_v I__6087 (
            .O(N__27254),
            .I(N__27246));
    Span12Mux_s5_v I__6086 (
            .O(N__27251),
            .I(N__27243));
    InMux I__6085 (
            .O(N__27250),
            .I(N__27240));
    InMux I__6084 (
            .O(N__27249),
            .I(N__27237));
    Span4Mux_v I__6083 (
            .O(N__27246),
            .I(N__27234));
    Span12Mux_v I__6082 (
            .O(N__27243),
            .I(N__27231));
    LocalMux I__6081 (
            .O(N__27240),
            .I(M_this_ppu_map_addr_8));
    LocalMux I__6080 (
            .O(N__27237),
            .I(M_this_ppu_map_addr_8));
    Odrv4 I__6079 (
            .O(N__27234),
            .I(M_this_ppu_map_addr_8));
    Odrv12 I__6078 (
            .O(N__27231),
            .I(M_this_ppu_map_addr_8));
    CascadeMux I__6077 (
            .O(N__27222),
            .I(N__27218));
    CascadeMux I__6076 (
            .O(N__27221),
            .I(N__27215));
    InMux I__6075 (
            .O(N__27218),
            .I(N__27212));
    InMux I__6074 (
            .O(N__27215),
            .I(N__27209));
    LocalMux I__6073 (
            .O(N__27212),
            .I(\this_ppu.M_this_ppu_map_addr_i_8 ));
    LocalMux I__6072 (
            .O(N__27209),
            .I(\this_ppu.M_this_ppu_map_addr_i_8 ));
    CascadeMux I__6071 (
            .O(N__27204),
            .I(N__27201));
    InMux I__6070 (
            .O(N__27201),
            .I(N__27198));
    LocalMux I__6069 (
            .O(N__27198),
            .I(N__27194));
    CascadeMux I__6068 (
            .O(N__27197),
            .I(N__27191));
    Span4Mux_v I__6067 (
            .O(N__27194),
            .I(N__27188));
    InMux I__6066 (
            .O(N__27191),
            .I(N__27185));
    Odrv4 I__6065 (
            .O(N__27188),
            .I(N_460_0));
    LocalMux I__6064 (
            .O(N__27185),
            .I(N_460_0));
    CascadeMux I__6063 (
            .O(N__27180),
            .I(N__27176));
    InMux I__6062 (
            .O(N__27179),
            .I(N__27173));
    InMux I__6061 (
            .O(N__27176),
            .I(N__27170));
    LocalMux I__6060 (
            .O(N__27173),
            .I(N__27165));
    LocalMux I__6059 (
            .O(N__27170),
            .I(N__27162));
    InMux I__6058 (
            .O(N__27169),
            .I(N__27155));
    InMux I__6057 (
            .O(N__27168),
            .I(N__27155));
    Span4Mux_v I__6056 (
            .O(N__27165),
            .I(N__27151));
    Span4Mux_v I__6055 (
            .O(N__27162),
            .I(N__27148));
    InMux I__6054 (
            .O(N__27161),
            .I(N__27143));
    InMux I__6053 (
            .O(N__27160),
            .I(N__27143));
    LocalMux I__6052 (
            .O(N__27155),
            .I(N__27140));
    InMux I__6051 (
            .O(N__27154),
            .I(N__27137));
    Odrv4 I__6050 (
            .O(N__27151),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__6049 (
            .O(N__27148),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__6048 (
            .O(N__27143),
            .I(M_this_state_qZ0Z_8));
    Odrv12 I__6047 (
            .O(N__27140),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__6046 (
            .O(N__27137),
            .I(M_this_state_qZ0Z_8));
    InMux I__6045 (
            .O(N__27126),
            .I(N__27118));
    InMux I__6044 (
            .O(N__27125),
            .I(N__27118));
    InMux I__6043 (
            .O(N__27124),
            .I(N__27115));
    InMux I__6042 (
            .O(N__27123),
            .I(N__27112));
    LocalMux I__6041 (
            .O(N__27118),
            .I(N__27107));
    LocalMux I__6040 (
            .O(N__27115),
            .I(N__27102));
    LocalMux I__6039 (
            .O(N__27112),
            .I(N__27102));
    InMux I__6038 (
            .O(N__27111),
            .I(N__27097));
    InMux I__6037 (
            .O(N__27110),
            .I(N__27097));
    Odrv4 I__6036 (
            .O(N__27107),
            .I(M_this_state_qZ0Z_3));
    Odrv12 I__6035 (
            .O(N__27102),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__6034 (
            .O(N__27097),
            .I(M_this_state_qZ0Z_3));
    InMux I__6033 (
            .O(N__27090),
            .I(N__27087));
    LocalMux I__6032 (
            .O(N__27087),
            .I(N__27084));
    Odrv4 I__6031 (
            .O(N__27084),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_2 ));
    InMux I__6030 (
            .O(N__27081),
            .I(N__27077));
    InMux I__6029 (
            .O(N__27080),
            .I(N__27074));
    LocalMux I__6028 (
            .O(N__27077),
            .I(N__27068));
    LocalMux I__6027 (
            .O(N__27074),
            .I(N__27068));
    InMux I__6026 (
            .O(N__27073),
            .I(N__27065));
    Span4Mux_h I__6025 (
            .O(N__27068),
            .I(N__27062));
    LocalMux I__6024 (
            .O(N__27065),
            .I(N__27059));
    Odrv4 I__6023 (
            .O(N__27062),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1 ));
    Odrv4 I__6022 (
            .O(N__27059),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1 ));
    InMux I__6021 (
            .O(N__27054),
            .I(N__27039));
    InMux I__6020 (
            .O(N__27053),
            .I(N__27033));
    InMux I__6019 (
            .O(N__27052),
            .I(N__27026));
    InMux I__6018 (
            .O(N__27051),
            .I(N__27026));
    InMux I__6017 (
            .O(N__27050),
            .I(N__27026));
    InMux I__6016 (
            .O(N__27049),
            .I(N__27023));
    InMux I__6015 (
            .O(N__27048),
            .I(N__27018));
    InMux I__6014 (
            .O(N__27047),
            .I(N__27018));
    InMux I__6013 (
            .O(N__27046),
            .I(N__27011));
    InMux I__6012 (
            .O(N__27045),
            .I(N__27011));
    InMux I__6011 (
            .O(N__27044),
            .I(N__27008));
    InMux I__6010 (
            .O(N__27043),
            .I(N__27002));
    InMux I__6009 (
            .O(N__27042),
            .I(N__26999));
    LocalMux I__6008 (
            .O(N__27039),
            .I(N__26996));
    InMux I__6007 (
            .O(N__27038),
            .I(N__26993));
    InMux I__6006 (
            .O(N__27037),
            .I(N__26990));
    CascadeMux I__6005 (
            .O(N__27036),
            .I(N__26986));
    LocalMux I__6004 (
            .O(N__27033),
            .I(N__26980));
    LocalMux I__6003 (
            .O(N__27026),
            .I(N__26980));
    LocalMux I__6002 (
            .O(N__27023),
            .I(N__26975));
    LocalMux I__6001 (
            .O(N__27018),
            .I(N__26975));
    InMux I__6000 (
            .O(N__27017),
            .I(N__26970));
    InMux I__5999 (
            .O(N__27016),
            .I(N__26970));
    LocalMux I__5998 (
            .O(N__27011),
            .I(N__26965));
    LocalMux I__5997 (
            .O(N__27008),
            .I(N__26965));
    InMux I__5996 (
            .O(N__27007),
            .I(N__26960));
    InMux I__5995 (
            .O(N__27006),
            .I(N__26960));
    InMux I__5994 (
            .O(N__27005),
            .I(N__26957));
    LocalMux I__5993 (
            .O(N__27002),
            .I(N__26954));
    LocalMux I__5992 (
            .O(N__26999),
            .I(N__26951));
    Span4Mux_v I__5991 (
            .O(N__26996),
            .I(N__26946));
    LocalMux I__5990 (
            .O(N__26993),
            .I(N__26946));
    LocalMux I__5989 (
            .O(N__26990),
            .I(N__26943));
    InMux I__5988 (
            .O(N__26989),
            .I(N__26936));
    InMux I__5987 (
            .O(N__26986),
            .I(N__26931));
    InMux I__5986 (
            .O(N__26985),
            .I(N__26931));
    Span4Mux_h I__5985 (
            .O(N__26980),
            .I(N__26920));
    Span4Mux_v I__5984 (
            .O(N__26975),
            .I(N__26920));
    LocalMux I__5983 (
            .O(N__26970),
            .I(N__26920));
    Span4Mux_v I__5982 (
            .O(N__26965),
            .I(N__26920));
    LocalMux I__5981 (
            .O(N__26960),
            .I(N__26920));
    LocalMux I__5980 (
            .O(N__26957),
            .I(N__26915));
    Span4Mux_h I__5979 (
            .O(N__26954),
            .I(N__26915));
    Span4Mux_v I__5978 (
            .O(N__26951),
            .I(N__26910));
    Span4Mux_h I__5977 (
            .O(N__26946),
            .I(N__26910));
    Span12Mux_v I__5976 (
            .O(N__26943),
            .I(N__26907));
    InMux I__5975 (
            .O(N__26942),
            .I(N__26898));
    InMux I__5974 (
            .O(N__26941),
            .I(N__26898));
    InMux I__5973 (
            .O(N__26940),
            .I(N__26898));
    InMux I__5972 (
            .O(N__26939),
            .I(N__26898));
    LocalMux I__5971 (
            .O(N__26936),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__5970 (
            .O(N__26931),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__5969 (
            .O(N__26920),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__5968 (
            .O(N__26915),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__5967 (
            .O(N__26910),
            .I(M_this_state_qZ0Z_2));
    Odrv12 I__5966 (
            .O(N__26907),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__5965 (
            .O(N__26898),
            .I(M_this_state_qZ0Z_2));
    InMux I__5964 (
            .O(N__26883),
            .I(N__26880));
    LocalMux I__5963 (
            .O(N__26880),
            .I(N__26874));
    InMux I__5962 (
            .O(N__26879),
            .I(N__26871));
    InMux I__5961 (
            .O(N__26878),
            .I(N__26868));
    InMux I__5960 (
            .O(N__26877),
            .I(N__26865));
    Span4Mux_v I__5959 (
            .O(N__26874),
            .I(N__26860));
    LocalMux I__5958 (
            .O(N__26871),
            .I(N__26860));
    LocalMux I__5957 (
            .O(N__26868),
            .I(N__26857));
    LocalMux I__5956 (
            .O(N__26865),
            .I(N__26850));
    Span4Mux_v I__5955 (
            .O(N__26860),
            .I(N__26845));
    Span4Mux_h I__5954 (
            .O(N__26857),
            .I(N__26845));
    InMux I__5953 (
            .O(N__26856),
            .I(N__26842));
    InMux I__5952 (
            .O(N__26855),
            .I(N__26839));
    InMux I__5951 (
            .O(N__26854),
            .I(N__26836));
    InMux I__5950 (
            .O(N__26853),
            .I(N__26833));
    Span4Mux_s3_v I__5949 (
            .O(N__26850),
            .I(N__26830));
    Span4Mux_v I__5948 (
            .O(N__26845),
            .I(N__26827));
    LocalMux I__5947 (
            .O(N__26842),
            .I(N__26824));
    LocalMux I__5946 (
            .O(N__26839),
            .I(N__26821));
    LocalMux I__5945 (
            .O(N__26836),
            .I(N__26818));
    LocalMux I__5944 (
            .O(N__26833),
            .I(N__26815));
    Span4Mux_v I__5943 (
            .O(N__26830),
            .I(N__26808));
    Span4Mux_v I__5942 (
            .O(N__26827),
            .I(N__26808));
    Span4Mux_h I__5941 (
            .O(N__26824),
            .I(N__26808));
    Span12Mux_h I__5940 (
            .O(N__26821),
            .I(N__26805));
    Span12Mux_h I__5939 (
            .O(N__26818),
            .I(N__26800));
    Span12Mux_h I__5938 (
            .O(N__26815),
            .I(N__26800));
    Span4Mux_h I__5937 (
            .O(N__26808),
            .I(N__26797));
    Odrv12 I__5936 (
            .O(N__26805),
            .I(N_250));
    Odrv12 I__5935 (
            .O(N__26800),
            .I(N_250));
    Odrv4 I__5934 (
            .O(N__26797),
            .I(N_250));
    CascadeMux I__5933 (
            .O(N__26790),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3Z0Z_0_cascade_ ));
    CascadeMux I__5932 (
            .O(N__26787),
            .I(N__26784));
    InMux I__5931 (
            .O(N__26784),
            .I(N__26780));
    CascadeMux I__5930 (
            .O(N__26783),
            .I(N__26777));
    LocalMux I__5929 (
            .O(N__26780),
            .I(N__26772));
    InMux I__5928 (
            .O(N__26777),
            .I(N__26765));
    InMux I__5927 (
            .O(N__26776),
            .I(N__26765));
    InMux I__5926 (
            .O(N__26775),
            .I(N__26765));
    Span4Mux_h I__5925 (
            .O(N__26772),
            .I(N__26762));
    LocalMux I__5924 (
            .O(N__26765),
            .I(N__26759));
    Odrv4 I__5923 (
            .O(N__26762),
            .I(\this_vga_signals.N_743 ));
    Odrv12 I__5922 (
            .O(N__26759),
            .I(\this_vga_signals.N_743 ));
    InMux I__5921 (
            .O(N__26754),
            .I(N__26750));
    InMux I__5920 (
            .O(N__26753),
            .I(N__26741));
    LocalMux I__5919 (
            .O(N__26750),
            .I(N__26738));
    InMux I__5918 (
            .O(N__26749),
            .I(N__26735));
    InMux I__5917 (
            .O(N__26748),
            .I(N__26732));
    InMux I__5916 (
            .O(N__26747),
            .I(N__26729));
    InMux I__5915 (
            .O(N__26746),
            .I(N__26726));
    InMux I__5914 (
            .O(N__26745),
            .I(N__26723));
    InMux I__5913 (
            .O(N__26744),
            .I(N__26720));
    LocalMux I__5912 (
            .O(N__26741),
            .I(N__26717));
    Span4Mux_v I__5911 (
            .O(N__26738),
            .I(N__26714));
    LocalMux I__5910 (
            .O(N__26735),
            .I(N__26709));
    LocalMux I__5909 (
            .O(N__26732),
            .I(N__26709));
    LocalMux I__5908 (
            .O(N__26729),
            .I(N__26706));
    LocalMux I__5907 (
            .O(N__26726),
            .I(N__26703));
    LocalMux I__5906 (
            .O(N__26723),
            .I(N__26698));
    LocalMux I__5905 (
            .O(N__26720),
            .I(N__26698));
    Span4Mux_v I__5904 (
            .O(N__26717),
            .I(N__26693));
    Span4Mux_v I__5903 (
            .O(N__26714),
            .I(N__26693));
    Span4Mux_v I__5902 (
            .O(N__26709),
            .I(N__26690));
    Span4Mux_v I__5901 (
            .O(N__26706),
            .I(N__26685));
    Span4Mux_v I__5900 (
            .O(N__26703),
            .I(N__26685));
    Span12Mux_v I__5899 (
            .O(N__26698),
            .I(N__26682));
    Sp12to4 I__5898 (
            .O(N__26693),
            .I(N__26679));
    Span4Mux_h I__5897 (
            .O(N__26690),
            .I(N__26674));
    Span4Mux_h I__5896 (
            .O(N__26685),
            .I(N__26674));
    Span12Mux_h I__5895 (
            .O(N__26682),
            .I(N__26669));
    Span12Mux_h I__5894 (
            .O(N__26679),
            .I(N__26669));
    Odrv4 I__5893 (
            .O(N__26674),
            .I(N_228));
    Odrv12 I__5892 (
            .O(N__26669),
            .I(N_228));
    InMux I__5891 (
            .O(N__26664),
            .I(N__26657));
    InMux I__5890 (
            .O(N__26663),
            .I(N__26654));
    InMux I__5889 (
            .O(N__26662),
            .I(N__26648));
    InMux I__5888 (
            .O(N__26661),
            .I(N__26645));
    InMux I__5887 (
            .O(N__26660),
            .I(N__26642));
    LocalMux I__5886 (
            .O(N__26657),
            .I(N__26639));
    LocalMux I__5885 (
            .O(N__26654),
            .I(N__26636));
    InMux I__5884 (
            .O(N__26653),
            .I(N__26633));
    InMux I__5883 (
            .O(N__26652),
            .I(N__26630));
    InMux I__5882 (
            .O(N__26651),
            .I(N__26627));
    LocalMux I__5881 (
            .O(N__26648),
            .I(N__26624));
    LocalMux I__5880 (
            .O(N__26645),
            .I(N__26621));
    LocalMux I__5879 (
            .O(N__26642),
            .I(N__26618));
    Span4Mux_v I__5878 (
            .O(N__26639),
            .I(N__26613));
    Span4Mux_v I__5877 (
            .O(N__26636),
            .I(N__26613));
    LocalMux I__5876 (
            .O(N__26633),
            .I(N__26610));
    LocalMux I__5875 (
            .O(N__26630),
            .I(N__26607));
    LocalMux I__5874 (
            .O(N__26627),
            .I(N__26604));
    Span4Mux_v I__5873 (
            .O(N__26624),
            .I(N__26599));
    Span4Mux_h I__5872 (
            .O(N__26621),
            .I(N__26599));
    Span4Mux_s2_v I__5871 (
            .O(N__26618),
            .I(N__26596));
    Span4Mux_h I__5870 (
            .O(N__26613),
            .I(N__26593));
    Span12Mux_s9_h I__5869 (
            .O(N__26610),
            .I(N__26590));
    Span4Mux_h I__5868 (
            .O(N__26607),
            .I(N__26583));
    Span4Mux_v I__5867 (
            .O(N__26604),
            .I(N__26583));
    Span4Mux_v I__5866 (
            .O(N__26599),
            .I(N__26583));
    Span4Mux_h I__5865 (
            .O(N__26596),
            .I(N__26580));
    Span4Mux_h I__5864 (
            .O(N__26593),
            .I(N__26577));
    Span12Mux_v I__5863 (
            .O(N__26590),
            .I(N__26574));
    Span4Mux_h I__5862 (
            .O(N__26583),
            .I(N__26569));
    Span4Mux_v I__5861 (
            .O(N__26580),
            .I(N__26569));
    Odrv4 I__5860 (
            .O(N__26577),
            .I(N_248));
    Odrv12 I__5859 (
            .O(N__26574),
            .I(N_248));
    Odrv4 I__5858 (
            .O(N__26569),
            .I(N_248));
    InMux I__5857 (
            .O(N__26562),
            .I(N__26559));
    LocalMux I__5856 (
            .O(N__26559),
            .I(M_this_sprites_address_qc_12_0));
    InMux I__5855 (
            .O(N__26556),
            .I(N__26545));
    InMux I__5854 (
            .O(N__26555),
            .I(N__26542));
    InMux I__5853 (
            .O(N__26554),
            .I(N__26539));
    InMux I__5852 (
            .O(N__26553),
            .I(N__26533));
    CascadeMux I__5851 (
            .O(N__26552),
            .I(N__26530));
    InMux I__5850 (
            .O(N__26551),
            .I(N__26523));
    InMux I__5849 (
            .O(N__26550),
            .I(N__26523));
    InMux I__5848 (
            .O(N__26549),
            .I(N__26523));
    InMux I__5847 (
            .O(N__26548),
            .I(N__26520));
    LocalMux I__5846 (
            .O(N__26545),
            .I(N__26515));
    LocalMux I__5845 (
            .O(N__26542),
            .I(N__26510));
    LocalMux I__5844 (
            .O(N__26539),
            .I(N__26510));
    InMux I__5843 (
            .O(N__26538),
            .I(N__26506));
    InMux I__5842 (
            .O(N__26537),
            .I(N__26501));
    InMux I__5841 (
            .O(N__26536),
            .I(N__26501));
    LocalMux I__5840 (
            .O(N__26533),
            .I(N__26498));
    InMux I__5839 (
            .O(N__26530),
            .I(N__26495));
    LocalMux I__5838 (
            .O(N__26523),
            .I(N__26492));
    LocalMux I__5837 (
            .O(N__26520),
            .I(N__26489));
    InMux I__5836 (
            .O(N__26519),
            .I(N__26486));
    InMux I__5835 (
            .O(N__26518),
            .I(N__26483));
    Span4Mux_h I__5834 (
            .O(N__26515),
            .I(N__26478));
    Span4Mux_h I__5833 (
            .O(N__26510),
            .I(N__26478));
    InMux I__5832 (
            .O(N__26509),
            .I(N__26475));
    LocalMux I__5831 (
            .O(N__26506),
            .I(N__26468));
    LocalMux I__5830 (
            .O(N__26501),
            .I(N__26468));
    Span4Mux_v I__5829 (
            .O(N__26498),
            .I(N__26468));
    LocalMux I__5828 (
            .O(N__26495),
            .I(N__26463));
    Span12Mux_s10_v I__5827 (
            .O(N__26492),
            .I(N__26463));
    Span4Mux_h I__5826 (
            .O(N__26489),
            .I(N__26460));
    LocalMux I__5825 (
            .O(N__26486),
            .I(N__26457));
    LocalMux I__5824 (
            .O(N__26483),
            .I(N__26454));
    Odrv4 I__5823 (
            .O(N__26478),
            .I(\this_vga_signals.N_427_0 ));
    LocalMux I__5822 (
            .O(N__26475),
            .I(\this_vga_signals.N_427_0 ));
    Odrv4 I__5821 (
            .O(N__26468),
            .I(\this_vga_signals.N_427_0 ));
    Odrv12 I__5820 (
            .O(N__26463),
            .I(\this_vga_signals.N_427_0 ));
    Odrv4 I__5819 (
            .O(N__26460),
            .I(\this_vga_signals.N_427_0 ));
    Odrv12 I__5818 (
            .O(N__26457),
            .I(\this_vga_signals.N_427_0 ));
    Odrv4 I__5817 (
            .O(N__26454),
            .I(\this_vga_signals.N_427_0 ));
    CascadeMux I__5816 (
            .O(N__26439),
            .I(N__26426));
    InMux I__5815 (
            .O(N__26438),
            .I(N__26405));
    InMux I__5814 (
            .O(N__26437),
            .I(N__26405));
    InMux I__5813 (
            .O(N__26436),
            .I(N__26405));
    InMux I__5812 (
            .O(N__26435),
            .I(N__26398));
    InMux I__5811 (
            .O(N__26434),
            .I(N__26398));
    InMux I__5810 (
            .O(N__26433),
            .I(N__26391));
    InMux I__5809 (
            .O(N__26432),
            .I(N__26391));
    InMux I__5808 (
            .O(N__26431),
            .I(N__26391));
    InMux I__5807 (
            .O(N__26430),
            .I(N__26388));
    InMux I__5806 (
            .O(N__26429),
            .I(N__26385));
    InMux I__5805 (
            .O(N__26426),
            .I(N__26382));
    InMux I__5804 (
            .O(N__26425),
            .I(N__26377));
    InMux I__5803 (
            .O(N__26424),
            .I(N__26377));
    InMux I__5802 (
            .O(N__26423),
            .I(N__26370));
    InMux I__5801 (
            .O(N__26422),
            .I(N__26370));
    InMux I__5800 (
            .O(N__26421),
            .I(N__26370));
    InMux I__5799 (
            .O(N__26420),
            .I(N__26365));
    InMux I__5798 (
            .O(N__26419),
            .I(N__26365));
    InMux I__5797 (
            .O(N__26418),
            .I(N__26358));
    InMux I__5796 (
            .O(N__26417),
            .I(N__26358));
    InMux I__5795 (
            .O(N__26416),
            .I(N__26358));
    InMux I__5794 (
            .O(N__26415),
            .I(N__26353));
    InMux I__5793 (
            .O(N__26414),
            .I(N__26353));
    InMux I__5792 (
            .O(N__26413),
            .I(N__26348));
    InMux I__5791 (
            .O(N__26412),
            .I(N__26348));
    LocalMux I__5790 (
            .O(N__26405),
            .I(N__26345));
    InMux I__5789 (
            .O(N__26404),
            .I(N__26340));
    InMux I__5788 (
            .O(N__26403),
            .I(N__26340));
    LocalMux I__5787 (
            .O(N__26398),
            .I(N__26335));
    LocalMux I__5786 (
            .O(N__26391),
            .I(N__26335));
    LocalMux I__5785 (
            .O(N__26388),
            .I(N__26332));
    LocalMux I__5784 (
            .O(N__26385),
            .I(N__26317));
    LocalMux I__5783 (
            .O(N__26382),
            .I(N__26317));
    LocalMux I__5782 (
            .O(N__26377),
            .I(N__26317));
    LocalMux I__5781 (
            .O(N__26370),
            .I(N__26317));
    LocalMux I__5780 (
            .O(N__26365),
            .I(N__26317));
    LocalMux I__5779 (
            .O(N__26358),
            .I(N__26317));
    LocalMux I__5778 (
            .O(N__26353),
            .I(N__26317));
    LocalMux I__5777 (
            .O(N__26348),
            .I(N__26302));
    Span4Mux_v I__5776 (
            .O(N__26345),
            .I(N__26302));
    LocalMux I__5775 (
            .O(N__26340),
            .I(N__26302));
    Span4Mux_v I__5774 (
            .O(N__26335),
            .I(N__26302));
    Span4Mux_h I__5773 (
            .O(N__26332),
            .I(N__26299));
    Span4Mux_v I__5772 (
            .O(N__26317),
            .I(N__26296));
    InMux I__5771 (
            .O(N__26316),
            .I(N__26291));
    InMux I__5770 (
            .O(N__26315),
            .I(N__26291));
    InMux I__5769 (
            .O(N__26314),
            .I(N__26282));
    InMux I__5768 (
            .O(N__26313),
            .I(N__26282));
    InMux I__5767 (
            .O(N__26312),
            .I(N__26282));
    InMux I__5766 (
            .O(N__26311),
            .I(N__26282));
    Odrv4 I__5765 (
            .O(N__26302),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5764 (
            .O(N__26299),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__5763 (
            .O(N__26296),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5762 (
            .O(N__26291),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__5761 (
            .O(N__26282),
            .I(M_this_state_qZ0Z_1));
    CascadeMux I__5760 (
            .O(N__26271),
            .I(\this_vga_signals.N_427_0_cascade_ ));
    CascadeMux I__5759 (
            .O(N__26268),
            .I(N__26265));
    InMux I__5758 (
            .O(N__26265),
            .I(N__26262));
    LocalMux I__5757 (
            .O(N__26262),
            .I(N__26259));
    Span12Mux_s10_v I__5756 (
            .O(N__26259),
            .I(N__26256));
    Odrv12 I__5755 (
            .O(N__26256),
            .I(N_1274_tz_0));
    InMux I__5754 (
            .O(N__26253),
            .I(N__26250));
    LocalMux I__5753 (
            .O(N__26250),
            .I(N__26247));
    Span4Mux_h I__5752 (
            .O(N__26247),
            .I(N__26244));
    Odrv4 I__5751 (
            .O(N__26244),
            .I(M_this_sprites_address_qc_0_2));
    InMux I__5750 (
            .O(N__26241),
            .I(N__26237));
    InMux I__5749 (
            .O(N__26240),
            .I(N__26234));
    LocalMux I__5748 (
            .O(N__26237),
            .I(N__26229));
    LocalMux I__5747 (
            .O(N__26234),
            .I(N__26229));
    Span4Mux_h I__5746 (
            .O(N__26229),
            .I(N__26226));
    Odrv4 I__5745 (
            .O(N__26226),
            .I(\this_vga_signals.N_889_0 ));
    CascadeMux I__5744 (
            .O(N__26223),
            .I(\this_vga_signals.N_889_0_cascade_ ));
    CascadeMux I__5743 (
            .O(N__26220),
            .I(N__26211));
    InMux I__5742 (
            .O(N__26219),
            .I(N__26208));
    InMux I__5741 (
            .O(N__26218),
            .I(N__26199));
    InMux I__5740 (
            .O(N__26217),
            .I(N__26199));
    InMux I__5739 (
            .O(N__26216),
            .I(N__26196));
    InMux I__5738 (
            .O(N__26215),
            .I(N__26191));
    InMux I__5737 (
            .O(N__26214),
            .I(N__26191));
    InMux I__5736 (
            .O(N__26211),
            .I(N__26188));
    LocalMux I__5735 (
            .O(N__26208),
            .I(N__26185));
    InMux I__5734 (
            .O(N__26207),
            .I(N__26179));
    InMux I__5733 (
            .O(N__26206),
            .I(N__26179));
    InMux I__5732 (
            .O(N__26205),
            .I(N__26174));
    InMux I__5731 (
            .O(N__26204),
            .I(N__26174));
    LocalMux I__5730 (
            .O(N__26199),
            .I(N__26170));
    LocalMux I__5729 (
            .O(N__26196),
            .I(N__26165));
    LocalMux I__5728 (
            .O(N__26191),
            .I(N__26165));
    LocalMux I__5727 (
            .O(N__26188),
            .I(N__26162));
    Span4Mux_v I__5726 (
            .O(N__26185),
            .I(N__26159));
    InMux I__5725 (
            .O(N__26184),
            .I(N__26156));
    LocalMux I__5724 (
            .O(N__26179),
            .I(N__26151));
    LocalMux I__5723 (
            .O(N__26174),
            .I(N__26151));
    InMux I__5722 (
            .O(N__26173),
            .I(N__26148));
    Span4Mux_h I__5721 (
            .O(N__26170),
            .I(N__26143));
    Span4Mux_h I__5720 (
            .O(N__26165),
            .I(N__26143));
    Odrv4 I__5719 (
            .O(N__26162),
            .I(N_750));
    Odrv4 I__5718 (
            .O(N__26159),
            .I(N_750));
    LocalMux I__5717 (
            .O(N__26156),
            .I(N_750));
    Odrv12 I__5716 (
            .O(N__26151),
            .I(N_750));
    LocalMux I__5715 (
            .O(N__26148),
            .I(N_750));
    Odrv4 I__5714 (
            .O(N__26143),
            .I(N_750));
    CascadeMux I__5713 (
            .O(N__26130),
            .I(N__26126));
    CascadeMux I__5712 (
            .O(N__26129),
            .I(N__26120));
    InMux I__5711 (
            .O(N__26126),
            .I(N__26115));
    InMux I__5710 (
            .O(N__26125),
            .I(N__26115));
    InMux I__5709 (
            .O(N__26124),
            .I(N__26112));
    InMux I__5708 (
            .O(N__26123),
            .I(N__26107));
    InMux I__5707 (
            .O(N__26120),
            .I(N__26107));
    LocalMux I__5706 (
            .O(N__26115),
            .I(N__26102));
    LocalMux I__5705 (
            .O(N__26112),
            .I(N__26099));
    LocalMux I__5704 (
            .O(N__26107),
            .I(N__26096));
    InMux I__5703 (
            .O(N__26106),
            .I(N__26091));
    InMux I__5702 (
            .O(N__26105),
            .I(N__26091));
    Span4Mux_h I__5701 (
            .O(N__26102),
            .I(N__26086));
    Span4Mux_h I__5700 (
            .O(N__26099),
            .I(N__26086));
    Span4Mux_v I__5699 (
            .O(N__26096),
            .I(N__26083));
    LocalMux I__5698 (
            .O(N__26091),
            .I(N_762));
    Odrv4 I__5697 (
            .O(N__26086),
            .I(N_762));
    Odrv4 I__5696 (
            .O(N__26083),
            .I(N_762));
    CascadeMux I__5695 (
            .O(N__26076),
            .I(N__26073));
    InMux I__5694 (
            .O(N__26073),
            .I(N__26069));
    CascadeMux I__5693 (
            .O(N__26072),
            .I(N__26066));
    LocalMux I__5692 (
            .O(N__26069),
            .I(N__26062));
    InMux I__5691 (
            .O(N__26066),
            .I(N__26059));
    CascadeMux I__5690 (
            .O(N__26065),
            .I(N__26056));
    Span4Mux_v I__5689 (
            .O(N__26062),
            .I(N__26050));
    LocalMux I__5688 (
            .O(N__26059),
            .I(N__26050));
    InMux I__5687 (
            .O(N__26056),
            .I(N__26047));
    CascadeMux I__5686 (
            .O(N__26055),
            .I(N__26044));
    Span4Mux_h I__5685 (
            .O(N__26050),
            .I(N__26036));
    LocalMux I__5684 (
            .O(N__26047),
            .I(N__26036));
    InMux I__5683 (
            .O(N__26044),
            .I(N__26033));
    CascadeMux I__5682 (
            .O(N__26043),
            .I(N__26030));
    CascadeMux I__5681 (
            .O(N__26042),
            .I(N__26025));
    CascadeMux I__5680 (
            .O(N__26041),
            .I(N__26021));
    Span4Mux_v I__5679 (
            .O(N__26036),
            .I(N__26012));
    LocalMux I__5678 (
            .O(N__26033),
            .I(N__26012));
    InMux I__5677 (
            .O(N__26030),
            .I(N__26009));
    CascadeMux I__5676 (
            .O(N__26029),
            .I(N__26006));
    CascadeMux I__5675 (
            .O(N__26028),
            .I(N__26003));
    InMux I__5674 (
            .O(N__26025),
            .I(N__26000));
    CascadeMux I__5673 (
            .O(N__26024),
            .I(N__25997));
    InMux I__5672 (
            .O(N__26021),
            .I(N__25994));
    CascadeMux I__5671 (
            .O(N__26020),
            .I(N__25991));
    CascadeMux I__5670 (
            .O(N__26019),
            .I(N__25987));
    CascadeMux I__5669 (
            .O(N__26018),
            .I(N__25984));
    CascadeMux I__5668 (
            .O(N__26017),
            .I(N__25981));
    Span4Mux_h I__5667 (
            .O(N__26012),
            .I(N__25975));
    LocalMux I__5666 (
            .O(N__26009),
            .I(N__25975));
    InMux I__5665 (
            .O(N__26006),
            .I(N__25972));
    InMux I__5664 (
            .O(N__26003),
            .I(N__25969));
    LocalMux I__5663 (
            .O(N__26000),
            .I(N__25966));
    InMux I__5662 (
            .O(N__25997),
            .I(N__25963));
    LocalMux I__5661 (
            .O(N__25994),
            .I(N__25960));
    InMux I__5660 (
            .O(N__25991),
            .I(N__25957));
    CascadeMux I__5659 (
            .O(N__25990),
            .I(N__25954));
    InMux I__5658 (
            .O(N__25987),
            .I(N__25948));
    InMux I__5657 (
            .O(N__25984),
            .I(N__25945));
    InMux I__5656 (
            .O(N__25981),
            .I(N__25942));
    CascadeMux I__5655 (
            .O(N__25980),
            .I(N__25939));
    Span4Mux_v I__5654 (
            .O(N__25975),
            .I(N__25934));
    LocalMux I__5653 (
            .O(N__25972),
            .I(N__25934));
    LocalMux I__5652 (
            .O(N__25969),
            .I(N__25931));
    Span4Mux_v I__5651 (
            .O(N__25966),
            .I(N__25926));
    LocalMux I__5650 (
            .O(N__25963),
            .I(N__25926));
    Span4Mux_v I__5649 (
            .O(N__25960),
            .I(N__25921));
    LocalMux I__5648 (
            .O(N__25957),
            .I(N__25921));
    InMux I__5647 (
            .O(N__25954),
            .I(N__25918));
    CascadeMux I__5646 (
            .O(N__25953),
            .I(N__25915));
    InMux I__5645 (
            .O(N__25952),
            .I(N__25912));
    InMux I__5644 (
            .O(N__25951),
            .I(N__25909));
    LocalMux I__5643 (
            .O(N__25948),
            .I(N__25904));
    LocalMux I__5642 (
            .O(N__25945),
            .I(N__25904));
    LocalMux I__5641 (
            .O(N__25942),
            .I(N__25901));
    InMux I__5640 (
            .O(N__25939),
            .I(N__25898));
    Span4Mux_h I__5639 (
            .O(N__25934),
            .I(N__25895));
    Span4Mux_v I__5638 (
            .O(N__25931),
            .I(N__25890));
    Span4Mux_v I__5637 (
            .O(N__25926),
            .I(N__25890));
    Span4Mux_v I__5636 (
            .O(N__25921),
            .I(N__25885));
    LocalMux I__5635 (
            .O(N__25918),
            .I(N__25885));
    InMux I__5634 (
            .O(N__25915),
            .I(N__25882));
    LocalMux I__5633 (
            .O(N__25912),
            .I(N__25879));
    LocalMux I__5632 (
            .O(N__25909),
            .I(N__25876));
    Span12Mux_v I__5631 (
            .O(N__25904),
            .I(N__25868));
    Span12Mux_s8_v I__5630 (
            .O(N__25901),
            .I(N__25868));
    LocalMux I__5629 (
            .O(N__25898),
            .I(N__25868));
    Span4Mux_v I__5628 (
            .O(N__25895),
            .I(N__25861));
    Span4Mux_h I__5627 (
            .O(N__25890),
            .I(N__25861));
    Span4Mux_h I__5626 (
            .O(N__25885),
            .I(N__25861));
    LocalMux I__5625 (
            .O(N__25882),
            .I(N__25854));
    Span4Mux_h I__5624 (
            .O(N__25879),
            .I(N__25854));
    Span4Mux_v I__5623 (
            .O(N__25876),
            .I(N__25854));
    InMux I__5622 (
            .O(N__25875),
            .I(N__25851));
    Odrv12 I__5621 (
            .O(N__25868),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv4 I__5620 (
            .O(N__25861),
            .I(M_this_sprites_address_qZ0Z_9));
    Odrv4 I__5619 (
            .O(N__25854),
            .I(M_this_sprites_address_qZ0Z_9));
    LocalMux I__5618 (
            .O(N__25851),
            .I(M_this_sprites_address_qZ0Z_9));
    CascadeMux I__5617 (
            .O(N__25842),
            .I(N_750_cascade_));
    InMux I__5616 (
            .O(N__25839),
            .I(N__25836));
    LocalMux I__5615 (
            .O(N__25836),
            .I(M_this_sprites_address_qc_9_0));
    CascadeMux I__5614 (
            .O(N__25833),
            .I(N__25830));
    InMux I__5613 (
            .O(N__25830),
            .I(N__25825));
    InMux I__5612 (
            .O(N__25829),
            .I(N__25822));
    InMux I__5611 (
            .O(N__25828),
            .I(N__25819));
    LocalMux I__5610 (
            .O(N__25825),
            .I(N__25810));
    LocalMux I__5609 (
            .O(N__25822),
            .I(N__25810));
    LocalMux I__5608 (
            .O(N__25819),
            .I(N__25807));
    InMux I__5607 (
            .O(N__25818),
            .I(N__25804));
    InMux I__5606 (
            .O(N__25817),
            .I(N__25798));
    InMux I__5605 (
            .O(N__25816),
            .I(N__25798));
    InMux I__5604 (
            .O(N__25815),
            .I(N__25795));
    Span4Mux_v I__5603 (
            .O(N__25810),
            .I(N__25790));
    Span4Mux_h I__5602 (
            .O(N__25807),
            .I(N__25790));
    LocalMux I__5601 (
            .O(N__25804),
            .I(N__25787));
    InMux I__5600 (
            .O(N__25803),
            .I(N__25784));
    LocalMux I__5599 (
            .O(N__25798),
            .I(N__25779));
    LocalMux I__5598 (
            .O(N__25795),
            .I(N__25779));
    Span4Mux_v I__5597 (
            .O(N__25790),
            .I(N__25776));
    Span4Mux_h I__5596 (
            .O(N__25787),
            .I(N__25771));
    LocalMux I__5595 (
            .O(N__25784),
            .I(N__25771));
    Span12Mux_h I__5594 (
            .O(N__25779),
            .I(N__25768));
    Span4Mux_v I__5593 (
            .O(N__25776),
            .I(N__25765));
    Sp12to4 I__5592 (
            .O(N__25771),
            .I(N__25762));
    Odrv12 I__5591 (
            .O(N__25768),
            .I(port_address_in_0));
    Odrv4 I__5590 (
            .O(N__25765),
            .I(port_address_in_0));
    Odrv12 I__5589 (
            .O(N__25762),
            .I(port_address_in_0));
    InMux I__5588 (
            .O(N__25755),
            .I(N__25752));
    LocalMux I__5587 (
            .O(N__25752),
            .I(N__25749));
    Odrv4 I__5586 (
            .O(N__25749),
            .I(\this_vga_signals.N_648 ));
    InMux I__5585 (
            .O(N__25746),
            .I(N__25739));
    InMux I__5584 (
            .O(N__25745),
            .I(N__25736));
    InMux I__5583 (
            .O(N__25744),
            .I(N__25733));
    InMux I__5582 (
            .O(N__25743),
            .I(N__25730));
    CascadeMux I__5581 (
            .O(N__25742),
            .I(N__25727));
    LocalMux I__5580 (
            .O(N__25739),
            .I(N__25723));
    LocalMux I__5579 (
            .O(N__25736),
            .I(N__25718));
    LocalMux I__5578 (
            .O(N__25733),
            .I(N__25718));
    LocalMux I__5577 (
            .O(N__25730),
            .I(N__25715));
    InMux I__5576 (
            .O(N__25727),
            .I(N__25712));
    CascadeMux I__5575 (
            .O(N__25726),
            .I(N__25708));
    Span4Mux_v I__5574 (
            .O(N__25723),
            .I(N__25704));
    Span4Mux_v I__5573 (
            .O(N__25718),
            .I(N__25697));
    Span4Mux_v I__5572 (
            .O(N__25715),
            .I(N__25697));
    LocalMux I__5571 (
            .O(N__25712),
            .I(N__25697));
    InMux I__5570 (
            .O(N__25711),
            .I(N__25694));
    InMux I__5569 (
            .O(N__25708),
            .I(N__25689));
    InMux I__5568 (
            .O(N__25707),
            .I(N__25689));
    Span4Mux_h I__5567 (
            .O(N__25704),
            .I(N__25684));
    Span4Mux_h I__5566 (
            .O(N__25697),
            .I(N__25684));
    LocalMux I__5565 (
            .O(N__25694),
            .I(N__25679));
    LocalMux I__5564 (
            .O(N__25689),
            .I(N__25679));
    Span4Mux_h I__5563 (
            .O(N__25684),
            .I(N__25676));
    Span12Mux_h I__5562 (
            .O(N__25679),
            .I(N__25673));
    Sp12to4 I__5561 (
            .O(N__25676),
            .I(N__25670));
    Odrv12 I__5560 (
            .O(N__25673),
            .I(port_address_in_1));
    Odrv12 I__5559 (
            .O(N__25670),
            .I(port_address_in_1));
    InMux I__5558 (
            .O(N__25665),
            .I(N__25659));
    InMux I__5557 (
            .O(N__25664),
            .I(N__25655));
    InMux I__5556 (
            .O(N__25663),
            .I(N__25650));
    InMux I__5555 (
            .O(N__25662),
            .I(N__25650));
    LocalMux I__5554 (
            .O(N__25659),
            .I(N__25646));
    InMux I__5553 (
            .O(N__25658),
            .I(N__25643));
    LocalMux I__5552 (
            .O(N__25655),
            .I(N__25640));
    LocalMux I__5551 (
            .O(N__25650),
            .I(N__25637));
    InMux I__5550 (
            .O(N__25649),
            .I(N__25634));
    Span4Mux_h I__5549 (
            .O(N__25646),
            .I(N__25629));
    LocalMux I__5548 (
            .O(N__25643),
            .I(N__25629));
    Span4Mux_v I__5547 (
            .O(N__25640),
            .I(N__25622));
    Span4Mux_h I__5546 (
            .O(N__25637),
            .I(N__25622));
    LocalMux I__5545 (
            .O(N__25634),
            .I(N__25622));
    Span4Mux_h I__5544 (
            .O(N__25629),
            .I(N__25619));
    Span4Mux_h I__5543 (
            .O(N__25622),
            .I(N__25616));
    Sp12to4 I__5542 (
            .O(N__25619),
            .I(N__25613));
    Span4Mux_v I__5541 (
            .O(N__25616),
            .I(N__25610));
    Span12Mux_v I__5540 (
            .O(N__25613),
            .I(N__25607));
    Span4Mux_v I__5539 (
            .O(N__25610),
            .I(N__25604));
    Odrv12 I__5538 (
            .O(N__25607),
            .I(port_address_in_2));
    Odrv4 I__5537 (
            .O(N__25604),
            .I(port_address_in_2));
    InMux I__5536 (
            .O(N__25599),
            .I(N__25596));
    LocalMux I__5535 (
            .O(N__25596),
            .I(N__25592));
    InMux I__5534 (
            .O(N__25595),
            .I(N__25589));
    Span4Mux_v I__5533 (
            .O(N__25592),
            .I(N__25584));
    LocalMux I__5532 (
            .O(N__25589),
            .I(N__25584));
    Span4Mux_h I__5531 (
            .O(N__25584),
            .I(N__25581));
    Sp12to4 I__5530 (
            .O(N__25581),
            .I(N__25578));
    Span12Mux_v I__5529 (
            .O(N__25578),
            .I(N__25575));
    Span12Mux_v I__5528 (
            .O(N__25575),
            .I(N__25572));
    Odrv12 I__5527 (
            .O(N__25572),
            .I(port_address_in_7));
    InMux I__5526 (
            .O(N__25569),
            .I(N__25565));
    InMux I__5525 (
            .O(N__25568),
            .I(N__25562));
    LocalMux I__5524 (
            .O(N__25565),
            .I(N__25559));
    LocalMux I__5523 (
            .O(N__25562),
            .I(N__25556));
    Span4Mux_h I__5522 (
            .O(N__25559),
            .I(N__25551));
    Span4Mux_v I__5521 (
            .O(N__25556),
            .I(N__25551));
    Sp12to4 I__5520 (
            .O(N__25551),
            .I(N__25548));
    Span12Mux_h I__5519 (
            .O(N__25548),
            .I(N__25544));
    InMux I__5518 (
            .O(N__25547),
            .I(N__25541));
    Odrv12 I__5517 (
            .O(N__25544),
            .I(port_rw_in));
    LocalMux I__5516 (
            .O(N__25541),
            .I(port_rw_in));
    CascadeMux I__5515 (
            .O(N__25536),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5LZ0Z8_cascade_ ));
    InMux I__5514 (
            .O(N__25533),
            .I(N__25530));
    LocalMux I__5513 (
            .O(N__25530),
            .I(N__25527));
    Span4Mux_h I__5512 (
            .O(N__25527),
            .I(N__25524));
    Odrv4 I__5511 (
            .O(N__25524),
            .I(M_this_substate_d_0_sqmuxa));
    CascadeMux I__5510 (
            .O(N__25521),
            .I(M_this_substate_d_0_sqmuxa_cascade_));
    InMux I__5509 (
            .O(N__25518),
            .I(N__25515));
    LocalMux I__5508 (
            .O(N__25515),
            .I(N__25512));
    Span4Mux_v I__5507 (
            .O(N__25512),
            .I(N__25509));
    Odrv4 I__5506 (
            .O(N__25509),
            .I(dma_c4_1_0));
    InMux I__5505 (
            .O(N__25506),
            .I(N__25495));
    InMux I__5504 (
            .O(N__25505),
            .I(N__25492));
    InMux I__5503 (
            .O(N__25504),
            .I(N__25487));
    InMux I__5502 (
            .O(N__25503),
            .I(N__25487));
    InMux I__5501 (
            .O(N__25502),
            .I(N__25479));
    InMux I__5500 (
            .O(N__25501),
            .I(N__25476));
    InMux I__5499 (
            .O(N__25500),
            .I(N__25473));
    CascadeMux I__5498 (
            .O(N__25499),
            .I(N__25469));
    InMux I__5497 (
            .O(N__25498),
            .I(N__25465));
    LocalMux I__5496 (
            .O(N__25495),
            .I(N__25462));
    LocalMux I__5495 (
            .O(N__25492),
            .I(N__25459));
    LocalMux I__5494 (
            .O(N__25487),
            .I(N__25456));
    InMux I__5493 (
            .O(N__25486),
            .I(N__25451));
    InMux I__5492 (
            .O(N__25485),
            .I(N__25451));
    InMux I__5491 (
            .O(N__25484),
            .I(N__25448));
    InMux I__5490 (
            .O(N__25483),
            .I(N__25443));
    InMux I__5489 (
            .O(N__25482),
            .I(N__25443));
    LocalMux I__5488 (
            .O(N__25479),
            .I(N__25436));
    LocalMux I__5487 (
            .O(N__25476),
            .I(N__25436));
    LocalMux I__5486 (
            .O(N__25473),
            .I(N__25436));
    InMux I__5485 (
            .O(N__25472),
            .I(N__25433));
    InMux I__5484 (
            .O(N__25469),
            .I(N__25430));
    InMux I__5483 (
            .O(N__25468),
            .I(N__25427));
    LocalMux I__5482 (
            .O(N__25465),
            .I(N__25424));
    Span4Mux_v I__5481 (
            .O(N__25462),
            .I(N__25419));
    Span4Mux_v I__5480 (
            .O(N__25459),
            .I(N__25419));
    Span4Mux_h I__5479 (
            .O(N__25456),
            .I(N__25408));
    LocalMux I__5478 (
            .O(N__25451),
            .I(N__25408));
    LocalMux I__5477 (
            .O(N__25448),
            .I(N__25408));
    LocalMux I__5476 (
            .O(N__25443),
            .I(N__25408));
    Span4Mux_v I__5475 (
            .O(N__25436),
            .I(N__25408));
    LocalMux I__5474 (
            .O(N__25433),
            .I(N__25403));
    LocalMux I__5473 (
            .O(N__25430),
            .I(N__25403));
    LocalMux I__5472 (
            .O(N__25427),
            .I(\this_vga_signals.N_732 ));
    Odrv4 I__5471 (
            .O(N__25424),
            .I(\this_vga_signals.N_732 ));
    Odrv4 I__5470 (
            .O(N__25419),
            .I(\this_vga_signals.N_732 ));
    Odrv4 I__5469 (
            .O(N__25408),
            .I(\this_vga_signals.N_732 ));
    Odrv12 I__5468 (
            .O(N__25403),
            .I(\this_vga_signals.N_732 ));
    InMux I__5467 (
            .O(N__25392),
            .I(N__25386));
    InMux I__5466 (
            .O(N__25391),
            .I(N__25386));
    LocalMux I__5465 (
            .O(N__25386),
            .I(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0));
    CascadeMux I__5464 (
            .O(N__25383),
            .I(N_622_cascade_));
    InMux I__5463 (
            .O(N__25380),
            .I(N__25377));
    LocalMux I__5462 (
            .O(N__25377),
            .I(N_1278_tz_0));
    CascadeMux I__5461 (
            .O(N__25374),
            .I(N__25371));
    InMux I__5460 (
            .O(N__25371),
            .I(N__25368));
    LocalMux I__5459 (
            .O(N__25368),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_12 ));
    CascadeMux I__5458 (
            .O(N__25365),
            .I(N_460_0_cascade_));
    CascadeMux I__5457 (
            .O(N__25362),
            .I(N__25359));
    InMux I__5456 (
            .O(N__25359),
            .I(N__25354));
    InMux I__5455 (
            .O(N__25358),
            .I(N__25341));
    InMux I__5454 (
            .O(N__25357),
            .I(N__25341));
    LocalMux I__5453 (
            .O(N__25354),
            .I(N__25338));
    InMux I__5452 (
            .O(N__25353),
            .I(N__25329));
    InMux I__5451 (
            .O(N__25352),
            .I(N__25329));
    InMux I__5450 (
            .O(N__25351),
            .I(N__25329));
    InMux I__5449 (
            .O(N__25350),
            .I(N__25329));
    InMux I__5448 (
            .O(N__25349),
            .I(N__25320));
    InMux I__5447 (
            .O(N__25348),
            .I(N__25320));
    InMux I__5446 (
            .O(N__25347),
            .I(N__25320));
    InMux I__5445 (
            .O(N__25346),
            .I(N__25320));
    LocalMux I__5444 (
            .O(N__25341),
            .I(N__25317));
    Span4Mux_v I__5443 (
            .O(N__25338),
            .I(N__25314));
    LocalMux I__5442 (
            .O(N__25329),
            .I(N__25307));
    LocalMux I__5441 (
            .O(N__25320),
            .I(N__25307));
    Span12Mux_s5_v I__5440 (
            .O(N__25317),
            .I(N__25307));
    Span4Mux_v I__5439 (
            .O(N__25314),
            .I(N__25304));
    Odrv12 I__5438 (
            .O(N__25307),
            .I(N_560));
    Odrv4 I__5437 (
            .O(N__25304),
            .I(N_560));
    CEMux I__5436 (
            .O(N__25299),
            .I(N__25296));
    LocalMux I__5435 (
            .O(N__25296),
            .I(N__25287));
    InMux I__5434 (
            .O(N__25295),
            .I(N__25284));
    InMux I__5433 (
            .O(N__25294),
            .I(N__25281));
    InMux I__5432 (
            .O(N__25293),
            .I(N__25278));
    CEMux I__5431 (
            .O(N__25292),
            .I(N__25273));
    CascadeMux I__5430 (
            .O(N__25291),
            .I(N__25270));
    InMux I__5429 (
            .O(N__25290),
            .I(N__25267));
    Span4Mux_h I__5428 (
            .O(N__25287),
            .I(N__25259));
    LocalMux I__5427 (
            .O(N__25284),
            .I(N__25259));
    LocalMux I__5426 (
            .O(N__25281),
            .I(N__25259));
    LocalMux I__5425 (
            .O(N__25278),
            .I(N__25256));
    InMux I__5424 (
            .O(N__25277),
            .I(N__25251));
    InMux I__5423 (
            .O(N__25276),
            .I(N__25251));
    LocalMux I__5422 (
            .O(N__25273),
            .I(N__25248));
    InMux I__5421 (
            .O(N__25270),
            .I(N__25245));
    LocalMux I__5420 (
            .O(N__25267),
            .I(N__25242));
    InMux I__5419 (
            .O(N__25266),
            .I(N__25239));
    Span4Mux_v I__5418 (
            .O(N__25259),
            .I(N__25236));
    Span4Mux_v I__5417 (
            .O(N__25256),
            .I(N__25231));
    LocalMux I__5416 (
            .O(N__25251),
            .I(N__25231));
    Span4Mux_v I__5415 (
            .O(N__25248),
            .I(N__25224));
    LocalMux I__5414 (
            .O(N__25245),
            .I(N__25224));
    Span4Mux_h I__5413 (
            .O(N__25242),
            .I(N__25219));
    LocalMux I__5412 (
            .O(N__25239),
            .I(N__25219));
    Span4Mux_h I__5411 (
            .O(N__25236),
            .I(N__25214));
    Span4Mux_v I__5410 (
            .O(N__25231),
            .I(N__25214));
    InMux I__5409 (
            .O(N__25230),
            .I(N__25209));
    InMux I__5408 (
            .O(N__25229),
            .I(N__25209));
    Span4Mux_h I__5407 (
            .O(N__25224),
            .I(N__25206));
    Span4Mux_h I__5406 (
            .O(N__25219),
            .I(N__25202));
    Span4Mux_v I__5405 (
            .O(N__25214),
            .I(N__25199));
    LocalMux I__5404 (
            .O(N__25209),
            .I(N__25194));
    Sp12to4 I__5403 (
            .O(N__25206),
            .I(N__25194));
    InMux I__5402 (
            .O(N__25205),
            .I(N__25191));
    Span4Mux_v I__5401 (
            .O(N__25202),
            .I(N__25188));
    Sp12to4 I__5400 (
            .O(N__25199),
            .I(N__25183));
    Span12Mux_v I__5399 (
            .O(N__25194),
            .I(N__25183));
    LocalMux I__5398 (
            .O(N__25191),
            .I(M_this_map_ram_write_en_0));
    Odrv4 I__5397 (
            .O(N__25188),
            .I(M_this_map_ram_write_en_0));
    Odrv12 I__5396 (
            .O(N__25183),
            .I(M_this_map_ram_write_en_0));
    CascadeMux I__5395 (
            .O(N__25176),
            .I(N_888_0_cascade_));
    CascadeMux I__5394 (
            .O(N__25173),
            .I(N__25170));
    InMux I__5393 (
            .O(N__25170),
            .I(N__25167));
    LocalMux I__5392 (
            .O(N__25167),
            .I(\this_vga_signals.N_779 ));
    InMux I__5391 (
            .O(N__25164),
            .I(N__25159));
    InMux I__5390 (
            .O(N__25163),
            .I(N__25156));
    InMux I__5389 (
            .O(N__25162),
            .I(N__25150));
    LocalMux I__5388 (
            .O(N__25159),
            .I(N__25145));
    LocalMux I__5387 (
            .O(N__25156),
            .I(N__25145));
    InMux I__5386 (
            .O(N__25155),
            .I(N__25142));
    InMux I__5385 (
            .O(N__25154),
            .I(N__25137));
    InMux I__5384 (
            .O(N__25153),
            .I(N__25137));
    LocalMux I__5383 (
            .O(N__25150),
            .I(this_start_data_delay_M_last_q));
    Odrv4 I__5382 (
            .O(N__25145),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__5381 (
            .O(N__25142),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__5380 (
            .O(N__25137),
            .I(this_start_data_delay_M_last_q));
    CascadeMux I__5379 (
            .O(N__25128),
            .I(N__25123));
    CascadeMux I__5378 (
            .O(N__25127),
            .I(N__25120));
    InMux I__5377 (
            .O(N__25126),
            .I(N__25112));
    InMux I__5376 (
            .O(N__25123),
            .I(N__25112));
    InMux I__5375 (
            .O(N__25120),
            .I(N__25109));
    InMux I__5374 (
            .O(N__25119),
            .I(N__25103));
    InMux I__5373 (
            .O(N__25118),
            .I(N__25103));
    CascadeMux I__5372 (
            .O(N__25117),
            .I(N__25100));
    LocalMux I__5371 (
            .O(N__25112),
            .I(N__25095));
    LocalMux I__5370 (
            .O(N__25109),
            .I(N__25095));
    InMux I__5369 (
            .O(N__25108),
            .I(N__25092));
    LocalMux I__5368 (
            .O(N__25103),
            .I(N__25089));
    InMux I__5367 (
            .O(N__25100),
            .I(N__25086));
    Span4Mux_v I__5366 (
            .O(N__25095),
            .I(N__25083));
    LocalMux I__5365 (
            .O(N__25092),
            .I(N__25080));
    Span4Mux_h I__5364 (
            .O(N__25089),
            .I(N__25075));
    LocalMux I__5363 (
            .O(N__25086),
            .I(N__25075));
    Span4Mux_h I__5362 (
            .O(N__25083),
            .I(N__25072));
    Span4Mux_v I__5361 (
            .O(N__25080),
            .I(N__25067));
    Span4Mux_v I__5360 (
            .O(N__25075),
            .I(N__25067));
    Sp12to4 I__5359 (
            .O(N__25072),
            .I(N__25062));
    Sp12to4 I__5358 (
            .O(N__25067),
            .I(N__25062));
    Span12Mux_h I__5357 (
            .O(N__25062),
            .I(N__25059));
    Odrv12 I__5356 (
            .O(N__25059),
            .I(port_enb_c));
    InMux I__5355 (
            .O(N__25056),
            .I(N__25051));
    InMux I__5354 (
            .O(N__25055),
            .I(N__25048));
    InMux I__5353 (
            .O(N__25054),
            .I(N__25041));
    LocalMux I__5352 (
            .O(N__25051),
            .I(N__25036));
    LocalMux I__5351 (
            .O(N__25048),
            .I(N__25036));
    InMux I__5350 (
            .O(N__25047),
            .I(N__25031));
    InMux I__5349 (
            .O(N__25046),
            .I(N__25031));
    InMux I__5348 (
            .O(N__25045),
            .I(N__25026));
    InMux I__5347 (
            .O(N__25044),
            .I(N__25026));
    LocalMux I__5346 (
            .O(N__25041),
            .I(M_this_delay_clk_out_0));
    Odrv4 I__5345 (
            .O(N__25036),
            .I(M_this_delay_clk_out_0));
    LocalMux I__5344 (
            .O(N__25031),
            .I(M_this_delay_clk_out_0));
    LocalMux I__5343 (
            .O(N__25026),
            .I(M_this_delay_clk_out_0));
    IoInMux I__5342 (
            .O(N__25017),
            .I(N__25014));
    LocalMux I__5341 (
            .O(N__25014),
            .I(N__25011));
    IoSpan4Mux I__5340 (
            .O(N__25011),
            .I(N__25008));
    Span4Mux_s2_v I__5339 (
            .O(N__25008),
            .I(N__25005));
    Span4Mux_v I__5338 (
            .O(N__25005),
            .I(N__25002));
    Span4Mux_v I__5337 (
            .O(N__25002),
            .I(N__24999));
    Odrv4 I__5336 (
            .O(N__24999),
            .I(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO));
    InMux I__5335 (
            .O(N__24996),
            .I(N__24993));
    LocalMux I__5334 (
            .O(N__24993),
            .I(N__24990));
    Odrv4 I__5333 (
            .O(N__24990),
            .I(M_this_state_q_RNI0A0EZ0Z_6));
    CascadeMux I__5332 (
            .O(N__24987),
            .I(M_this_state_q_RNI244K2Z0Z_6_cascade_));
    IoInMux I__5331 (
            .O(N__24984),
            .I(N__24981));
    LocalMux I__5330 (
            .O(N__24981),
            .I(N__24976));
    InMux I__5329 (
            .O(N__24980),
            .I(N__24973));
    InMux I__5328 (
            .O(N__24979),
            .I(N__24970));
    IoSpan4Mux I__5327 (
            .O(N__24976),
            .I(N__24967));
    LocalMux I__5326 (
            .O(N__24973),
            .I(N__24964));
    LocalMux I__5325 (
            .O(N__24970),
            .I(N__24961));
    Span4Mux_s2_h I__5324 (
            .O(N__24967),
            .I(N__24958));
    Span4Mux_h I__5323 (
            .O(N__24964),
            .I(N__24955));
    Span4Mux_v I__5322 (
            .O(N__24961),
            .I(N__24952));
    Sp12to4 I__5321 (
            .O(N__24958),
            .I(N__24948));
    Span4Mux_v I__5320 (
            .O(N__24955),
            .I(N__24943));
    Span4Mux_v I__5319 (
            .O(N__24952),
            .I(N__24943));
    InMux I__5318 (
            .O(N__24951),
            .I(N__24940));
    Span12Mux_h I__5317 (
            .O(N__24948),
            .I(N__24936));
    Sp12to4 I__5316 (
            .O(N__24943),
            .I(N__24933));
    LocalMux I__5315 (
            .O(N__24940),
            .I(N__24930));
    CascadeMux I__5314 (
            .O(N__24939),
            .I(N__24927));
    Span12Mux_v I__5313 (
            .O(N__24936),
            .I(N__24922));
    Span12Mux_h I__5312 (
            .O(N__24933),
            .I(N__24922));
    Span4Mux_v I__5311 (
            .O(N__24930),
            .I(N__24919));
    InMux I__5310 (
            .O(N__24927),
            .I(N__24916));
    Odrv12 I__5309 (
            .O(N__24922),
            .I(dma_0));
    Odrv4 I__5308 (
            .O(N__24919),
            .I(dma_0));
    LocalMux I__5307 (
            .O(N__24916),
            .I(dma_0));
    InMux I__5306 (
            .O(N__24909),
            .I(N__24906));
    LocalMux I__5305 (
            .O(N__24906),
            .I(N__24903));
    Odrv4 I__5304 (
            .O(N__24903),
            .I(M_this_state_q_fastZ0Z_9));
    InMux I__5303 (
            .O(N__24900),
            .I(N__24897));
    LocalMux I__5302 (
            .O(N__24897),
            .I(N__24894));
    Span4Mux_v I__5301 (
            .O(N__24894),
            .I(N__24891));
    Odrv4 I__5300 (
            .O(N__24891),
            .I(N_861));
    CascadeMux I__5299 (
            .O(N__24888),
            .I(N_861_cascade_));
    InMux I__5298 (
            .O(N__24885),
            .I(N__24882));
    LocalMux I__5297 (
            .O(N__24882),
            .I(dma_c4_1));
    CascadeMux I__5296 (
            .O(N__24879),
            .I(N__24876));
    InMux I__5295 (
            .O(N__24876),
            .I(N__24873));
    LocalMux I__5294 (
            .O(N__24873),
            .I(this_vga_signals_un20_i_a2_4_a3_0_a4_2_1));
    InMux I__5293 (
            .O(N__24870),
            .I(N__24867));
    LocalMux I__5292 (
            .O(N__24867),
            .I(\this_ppu.un1_M_haddress_q_2_cry_7_THRU_CO ));
    CascadeMux I__5291 (
            .O(N__24864),
            .I(N__24861));
    InMux I__5290 (
            .O(N__24861),
            .I(N__24858));
    LocalMux I__5289 (
            .O(N__24858),
            .I(\this_ppu.un1_M_haddress_q_cry_7_THRU_CO ));
    InMux I__5288 (
            .O(N__24855),
            .I(bfn_20_7_0_));
    InMux I__5287 (
            .O(N__24852),
            .I(N__24849));
    LocalMux I__5286 (
            .O(N__24849),
            .I(N__24845));
    InMux I__5285 (
            .O(N__24848),
            .I(N__24842));
    Span4Mux_v I__5284 (
            .O(N__24845),
            .I(N__24839));
    LocalMux I__5283 (
            .O(N__24842),
            .I(N__24836));
    Span4Mux_v I__5282 (
            .O(N__24839),
            .I(N__24833));
    Span4Mux_v I__5281 (
            .O(N__24836),
            .I(N__24830));
    Odrv4 I__5280 (
            .O(N__24833),
            .I(\this_ppu.vscroll8 ));
    Odrv4 I__5279 (
            .O(N__24830),
            .I(\this_ppu.vscroll8 ));
    InMux I__5278 (
            .O(N__24825),
            .I(N__24822));
    LocalMux I__5277 (
            .O(N__24822),
            .I(M_this_oam_ram_read_data_i_11));
    InMux I__5276 (
            .O(N__24819),
            .I(N__24816));
    LocalMux I__5275 (
            .O(N__24816),
            .I(\this_ppu.un2_vscroll_axb_0 ));
    CascadeMux I__5274 (
            .O(N__24813),
            .I(N__24805));
    CascadeMux I__5273 (
            .O(N__24812),
            .I(N__24799));
    CascadeMux I__5272 (
            .O(N__24811),
            .I(N__24796));
    CascadeMux I__5271 (
            .O(N__24810),
            .I(N__24793));
    CascadeMux I__5270 (
            .O(N__24809),
            .I(N__24790));
    CascadeMux I__5269 (
            .O(N__24808),
            .I(N__24787));
    InMux I__5268 (
            .O(N__24805),
            .I(N__24784));
    CascadeMux I__5267 (
            .O(N__24804),
            .I(N__24781));
    CascadeMux I__5266 (
            .O(N__24803),
            .I(N__24777));
    CascadeMux I__5265 (
            .O(N__24802),
            .I(N__24769));
    InMux I__5264 (
            .O(N__24799),
            .I(N__24765));
    InMux I__5263 (
            .O(N__24796),
            .I(N__24762));
    InMux I__5262 (
            .O(N__24793),
            .I(N__24759));
    InMux I__5261 (
            .O(N__24790),
            .I(N__24756));
    InMux I__5260 (
            .O(N__24787),
            .I(N__24753));
    LocalMux I__5259 (
            .O(N__24784),
            .I(N__24750));
    InMux I__5258 (
            .O(N__24781),
            .I(N__24747));
    CascadeMux I__5257 (
            .O(N__24780),
            .I(N__24744));
    InMux I__5256 (
            .O(N__24777),
            .I(N__24741));
    CascadeMux I__5255 (
            .O(N__24776),
            .I(N__24738));
    CascadeMux I__5254 (
            .O(N__24775),
            .I(N__24735));
    CascadeMux I__5253 (
            .O(N__24774),
            .I(N__24732));
    CascadeMux I__5252 (
            .O(N__24773),
            .I(N__24729));
    CascadeMux I__5251 (
            .O(N__24772),
            .I(N__24726));
    InMux I__5250 (
            .O(N__24769),
            .I(N__24723));
    CascadeMux I__5249 (
            .O(N__24768),
            .I(N__24720));
    LocalMux I__5248 (
            .O(N__24765),
            .I(N__24711));
    LocalMux I__5247 (
            .O(N__24762),
            .I(N__24711));
    LocalMux I__5246 (
            .O(N__24759),
            .I(N__24711));
    LocalMux I__5245 (
            .O(N__24756),
            .I(N__24711));
    LocalMux I__5244 (
            .O(N__24753),
            .I(N__24708));
    Span4Mux_v I__5243 (
            .O(N__24750),
            .I(N__24703));
    LocalMux I__5242 (
            .O(N__24747),
            .I(N__24703));
    InMux I__5241 (
            .O(N__24744),
            .I(N__24700));
    LocalMux I__5240 (
            .O(N__24741),
            .I(N__24697));
    InMux I__5239 (
            .O(N__24738),
            .I(N__24694));
    InMux I__5238 (
            .O(N__24735),
            .I(N__24691));
    InMux I__5237 (
            .O(N__24732),
            .I(N__24688));
    InMux I__5236 (
            .O(N__24729),
            .I(N__24685));
    InMux I__5235 (
            .O(N__24726),
            .I(N__24682));
    LocalMux I__5234 (
            .O(N__24723),
            .I(N__24679));
    InMux I__5233 (
            .O(N__24720),
            .I(N__24676));
    Span12Mux_v I__5232 (
            .O(N__24711),
            .I(N__24673));
    Span12Mux_s5_v I__5231 (
            .O(N__24708),
            .I(N__24658));
    Sp12to4 I__5230 (
            .O(N__24703),
            .I(N__24658));
    LocalMux I__5229 (
            .O(N__24700),
            .I(N__24658));
    Sp12to4 I__5228 (
            .O(N__24697),
            .I(N__24658));
    LocalMux I__5227 (
            .O(N__24694),
            .I(N__24658));
    LocalMux I__5226 (
            .O(N__24691),
            .I(N__24658));
    LocalMux I__5225 (
            .O(N__24688),
            .I(N__24658));
    LocalMux I__5224 (
            .O(N__24685),
            .I(N__24653));
    LocalMux I__5223 (
            .O(N__24682),
            .I(N__24653));
    Span4Mux_h I__5222 (
            .O(N__24679),
            .I(N__24650));
    LocalMux I__5221 (
            .O(N__24676),
            .I(N__24647));
    Span12Mux_h I__5220 (
            .O(N__24673),
            .I(N__24644));
    Span12Mux_v I__5219 (
            .O(N__24658),
            .I(N__24639));
    Span12Mux_v I__5218 (
            .O(N__24653),
            .I(N__24639));
    Span4Mux_v I__5217 (
            .O(N__24650),
            .I(N__24634));
    Span4Mux_h I__5216 (
            .O(N__24647),
            .I(N__24634));
    Odrv12 I__5215 (
            .O(N__24644),
            .I(M_this_ppu_sprites_addr_3));
    Odrv12 I__5214 (
            .O(N__24639),
            .I(M_this_ppu_sprites_addr_3));
    Odrv4 I__5213 (
            .O(N__24634),
            .I(M_this_ppu_sprites_addr_3));
    CascadeMux I__5212 (
            .O(N__24627),
            .I(N__24624));
    InMux I__5211 (
            .O(N__24624),
            .I(N__24620));
    CascadeMux I__5210 (
            .O(N__24623),
            .I(N__24617));
    LocalMux I__5209 (
            .O(N__24620),
            .I(N__24612));
    InMux I__5208 (
            .O(N__24617),
            .I(N__24609));
    CascadeMux I__5207 (
            .O(N__24616),
            .I(N__24606));
    CascadeMux I__5206 (
            .O(N__24615),
            .I(N__24602));
    Span4Mux_v I__5205 (
            .O(N__24612),
            .I(N__24597));
    LocalMux I__5204 (
            .O(N__24609),
            .I(N__24597));
    InMux I__5203 (
            .O(N__24606),
            .I(N__24594));
    CascadeMux I__5202 (
            .O(N__24605),
            .I(N__24590));
    InMux I__5201 (
            .O(N__24602),
            .I(N__24577));
    Span4Mux_h I__5200 (
            .O(N__24597),
            .I(N__24572));
    LocalMux I__5199 (
            .O(N__24594),
            .I(N__24572));
    CascadeMux I__5198 (
            .O(N__24593),
            .I(N__24569));
    InMux I__5197 (
            .O(N__24590),
            .I(N__24566));
    CascadeMux I__5196 (
            .O(N__24589),
            .I(N__24563));
    CascadeMux I__5195 (
            .O(N__24588),
            .I(N__24560));
    CascadeMux I__5194 (
            .O(N__24587),
            .I(N__24557));
    CascadeMux I__5193 (
            .O(N__24586),
            .I(N__24554));
    CascadeMux I__5192 (
            .O(N__24585),
            .I(N__24551));
    CascadeMux I__5191 (
            .O(N__24584),
            .I(N__24548));
    CascadeMux I__5190 (
            .O(N__24583),
            .I(N__24545));
    CascadeMux I__5189 (
            .O(N__24582),
            .I(N__24542));
    CascadeMux I__5188 (
            .O(N__24581),
            .I(N__24539));
    CascadeMux I__5187 (
            .O(N__24580),
            .I(N__24536));
    LocalMux I__5186 (
            .O(N__24577),
            .I(N__24533));
    Span4Mux_v I__5185 (
            .O(N__24572),
            .I(N__24530));
    InMux I__5184 (
            .O(N__24569),
            .I(N__24527));
    LocalMux I__5183 (
            .O(N__24566),
            .I(N__24524));
    InMux I__5182 (
            .O(N__24563),
            .I(N__24521));
    InMux I__5181 (
            .O(N__24560),
            .I(N__24518));
    InMux I__5180 (
            .O(N__24557),
            .I(N__24515));
    InMux I__5179 (
            .O(N__24554),
            .I(N__24512));
    InMux I__5178 (
            .O(N__24551),
            .I(N__24509));
    InMux I__5177 (
            .O(N__24548),
            .I(N__24506));
    InMux I__5176 (
            .O(N__24545),
            .I(N__24503));
    InMux I__5175 (
            .O(N__24542),
            .I(N__24500));
    InMux I__5174 (
            .O(N__24539),
            .I(N__24497));
    InMux I__5173 (
            .O(N__24536),
            .I(N__24494));
    Span12Mux_h I__5172 (
            .O(N__24533),
            .I(N__24489));
    Sp12to4 I__5171 (
            .O(N__24530),
            .I(N__24484));
    LocalMux I__5170 (
            .O(N__24527),
            .I(N__24484));
    Span12Mux_v I__5169 (
            .O(N__24524),
            .I(N__24469));
    LocalMux I__5168 (
            .O(N__24521),
            .I(N__24469));
    LocalMux I__5167 (
            .O(N__24518),
            .I(N__24469));
    LocalMux I__5166 (
            .O(N__24515),
            .I(N__24469));
    LocalMux I__5165 (
            .O(N__24512),
            .I(N__24469));
    LocalMux I__5164 (
            .O(N__24509),
            .I(N__24469));
    LocalMux I__5163 (
            .O(N__24506),
            .I(N__24469));
    LocalMux I__5162 (
            .O(N__24503),
            .I(N__24460));
    LocalMux I__5161 (
            .O(N__24500),
            .I(N__24460));
    LocalMux I__5160 (
            .O(N__24497),
            .I(N__24460));
    LocalMux I__5159 (
            .O(N__24494),
            .I(N__24460));
    CascadeMux I__5158 (
            .O(N__24493),
            .I(N__24456));
    InMux I__5157 (
            .O(N__24492),
            .I(N__24452));
    Span12Mux_v I__5156 (
            .O(N__24489),
            .I(N__24449));
    Span12Mux_h I__5155 (
            .O(N__24484),
            .I(N__24446));
    Span12Mux_v I__5154 (
            .O(N__24469),
            .I(N__24441));
    Span12Mux_s7_v I__5153 (
            .O(N__24460),
            .I(N__24441));
    InMux I__5152 (
            .O(N__24459),
            .I(N__24438));
    InMux I__5151 (
            .O(N__24456),
            .I(N__24435));
    InMux I__5150 (
            .O(N__24455),
            .I(N__24432));
    LocalMux I__5149 (
            .O(N__24452),
            .I(N__24429));
    Odrv12 I__5148 (
            .O(N__24449),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv12 I__5147 (
            .O(N__24446),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv12 I__5146 (
            .O(N__24441),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5145 (
            .O(N__24438),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5144 (
            .O(N__24435),
            .I(M_this_sprites_address_qZ0Z_10));
    LocalMux I__5143 (
            .O(N__24432),
            .I(M_this_sprites_address_qZ0Z_10));
    Odrv4 I__5142 (
            .O(N__24429),
            .I(M_this_sprites_address_qZ0Z_10));
    InMux I__5141 (
            .O(N__24414),
            .I(N__24410));
    InMux I__5140 (
            .O(N__24413),
            .I(N__24407));
    LocalMux I__5139 (
            .O(N__24410),
            .I(N__24402));
    LocalMux I__5138 (
            .O(N__24407),
            .I(N__24402));
    Odrv4 I__5137 (
            .O(N__24402),
            .I(un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0));
    CascadeMux I__5136 (
            .O(N__24399),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_10_cascade_ ));
    InMux I__5135 (
            .O(N__24396),
            .I(N__24393));
    LocalMux I__5134 (
            .O(N__24393),
            .I(N_612));
    CascadeMux I__5133 (
            .O(N__24390),
            .I(N__24387));
    InMux I__5132 (
            .O(N__24387),
            .I(N__24384));
    LocalMux I__5131 (
            .O(N__24384),
            .I(N__24381));
    Odrv4 I__5130 (
            .O(N__24381),
            .I(\this_ppu.un1_M_haddress_q_2_4 ));
    InMux I__5129 (
            .O(N__24378),
            .I(N__24375));
    LocalMux I__5128 (
            .O(N__24375),
            .I(N_627));
    CascadeMux I__5127 (
            .O(N__24372),
            .I(N_509_0_cascade_));
    CascadeMux I__5126 (
            .O(N__24369),
            .I(N__24363));
    CascadeMux I__5125 (
            .O(N__24368),
            .I(N__24360));
    CascadeMux I__5124 (
            .O(N__24367),
            .I(N__24355));
    InMux I__5123 (
            .O(N__24366),
            .I(N__24352));
    InMux I__5122 (
            .O(N__24363),
            .I(N__24349));
    InMux I__5121 (
            .O(N__24360),
            .I(N__24346));
    InMux I__5120 (
            .O(N__24359),
            .I(N__24342));
    InMux I__5119 (
            .O(N__24358),
            .I(N__24337));
    InMux I__5118 (
            .O(N__24355),
            .I(N__24337));
    LocalMux I__5117 (
            .O(N__24352),
            .I(N__24334));
    LocalMux I__5116 (
            .O(N__24349),
            .I(N__24329));
    LocalMux I__5115 (
            .O(N__24346),
            .I(N__24329));
    InMux I__5114 (
            .O(N__24345),
            .I(N__24326));
    LocalMux I__5113 (
            .O(N__24342),
            .I(N__24323));
    LocalMux I__5112 (
            .O(N__24337),
            .I(N__24320));
    Span4Mux_h I__5111 (
            .O(N__24334),
            .I(N__24313));
    Span4Mux_v I__5110 (
            .O(N__24329),
            .I(N__24313));
    LocalMux I__5109 (
            .O(N__24326),
            .I(N__24313));
    Odrv4 I__5108 (
            .O(N__24323),
            .I(\this_vga_signals.N_415_0 ));
    Odrv4 I__5107 (
            .O(N__24320),
            .I(\this_vga_signals.N_415_0 ));
    Odrv4 I__5106 (
            .O(N__24313),
            .I(\this_vga_signals.N_415_0 ));
    InMux I__5105 (
            .O(N__24306),
            .I(N__24300));
    InMux I__5104 (
            .O(N__24305),
            .I(N__24300));
    LocalMux I__5103 (
            .O(N__24300),
            .I(N__24297));
    Odrv4 I__5102 (
            .O(N__24297),
            .I(un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0));
    InMux I__5101 (
            .O(N__24294),
            .I(N__24291));
    LocalMux I__5100 (
            .O(N__24291),
            .I(M_this_sprites_address_q_0_0_i_472));
    InMux I__5099 (
            .O(N__24288),
            .I(N__24285));
    LocalMux I__5098 (
            .O(N__24285),
            .I(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_6));
    InMux I__5097 (
            .O(N__24282),
            .I(N__24276));
    CascadeMux I__5096 (
            .O(N__24281),
            .I(N__24272));
    CascadeMux I__5095 (
            .O(N__24280),
            .I(N__24269));
    InMux I__5094 (
            .O(N__24279),
            .I(N__24265));
    LocalMux I__5093 (
            .O(N__24276),
            .I(N__24262));
    InMux I__5092 (
            .O(N__24275),
            .I(N__24259));
    InMux I__5091 (
            .O(N__24272),
            .I(N__24254));
    InMux I__5090 (
            .O(N__24269),
            .I(N__24254));
    InMux I__5089 (
            .O(N__24268),
            .I(N__24251));
    LocalMux I__5088 (
            .O(N__24265),
            .I(N_773));
    Odrv4 I__5087 (
            .O(N__24262),
            .I(N_773));
    LocalMux I__5086 (
            .O(N__24259),
            .I(N_773));
    LocalMux I__5085 (
            .O(N__24254),
            .I(N_773));
    LocalMux I__5084 (
            .O(N__24251),
            .I(N_773));
    CascadeMux I__5083 (
            .O(N__24240),
            .I(N__24229));
    CascadeMux I__5082 (
            .O(N__24239),
            .I(N__24226));
    CascadeMux I__5081 (
            .O(N__24238),
            .I(N__24219));
    CascadeMux I__5080 (
            .O(N__24237),
            .I(N__24216));
    CascadeMux I__5079 (
            .O(N__24236),
            .I(N__24213));
    CascadeMux I__5078 (
            .O(N__24235),
            .I(N__24210));
    CascadeMux I__5077 (
            .O(N__24234),
            .I(N__24207));
    CascadeMux I__5076 (
            .O(N__24233),
            .I(N__24202));
    CascadeMux I__5075 (
            .O(N__24232),
            .I(N__24199));
    InMux I__5074 (
            .O(N__24229),
            .I(N__24196));
    InMux I__5073 (
            .O(N__24226),
            .I(N__24193));
    CascadeMux I__5072 (
            .O(N__24225),
            .I(N__24190));
    CascadeMux I__5071 (
            .O(N__24224),
            .I(N__24187));
    CascadeMux I__5070 (
            .O(N__24223),
            .I(N__24184));
    CascadeMux I__5069 (
            .O(N__24222),
            .I(N__24181));
    InMux I__5068 (
            .O(N__24219),
            .I(N__24178));
    InMux I__5067 (
            .O(N__24216),
            .I(N__24175));
    InMux I__5066 (
            .O(N__24213),
            .I(N__24172));
    InMux I__5065 (
            .O(N__24210),
            .I(N__24169));
    InMux I__5064 (
            .O(N__24207),
            .I(N__24166));
    CascadeMux I__5063 (
            .O(N__24206),
            .I(N__24163));
    CascadeMux I__5062 (
            .O(N__24205),
            .I(N__24160));
    InMux I__5061 (
            .O(N__24202),
            .I(N__24157));
    InMux I__5060 (
            .O(N__24199),
            .I(N__24154));
    LocalMux I__5059 (
            .O(N__24196),
            .I(N__24150));
    LocalMux I__5058 (
            .O(N__24193),
            .I(N__24146));
    InMux I__5057 (
            .O(N__24190),
            .I(N__24143));
    InMux I__5056 (
            .O(N__24187),
            .I(N__24140));
    InMux I__5055 (
            .O(N__24184),
            .I(N__24137));
    InMux I__5054 (
            .O(N__24181),
            .I(N__24134));
    LocalMux I__5053 (
            .O(N__24178),
            .I(N__24129));
    LocalMux I__5052 (
            .O(N__24175),
            .I(N__24129));
    LocalMux I__5051 (
            .O(N__24172),
            .I(N__24126));
    LocalMux I__5050 (
            .O(N__24169),
            .I(N__24121));
    LocalMux I__5049 (
            .O(N__24166),
            .I(N__24121));
    InMux I__5048 (
            .O(N__24163),
            .I(N__24118));
    InMux I__5047 (
            .O(N__24160),
            .I(N__24115));
    LocalMux I__5046 (
            .O(N__24157),
            .I(N__24110));
    LocalMux I__5045 (
            .O(N__24154),
            .I(N__24110));
    CascadeMux I__5044 (
            .O(N__24153),
            .I(N__24105));
    Span4Mux_h I__5043 (
            .O(N__24150),
            .I(N__24102));
    CascadeMux I__5042 (
            .O(N__24149),
            .I(N__24099));
    Span4Mux_v I__5041 (
            .O(N__24146),
            .I(N__24092));
    LocalMux I__5040 (
            .O(N__24143),
            .I(N__24092));
    LocalMux I__5039 (
            .O(N__24140),
            .I(N__24092));
    LocalMux I__5038 (
            .O(N__24137),
            .I(N__24089));
    LocalMux I__5037 (
            .O(N__24134),
            .I(N__24086));
    Span4Mux_v I__5036 (
            .O(N__24129),
            .I(N__24081));
    Span4Mux_v I__5035 (
            .O(N__24126),
            .I(N__24081));
    Span4Mux_v I__5034 (
            .O(N__24121),
            .I(N__24072));
    LocalMux I__5033 (
            .O(N__24118),
            .I(N__24072));
    LocalMux I__5032 (
            .O(N__24115),
            .I(N__24072));
    Span4Mux_v I__5031 (
            .O(N__24110),
            .I(N__24072));
    CascadeMux I__5030 (
            .O(N__24109),
            .I(N__24068));
    InMux I__5029 (
            .O(N__24108),
            .I(N__24063));
    InMux I__5028 (
            .O(N__24105),
            .I(N__24063));
    Span4Mux_h I__5027 (
            .O(N__24102),
            .I(N__24060));
    InMux I__5026 (
            .O(N__24099),
            .I(N__24057));
    Sp12to4 I__5025 (
            .O(N__24092),
            .I(N__24050));
    Sp12to4 I__5024 (
            .O(N__24089),
            .I(N__24050));
    Sp12to4 I__5023 (
            .O(N__24086),
            .I(N__24050));
    Sp12to4 I__5022 (
            .O(N__24081),
            .I(N__24047));
    Sp12to4 I__5021 (
            .O(N__24072),
            .I(N__24044));
    InMux I__5020 (
            .O(N__24071),
            .I(N__24041));
    InMux I__5019 (
            .O(N__24068),
            .I(N__24038));
    LocalMux I__5018 (
            .O(N__24063),
            .I(N__24035));
    Span4Mux_h I__5017 (
            .O(N__24060),
            .I(N__24032));
    LocalMux I__5016 (
            .O(N__24057),
            .I(N__24023));
    Span12Mux_s8_v I__5015 (
            .O(N__24050),
            .I(N__24023));
    Span12Mux_h I__5014 (
            .O(N__24047),
            .I(N__24023));
    Span12Mux_v I__5013 (
            .O(N__24044),
            .I(N__24023));
    LocalMux I__5012 (
            .O(N__24041),
            .I(N__24020));
    LocalMux I__5011 (
            .O(N__24038),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv4 I__5010 (
            .O(N__24035),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv4 I__5009 (
            .O(N__24032),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv12 I__5008 (
            .O(N__24023),
            .I(M_this_sprites_address_qZ0Z_6));
    Odrv4 I__5007 (
            .O(N__24020),
            .I(M_this_sprites_address_qZ0Z_6));
    InMux I__5006 (
            .O(N__24009),
            .I(N__24006));
    LocalMux I__5005 (
            .O(N__24006),
            .I(M_this_sprites_address_qc_6_0));
    CascadeMux I__5004 (
            .O(N__24003),
            .I(N__24000));
    InMux I__5003 (
            .O(N__24000),
            .I(N__23997));
    LocalMux I__5002 (
            .O(N__23997),
            .I(N__23994));
    Odrv4 I__5001 (
            .O(N__23994),
            .I(N_1282_tz_0));
    InMux I__5000 (
            .O(N__23991),
            .I(N__23987));
    InMux I__4999 (
            .O(N__23990),
            .I(N__23984));
    LocalMux I__4998 (
            .O(N__23987),
            .I(un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0));
    LocalMux I__4997 (
            .O(N__23984),
            .I(un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0));
    CascadeMux I__4996 (
            .O(N__23979),
            .I(N_1290_tz_0_cascade_));
    InMux I__4995 (
            .O(N__23976),
            .I(N__23973));
    LocalMux I__4994 (
            .O(N__23973),
            .I(N_607));
    CascadeMux I__4993 (
            .O(N__23970),
            .I(N__23965));
    CascadeMux I__4992 (
            .O(N__23969),
            .I(N__23958));
    CascadeMux I__4991 (
            .O(N__23968),
            .I(N__23955));
    InMux I__4990 (
            .O(N__23965),
            .I(N__23951));
    CascadeMux I__4989 (
            .O(N__23964),
            .I(N__23948));
    CascadeMux I__4988 (
            .O(N__23963),
            .I(N__23943));
    CascadeMux I__4987 (
            .O(N__23962),
            .I(N__23939));
    CascadeMux I__4986 (
            .O(N__23961),
            .I(N__23934));
    InMux I__4985 (
            .O(N__23958),
            .I(N__23931));
    InMux I__4984 (
            .O(N__23955),
            .I(N__23928));
    CascadeMux I__4983 (
            .O(N__23954),
            .I(N__23925));
    LocalMux I__4982 (
            .O(N__23951),
            .I(N__23922));
    InMux I__4981 (
            .O(N__23948),
            .I(N__23919));
    CascadeMux I__4980 (
            .O(N__23947),
            .I(N__23916));
    CascadeMux I__4979 (
            .O(N__23946),
            .I(N__23913));
    InMux I__4978 (
            .O(N__23943),
            .I(N__23910));
    CascadeMux I__4977 (
            .O(N__23942),
            .I(N__23907));
    InMux I__4976 (
            .O(N__23939),
            .I(N__23903));
    CascadeMux I__4975 (
            .O(N__23938),
            .I(N__23900));
    CascadeMux I__4974 (
            .O(N__23937),
            .I(N__23897));
    InMux I__4973 (
            .O(N__23934),
            .I(N__23894));
    LocalMux I__4972 (
            .O(N__23931),
            .I(N__23890));
    LocalMux I__4971 (
            .O(N__23928),
            .I(N__23887));
    InMux I__4970 (
            .O(N__23925),
            .I(N__23884));
    Span4Mux_h I__4969 (
            .O(N__23922),
            .I(N__23880));
    LocalMux I__4968 (
            .O(N__23919),
            .I(N__23877));
    InMux I__4967 (
            .O(N__23916),
            .I(N__23874));
    InMux I__4966 (
            .O(N__23913),
            .I(N__23871));
    LocalMux I__4965 (
            .O(N__23910),
            .I(N__23868));
    InMux I__4964 (
            .O(N__23907),
            .I(N__23865));
    CascadeMux I__4963 (
            .O(N__23906),
            .I(N__23862));
    LocalMux I__4962 (
            .O(N__23903),
            .I(N__23859));
    InMux I__4961 (
            .O(N__23900),
            .I(N__23856));
    InMux I__4960 (
            .O(N__23897),
            .I(N__23853));
    LocalMux I__4959 (
            .O(N__23894),
            .I(N__23850));
    CascadeMux I__4958 (
            .O(N__23893),
            .I(N__23847));
    Span4Mux_s2_v I__4957 (
            .O(N__23890),
            .I(N__23840));
    Span4Mux_h I__4956 (
            .O(N__23887),
            .I(N__23840));
    LocalMux I__4955 (
            .O(N__23884),
            .I(N__23840));
    CascadeMux I__4954 (
            .O(N__23883),
            .I(N__23837));
    Span4Mux_v I__4953 (
            .O(N__23880),
            .I(N__23832));
    Span4Mux_h I__4952 (
            .O(N__23877),
            .I(N__23832));
    LocalMux I__4951 (
            .O(N__23874),
            .I(N__23829));
    LocalMux I__4950 (
            .O(N__23871),
            .I(N__23826));
    Span4Mux_h I__4949 (
            .O(N__23868),
            .I(N__23821));
    LocalMux I__4948 (
            .O(N__23865),
            .I(N__23821));
    InMux I__4947 (
            .O(N__23862),
            .I(N__23818));
    Span4Mux_h I__4946 (
            .O(N__23859),
            .I(N__23815));
    LocalMux I__4945 (
            .O(N__23856),
            .I(N__23812));
    LocalMux I__4944 (
            .O(N__23853),
            .I(N__23808));
    Span4Mux_v I__4943 (
            .O(N__23850),
            .I(N__23805));
    InMux I__4942 (
            .O(N__23847),
            .I(N__23802));
    Span4Mux_v I__4941 (
            .O(N__23840),
            .I(N__23799));
    InMux I__4940 (
            .O(N__23837),
            .I(N__23796));
    Span4Mux_v I__4939 (
            .O(N__23832),
            .I(N__23791));
    Span4Mux_h I__4938 (
            .O(N__23829),
            .I(N__23791));
    Span4Mux_v I__4937 (
            .O(N__23826),
            .I(N__23784));
    Span4Mux_v I__4936 (
            .O(N__23821),
            .I(N__23784));
    LocalMux I__4935 (
            .O(N__23818),
            .I(N__23784));
    Span4Mux_v I__4934 (
            .O(N__23815),
            .I(N__23777));
    Span4Mux_h I__4933 (
            .O(N__23812),
            .I(N__23777));
    InMux I__4932 (
            .O(N__23811),
            .I(N__23774));
    Span12Mux_h I__4931 (
            .O(N__23808),
            .I(N__23771));
    Sp12to4 I__4930 (
            .O(N__23805),
            .I(N__23766));
    LocalMux I__4929 (
            .O(N__23802),
            .I(N__23766));
    Sp12to4 I__4928 (
            .O(N__23799),
            .I(N__23761));
    LocalMux I__4927 (
            .O(N__23796),
            .I(N__23761));
    Span4Mux_h I__4926 (
            .O(N__23791),
            .I(N__23758));
    Span4Mux_h I__4925 (
            .O(N__23784),
            .I(N__23755));
    CascadeMux I__4924 (
            .O(N__23783),
            .I(N__23752));
    CascadeMux I__4923 (
            .O(N__23782),
            .I(N__23749));
    Span4Mux_h I__4922 (
            .O(N__23777),
            .I(N__23743));
    LocalMux I__4921 (
            .O(N__23774),
            .I(N__23743));
    Span12Mux_v I__4920 (
            .O(N__23771),
            .I(N__23740));
    Span12Mux_h I__4919 (
            .O(N__23766),
            .I(N__23735));
    Span12Mux_h I__4918 (
            .O(N__23761),
            .I(N__23735));
    Span4Mux_h I__4917 (
            .O(N__23758),
            .I(N__23730));
    Span4Mux_h I__4916 (
            .O(N__23755),
            .I(N__23730));
    InMux I__4915 (
            .O(N__23752),
            .I(N__23725));
    InMux I__4914 (
            .O(N__23749),
            .I(N__23725));
    InMux I__4913 (
            .O(N__23748),
            .I(N__23722));
    Span4Mux_h I__4912 (
            .O(N__23743),
            .I(N__23719));
    Odrv12 I__4911 (
            .O(N__23740),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv12 I__4910 (
            .O(N__23735),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv4 I__4909 (
            .O(N__23730),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__4908 (
            .O(N__23725),
            .I(M_this_sprites_address_qZ0Z_7));
    LocalMux I__4907 (
            .O(N__23722),
            .I(M_this_sprites_address_qZ0Z_7));
    Odrv4 I__4906 (
            .O(N__23719),
            .I(M_this_sprites_address_qZ0Z_7));
    InMux I__4905 (
            .O(N__23706),
            .I(N__23700));
    InMux I__4904 (
            .O(N__23705),
            .I(N__23700));
    LocalMux I__4903 (
            .O(N__23700),
            .I(N__23697));
    Span4Mux_h I__4902 (
            .O(N__23697),
            .I(N__23694));
    Odrv4 I__4901 (
            .O(N__23694),
            .I(un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0));
    InMux I__4900 (
            .O(N__23691),
            .I(un1_M_this_sprites_address_q_cry_6));
    CascadeMux I__4899 (
            .O(N__23688),
            .I(N__23684));
    CascadeMux I__4898 (
            .O(N__23687),
            .I(N__23678));
    InMux I__4897 (
            .O(N__23684),
            .I(N__23674));
    CascadeMux I__4896 (
            .O(N__23683),
            .I(N__23671));
    CascadeMux I__4895 (
            .O(N__23682),
            .I(N__23668));
    CascadeMux I__4894 (
            .O(N__23681),
            .I(N__23661));
    InMux I__4893 (
            .O(N__23678),
            .I(N__23658));
    CascadeMux I__4892 (
            .O(N__23677),
            .I(N__23655));
    LocalMux I__4891 (
            .O(N__23674),
            .I(N__23650));
    InMux I__4890 (
            .O(N__23671),
            .I(N__23647));
    InMux I__4889 (
            .O(N__23668),
            .I(N__23644));
    CascadeMux I__4888 (
            .O(N__23667),
            .I(N__23641));
    CascadeMux I__4887 (
            .O(N__23666),
            .I(N__23638));
    CascadeMux I__4886 (
            .O(N__23665),
            .I(N__23633));
    CascadeMux I__4885 (
            .O(N__23664),
            .I(N__23630));
    InMux I__4884 (
            .O(N__23661),
            .I(N__23625));
    LocalMux I__4883 (
            .O(N__23658),
            .I(N__23622));
    InMux I__4882 (
            .O(N__23655),
            .I(N__23619));
    CascadeMux I__4881 (
            .O(N__23654),
            .I(N__23616));
    CascadeMux I__4880 (
            .O(N__23653),
            .I(N__23613));
    Span4Mux_v I__4879 (
            .O(N__23650),
            .I(N__23606));
    LocalMux I__4878 (
            .O(N__23647),
            .I(N__23606));
    LocalMux I__4877 (
            .O(N__23644),
            .I(N__23606));
    InMux I__4876 (
            .O(N__23641),
            .I(N__23603));
    InMux I__4875 (
            .O(N__23638),
            .I(N__23600));
    CascadeMux I__4874 (
            .O(N__23637),
            .I(N__23597));
    CascadeMux I__4873 (
            .O(N__23636),
            .I(N__23594));
    InMux I__4872 (
            .O(N__23633),
            .I(N__23591));
    InMux I__4871 (
            .O(N__23630),
            .I(N__23588));
    CascadeMux I__4870 (
            .O(N__23629),
            .I(N__23585));
    CascadeMux I__4869 (
            .O(N__23628),
            .I(N__23582));
    LocalMux I__4868 (
            .O(N__23625),
            .I(N__23579));
    Span4Mux_h I__4867 (
            .O(N__23622),
            .I(N__23574));
    LocalMux I__4866 (
            .O(N__23619),
            .I(N__23574));
    InMux I__4865 (
            .O(N__23616),
            .I(N__23571));
    InMux I__4864 (
            .O(N__23613),
            .I(N__23568));
    Span4Mux_v I__4863 (
            .O(N__23606),
            .I(N__23561));
    LocalMux I__4862 (
            .O(N__23603),
            .I(N__23561));
    LocalMux I__4861 (
            .O(N__23600),
            .I(N__23561));
    InMux I__4860 (
            .O(N__23597),
            .I(N__23558));
    InMux I__4859 (
            .O(N__23594),
            .I(N__23555));
    LocalMux I__4858 (
            .O(N__23591),
            .I(N__23550));
    LocalMux I__4857 (
            .O(N__23588),
            .I(N__23550));
    InMux I__4856 (
            .O(N__23585),
            .I(N__23547));
    InMux I__4855 (
            .O(N__23582),
            .I(N__23544));
    Span4Mux_v I__4854 (
            .O(N__23579),
            .I(N__23537));
    Span4Mux_v I__4853 (
            .O(N__23574),
            .I(N__23537));
    LocalMux I__4852 (
            .O(N__23571),
            .I(N__23537));
    LocalMux I__4851 (
            .O(N__23568),
            .I(N__23533));
    Span4Mux_v I__4850 (
            .O(N__23561),
            .I(N__23526));
    LocalMux I__4849 (
            .O(N__23558),
            .I(N__23526));
    LocalMux I__4848 (
            .O(N__23555),
            .I(N__23526));
    Span4Mux_v I__4847 (
            .O(N__23550),
            .I(N__23519));
    LocalMux I__4846 (
            .O(N__23547),
            .I(N__23519));
    LocalMux I__4845 (
            .O(N__23544),
            .I(N__23519));
    Span4Mux_h I__4844 (
            .O(N__23537),
            .I(N__23514));
    CascadeMux I__4843 (
            .O(N__23536),
            .I(N__23511));
    Sp12to4 I__4842 (
            .O(N__23533),
            .I(N__23507));
    Span4Mux_v I__4841 (
            .O(N__23526),
            .I(N__23502));
    Span4Mux_v I__4840 (
            .O(N__23519),
            .I(N__23502));
    InMux I__4839 (
            .O(N__23518),
            .I(N__23499));
    InMux I__4838 (
            .O(N__23517),
            .I(N__23496));
    Span4Mux_h I__4837 (
            .O(N__23514),
            .I(N__23493));
    InMux I__4836 (
            .O(N__23511),
            .I(N__23490));
    InMux I__4835 (
            .O(N__23510),
            .I(N__23487));
    Span12Mux_s9_v I__4834 (
            .O(N__23507),
            .I(N__23478));
    Sp12to4 I__4833 (
            .O(N__23502),
            .I(N__23478));
    LocalMux I__4832 (
            .O(N__23499),
            .I(N__23478));
    LocalMux I__4831 (
            .O(N__23496),
            .I(N__23478));
    Odrv4 I__4830 (
            .O(N__23493),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__4829 (
            .O(N__23490),
            .I(M_this_sprites_address_qZ0Z_8));
    LocalMux I__4828 (
            .O(N__23487),
            .I(M_this_sprites_address_qZ0Z_8));
    Odrv12 I__4827 (
            .O(N__23478),
            .I(M_this_sprites_address_qZ0Z_8));
    InMux I__4826 (
            .O(N__23469),
            .I(N__23463));
    InMux I__4825 (
            .O(N__23468),
            .I(N__23463));
    LocalMux I__4824 (
            .O(N__23463),
            .I(N__23460));
    Odrv12 I__4823 (
            .O(N__23460),
            .I(un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0));
    InMux I__4822 (
            .O(N__23457),
            .I(bfn_19_23_0_));
    InMux I__4821 (
            .O(N__23454),
            .I(un1_M_this_sprites_address_q_cry_8));
    InMux I__4820 (
            .O(N__23451),
            .I(un1_M_this_sprites_address_q_cry_9));
    InMux I__4819 (
            .O(N__23448),
            .I(N__23445));
    LocalMux I__4818 (
            .O(N__23445),
            .I(N__23441));
    InMux I__4817 (
            .O(N__23444),
            .I(N__23438));
    Odrv4 I__4816 (
            .O(N__23441),
            .I(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0));
    LocalMux I__4815 (
            .O(N__23438),
            .I(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0));
    InMux I__4814 (
            .O(N__23433),
            .I(un1_M_this_sprites_address_q_cry_10));
    InMux I__4813 (
            .O(N__23430),
            .I(un1_M_this_sprites_address_q_cry_11));
    InMux I__4812 (
            .O(N__23427),
            .I(un1_M_this_sprites_address_q_cry_12));
    CascadeMux I__4811 (
            .O(N__23424),
            .I(N__23421));
    InMux I__4810 (
            .O(N__23421),
            .I(N__23418));
    LocalMux I__4809 (
            .O(N__23418),
            .I(N__23415));
    Span4Mux_v I__4808 (
            .O(N__23415),
            .I(N__23412));
    Odrv4 I__4807 (
            .O(N__23412),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_9 ));
    CascadeMux I__4806 (
            .O(N__23409),
            .I(N__23406));
    InMux I__4805 (
            .O(N__23406),
            .I(N__23403));
    LocalMux I__4804 (
            .O(N__23403),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_13 ));
    InMux I__4803 (
            .O(N__23400),
            .I(N__23396));
    InMux I__4802 (
            .O(N__23399),
            .I(N__23393));
    LocalMux I__4801 (
            .O(N__23396),
            .I(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0));
    LocalMux I__4800 (
            .O(N__23393),
            .I(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0));
    InMux I__4799 (
            .O(N__23388),
            .I(N__23385));
    LocalMux I__4798 (
            .O(N__23385),
            .I(\this_vga_signals.N_459_0 ));
    InMux I__4797 (
            .O(N__23382),
            .I(N__23378));
    CascadeMux I__4796 (
            .O(N__23381),
            .I(N__23374));
    LocalMux I__4795 (
            .O(N__23378),
            .I(N__23371));
    InMux I__4794 (
            .O(N__23377),
            .I(N__23368));
    InMux I__4793 (
            .O(N__23374),
            .I(N__23365));
    Span4Mux_v I__4792 (
            .O(N__23371),
            .I(N__23362));
    LocalMux I__4791 (
            .O(N__23368),
            .I(N_440_0));
    LocalMux I__4790 (
            .O(N__23365),
            .I(N_440_0));
    Odrv4 I__4789 (
            .O(N__23362),
            .I(N_440_0));
    CascadeMux I__4788 (
            .O(N__23355),
            .I(N__23348));
    CascadeMux I__4787 (
            .O(N__23354),
            .I(N__23345));
    CascadeMux I__4786 (
            .O(N__23353),
            .I(N__23342));
    CascadeMux I__4785 (
            .O(N__23352),
            .I(N__23338));
    CascadeMux I__4784 (
            .O(N__23351),
            .I(N__23331));
    InMux I__4783 (
            .O(N__23348),
            .I(N__23324));
    InMux I__4782 (
            .O(N__23345),
            .I(N__23321));
    InMux I__4781 (
            .O(N__23342),
            .I(N__23318));
    CascadeMux I__4780 (
            .O(N__23341),
            .I(N__23314));
    InMux I__4779 (
            .O(N__23338),
            .I(N__23311));
    CascadeMux I__4778 (
            .O(N__23337),
            .I(N__23308));
    CascadeMux I__4777 (
            .O(N__23336),
            .I(N__23304));
    CascadeMux I__4776 (
            .O(N__23335),
            .I(N__23301));
    CascadeMux I__4775 (
            .O(N__23334),
            .I(N__23298));
    InMux I__4774 (
            .O(N__23331),
            .I(N__23295));
    CascadeMux I__4773 (
            .O(N__23330),
            .I(N__23292));
    CascadeMux I__4772 (
            .O(N__23329),
            .I(N__23289));
    CascadeMux I__4771 (
            .O(N__23328),
            .I(N__23286));
    CascadeMux I__4770 (
            .O(N__23327),
            .I(N__23283));
    LocalMux I__4769 (
            .O(N__23324),
            .I(N__23280));
    LocalMux I__4768 (
            .O(N__23321),
            .I(N__23275));
    LocalMux I__4767 (
            .O(N__23318),
            .I(N__23275));
    CascadeMux I__4766 (
            .O(N__23317),
            .I(N__23272));
    InMux I__4765 (
            .O(N__23314),
            .I(N__23269));
    LocalMux I__4764 (
            .O(N__23311),
            .I(N__23266));
    InMux I__4763 (
            .O(N__23308),
            .I(N__23263));
    CascadeMux I__4762 (
            .O(N__23307),
            .I(N__23260));
    InMux I__4761 (
            .O(N__23304),
            .I(N__23257));
    InMux I__4760 (
            .O(N__23301),
            .I(N__23254));
    InMux I__4759 (
            .O(N__23298),
            .I(N__23251));
    LocalMux I__4758 (
            .O(N__23295),
            .I(N__23248));
    InMux I__4757 (
            .O(N__23292),
            .I(N__23245));
    InMux I__4756 (
            .O(N__23289),
            .I(N__23242));
    InMux I__4755 (
            .O(N__23286),
            .I(N__23239));
    InMux I__4754 (
            .O(N__23283),
            .I(N__23236));
    Span4Mux_v I__4753 (
            .O(N__23280),
            .I(N__23231));
    Span4Mux_v I__4752 (
            .O(N__23275),
            .I(N__23231));
    InMux I__4751 (
            .O(N__23272),
            .I(N__23228));
    LocalMux I__4750 (
            .O(N__23269),
            .I(N__23225));
    Span4Mux_h I__4749 (
            .O(N__23266),
            .I(N__23220));
    LocalMux I__4748 (
            .O(N__23263),
            .I(N__23220));
    InMux I__4747 (
            .O(N__23260),
            .I(N__23217));
    LocalMux I__4746 (
            .O(N__23257),
            .I(N__23210));
    LocalMux I__4745 (
            .O(N__23254),
            .I(N__23210));
    LocalMux I__4744 (
            .O(N__23251),
            .I(N__23210));
    Span12Mux_s7_h I__4743 (
            .O(N__23248),
            .I(N__23199));
    LocalMux I__4742 (
            .O(N__23245),
            .I(N__23199));
    LocalMux I__4741 (
            .O(N__23242),
            .I(N__23199));
    LocalMux I__4740 (
            .O(N__23239),
            .I(N__23199));
    LocalMux I__4739 (
            .O(N__23236),
            .I(N__23199));
    Span4Mux_h I__4738 (
            .O(N__23231),
            .I(N__23196));
    LocalMux I__4737 (
            .O(N__23228),
            .I(N__23193));
    Span4Mux_v I__4736 (
            .O(N__23225),
            .I(N__23186));
    Span4Mux_v I__4735 (
            .O(N__23220),
            .I(N__23186));
    LocalMux I__4734 (
            .O(N__23217),
            .I(N__23186));
    Span12Mux_s10_v I__4733 (
            .O(N__23210),
            .I(N__23172));
    Span12Mux_v I__4732 (
            .O(N__23199),
            .I(N__23172));
    Sp12to4 I__4731 (
            .O(N__23196),
            .I(N__23172));
    Span12Mux_h I__4730 (
            .O(N__23193),
            .I(N__23172));
    Span4Mux_h I__4729 (
            .O(N__23186),
            .I(N__23169));
    InMux I__4728 (
            .O(N__23185),
            .I(N__23166));
    InMux I__4727 (
            .O(N__23184),
            .I(N__23163));
    InMux I__4726 (
            .O(N__23183),
            .I(N__23158));
    InMux I__4725 (
            .O(N__23182),
            .I(N__23158));
    InMux I__4724 (
            .O(N__23181),
            .I(N__23155));
    Odrv12 I__4723 (
            .O(N__23172),
            .I(M_this_sprites_address_qZ0Z_0));
    Odrv4 I__4722 (
            .O(N__23169),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__4721 (
            .O(N__23166),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__4720 (
            .O(N__23163),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__4719 (
            .O(N__23158),
            .I(M_this_sprites_address_qZ0Z_0));
    LocalMux I__4718 (
            .O(N__23155),
            .I(M_this_sprites_address_qZ0Z_0));
    CascadeMux I__4717 (
            .O(N__23142),
            .I(N__23138));
    InMux I__4716 (
            .O(N__23141),
            .I(N__23135));
    InMux I__4715 (
            .O(N__23138),
            .I(N__23132));
    LocalMux I__4714 (
            .O(N__23135),
            .I(un1_M_this_state_q_6_0));
    LocalMux I__4713 (
            .O(N__23132),
            .I(un1_M_this_state_q_6_0));
    InMux I__4712 (
            .O(N__23127),
            .I(N__23124));
    LocalMux I__4711 (
            .O(N__23124),
            .I(N__23120));
    InMux I__4710 (
            .O(N__23123),
            .I(N__23117));
    Odrv4 I__4709 (
            .O(N__23120),
            .I(M_this_sprites_address_q_RNIRO0N6Z0Z_0));
    LocalMux I__4708 (
            .O(N__23117),
            .I(M_this_sprites_address_q_RNIRO0N6Z0Z_0));
    CascadeMux I__4707 (
            .O(N__23112),
            .I(N__23105));
    CascadeMux I__4706 (
            .O(N__23111),
            .I(N__23102));
    CascadeMux I__4705 (
            .O(N__23110),
            .I(N__23098));
    CascadeMux I__4704 (
            .O(N__23109),
            .I(N__23095));
    CascadeMux I__4703 (
            .O(N__23108),
            .I(N__23090));
    InMux I__4702 (
            .O(N__23105),
            .I(N__23084));
    InMux I__4701 (
            .O(N__23102),
            .I(N__23081));
    CascadeMux I__4700 (
            .O(N__23101),
            .I(N__23078));
    InMux I__4699 (
            .O(N__23098),
            .I(N__23075));
    InMux I__4698 (
            .O(N__23095),
            .I(N__23072));
    CascadeMux I__4697 (
            .O(N__23094),
            .I(N__23069));
    CascadeMux I__4696 (
            .O(N__23093),
            .I(N__23066));
    InMux I__4695 (
            .O(N__23090),
            .I(N__23062));
    CascadeMux I__4694 (
            .O(N__23089),
            .I(N__23059));
    CascadeMux I__4693 (
            .O(N__23088),
            .I(N__23056));
    CascadeMux I__4692 (
            .O(N__23087),
            .I(N__23051));
    LocalMux I__4691 (
            .O(N__23084),
            .I(N__23048));
    LocalMux I__4690 (
            .O(N__23081),
            .I(N__23045));
    InMux I__4689 (
            .O(N__23078),
            .I(N__23042));
    LocalMux I__4688 (
            .O(N__23075),
            .I(N__23039));
    LocalMux I__4687 (
            .O(N__23072),
            .I(N__23036));
    InMux I__4686 (
            .O(N__23069),
            .I(N__23033));
    InMux I__4685 (
            .O(N__23066),
            .I(N__23030));
    CascadeMux I__4684 (
            .O(N__23065),
            .I(N__23027));
    LocalMux I__4683 (
            .O(N__23062),
            .I(N__23024));
    InMux I__4682 (
            .O(N__23059),
            .I(N__23021));
    InMux I__4681 (
            .O(N__23056),
            .I(N__23018));
    CascadeMux I__4680 (
            .O(N__23055),
            .I(N__23015));
    CascadeMux I__4679 (
            .O(N__23054),
            .I(N__23012));
    InMux I__4678 (
            .O(N__23051),
            .I(N__23008));
    Span4Mux_h I__4677 (
            .O(N__23048),
            .I(N__23001));
    Span4Mux_v I__4676 (
            .O(N__23045),
            .I(N__23001));
    LocalMux I__4675 (
            .O(N__23042),
            .I(N__23001));
    Span4Mux_v I__4674 (
            .O(N__23039),
            .I(N__22994));
    Span4Mux_h I__4673 (
            .O(N__23036),
            .I(N__22994));
    LocalMux I__4672 (
            .O(N__23033),
            .I(N__22994));
    LocalMux I__4671 (
            .O(N__23030),
            .I(N__22991));
    InMux I__4670 (
            .O(N__23027),
            .I(N__22988));
    Span4Mux_s2_v I__4669 (
            .O(N__23024),
            .I(N__22981));
    LocalMux I__4668 (
            .O(N__23021),
            .I(N__22981));
    LocalMux I__4667 (
            .O(N__23018),
            .I(N__22981));
    InMux I__4666 (
            .O(N__23015),
            .I(N__22978));
    InMux I__4665 (
            .O(N__23012),
            .I(N__22975));
    CascadeMux I__4664 (
            .O(N__23011),
            .I(N__22971));
    LocalMux I__4663 (
            .O(N__23008),
            .I(N__22968));
    Span4Mux_v I__4662 (
            .O(N__23001),
            .I(N__22965));
    Span4Mux_v I__4661 (
            .O(N__22994),
            .I(N__22958));
    Span4Mux_h I__4660 (
            .O(N__22991),
            .I(N__22958));
    LocalMux I__4659 (
            .O(N__22988),
            .I(N__22958));
    Span4Mux_v I__4658 (
            .O(N__22981),
            .I(N__22951));
    LocalMux I__4657 (
            .O(N__22978),
            .I(N__22951));
    LocalMux I__4656 (
            .O(N__22975),
            .I(N__22951));
    CascadeMux I__4655 (
            .O(N__22974),
            .I(N__22948));
    InMux I__4654 (
            .O(N__22971),
            .I(N__22944));
    Span12Mux_h I__4653 (
            .O(N__22968),
            .I(N__22941));
    Sp12to4 I__4652 (
            .O(N__22965),
            .I(N__22938));
    Span4Mux_v I__4651 (
            .O(N__22958),
            .I(N__22933));
    Span4Mux_v I__4650 (
            .O(N__22951),
            .I(N__22933));
    InMux I__4649 (
            .O(N__22948),
            .I(N__22930));
    InMux I__4648 (
            .O(N__22947),
            .I(N__22927));
    LocalMux I__4647 (
            .O(N__22944),
            .I(N__22921));
    Span12Mux_v I__4646 (
            .O(N__22941),
            .I(N__22912));
    Span12Mux_h I__4645 (
            .O(N__22938),
            .I(N__22912));
    Sp12to4 I__4644 (
            .O(N__22933),
            .I(N__22912));
    LocalMux I__4643 (
            .O(N__22930),
            .I(N__22912));
    LocalMux I__4642 (
            .O(N__22927),
            .I(N__22909));
    InMux I__4641 (
            .O(N__22926),
            .I(N__22906));
    InMux I__4640 (
            .O(N__22925),
            .I(N__22903));
    InMux I__4639 (
            .O(N__22924),
            .I(N__22900));
    Odrv12 I__4638 (
            .O(N__22921),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv12 I__4637 (
            .O(N__22912),
            .I(M_this_sprites_address_qZ0Z_1));
    Odrv4 I__4636 (
            .O(N__22909),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__4635 (
            .O(N__22906),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__4634 (
            .O(N__22903),
            .I(M_this_sprites_address_qZ0Z_1));
    LocalMux I__4633 (
            .O(N__22900),
            .I(M_this_sprites_address_qZ0Z_1));
    InMux I__4632 (
            .O(N__22887),
            .I(N__22884));
    LocalMux I__4631 (
            .O(N__22884),
            .I(N__22880));
    InMux I__4630 (
            .O(N__22883),
            .I(N__22877));
    Odrv4 I__4629 (
            .O(N__22880),
            .I(un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0));
    LocalMux I__4628 (
            .O(N__22877),
            .I(un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0));
    InMux I__4627 (
            .O(N__22872),
            .I(un1_M_this_sprites_address_q_cry_0));
    CascadeMux I__4626 (
            .O(N__22869),
            .I(N__22865));
    CascadeMux I__4625 (
            .O(N__22868),
            .I(N__22860));
    InMux I__4624 (
            .O(N__22865),
            .I(N__22849));
    CascadeMux I__4623 (
            .O(N__22864),
            .I(N__22846));
    CascadeMux I__4622 (
            .O(N__22863),
            .I(N__22842));
    InMux I__4621 (
            .O(N__22860),
            .I(N__22839));
    CascadeMux I__4620 (
            .O(N__22859),
            .I(N__22836));
    CascadeMux I__4619 (
            .O(N__22858),
            .I(N__22833));
    CascadeMux I__4618 (
            .O(N__22857),
            .I(N__22830));
    CascadeMux I__4617 (
            .O(N__22856),
            .I(N__22827));
    CascadeMux I__4616 (
            .O(N__22855),
            .I(N__22824));
    CascadeMux I__4615 (
            .O(N__22854),
            .I(N__22821));
    CascadeMux I__4614 (
            .O(N__22853),
            .I(N__22818));
    CascadeMux I__4613 (
            .O(N__22852),
            .I(N__22814));
    LocalMux I__4612 (
            .O(N__22849),
            .I(N__22811));
    InMux I__4611 (
            .O(N__22846),
            .I(N__22808));
    CascadeMux I__4610 (
            .O(N__22845),
            .I(N__22805));
    InMux I__4609 (
            .O(N__22842),
            .I(N__22802));
    LocalMux I__4608 (
            .O(N__22839),
            .I(N__22797));
    InMux I__4607 (
            .O(N__22836),
            .I(N__22794));
    InMux I__4606 (
            .O(N__22833),
            .I(N__22791));
    InMux I__4605 (
            .O(N__22830),
            .I(N__22788));
    InMux I__4604 (
            .O(N__22827),
            .I(N__22785));
    InMux I__4603 (
            .O(N__22824),
            .I(N__22782));
    InMux I__4602 (
            .O(N__22821),
            .I(N__22779));
    InMux I__4601 (
            .O(N__22818),
            .I(N__22776));
    CascadeMux I__4600 (
            .O(N__22817),
            .I(N__22772));
    InMux I__4599 (
            .O(N__22814),
            .I(N__22769));
    Span4Mux_v I__4598 (
            .O(N__22811),
            .I(N__22764));
    LocalMux I__4597 (
            .O(N__22808),
            .I(N__22764));
    InMux I__4596 (
            .O(N__22805),
            .I(N__22761));
    LocalMux I__4595 (
            .O(N__22802),
            .I(N__22758));
    CascadeMux I__4594 (
            .O(N__22801),
            .I(N__22755));
    CascadeMux I__4593 (
            .O(N__22800),
            .I(N__22752));
    Span4Mux_v I__4592 (
            .O(N__22797),
            .I(N__22745));
    LocalMux I__4591 (
            .O(N__22794),
            .I(N__22745));
    LocalMux I__4590 (
            .O(N__22791),
            .I(N__22745));
    LocalMux I__4589 (
            .O(N__22788),
            .I(N__22742));
    LocalMux I__4588 (
            .O(N__22785),
            .I(N__22737));
    LocalMux I__4587 (
            .O(N__22782),
            .I(N__22737));
    LocalMux I__4586 (
            .O(N__22779),
            .I(N__22732));
    LocalMux I__4585 (
            .O(N__22776),
            .I(N__22732));
    CascadeMux I__4584 (
            .O(N__22775),
            .I(N__22729));
    InMux I__4583 (
            .O(N__22772),
            .I(N__22726));
    LocalMux I__4582 (
            .O(N__22769),
            .I(N__22719));
    Span4Mux_v I__4581 (
            .O(N__22764),
            .I(N__22719));
    LocalMux I__4580 (
            .O(N__22761),
            .I(N__22719));
    Span4Mux_v I__4579 (
            .O(N__22758),
            .I(N__22716));
    InMux I__4578 (
            .O(N__22755),
            .I(N__22713));
    InMux I__4577 (
            .O(N__22752),
            .I(N__22710));
    Span4Mux_v I__4576 (
            .O(N__22745),
            .I(N__22707));
    Span4Mux_v I__4575 (
            .O(N__22742),
            .I(N__22704));
    Span4Mux_v I__4574 (
            .O(N__22737),
            .I(N__22698));
    Span4Mux_v I__4573 (
            .O(N__22732),
            .I(N__22698));
    InMux I__4572 (
            .O(N__22729),
            .I(N__22695));
    LocalMux I__4571 (
            .O(N__22726),
            .I(N__22692));
    Span4Mux_v I__4570 (
            .O(N__22719),
            .I(N__22687));
    Span4Mux_h I__4569 (
            .O(N__22716),
            .I(N__22684));
    LocalMux I__4568 (
            .O(N__22713),
            .I(N__22681));
    LocalMux I__4567 (
            .O(N__22710),
            .I(N__22674));
    Sp12to4 I__4566 (
            .O(N__22707),
            .I(N__22674));
    Sp12to4 I__4565 (
            .O(N__22704),
            .I(N__22674));
    InMux I__4564 (
            .O(N__22703),
            .I(N__22671));
    Span4Mux_h I__4563 (
            .O(N__22698),
            .I(N__22668));
    LocalMux I__4562 (
            .O(N__22695),
            .I(N__22665));
    Span12Mux_h I__4561 (
            .O(N__22692),
            .I(N__22662));
    InMux I__4560 (
            .O(N__22691),
            .I(N__22659));
    InMux I__4559 (
            .O(N__22690),
            .I(N__22656));
    Span4Mux_h I__4558 (
            .O(N__22687),
            .I(N__22651));
    Span4Mux_v I__4557 (
            .O(N__22684),
            .I(N__22651));
    Span12Mux_h I__4556 (
            .O(N__22681),
            .I(N__22646));
    Span12Mux_h I__4555 (
            .O(N__22674),
            .I(N__22646));
    LocalMux I__4554 (
            .O(N__22671),
            .I(N__22639));
    Span4Mux_h I__4553 (
            .O(N__22668),
            .I(N__22639));
    Span4Mux_v I__4552 (
            .O(N__22665),
            .I(N__22639));
    Odrv12 I__4551 (
            .O(N__22662),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__4550 (
            .O(N__22659),
            .I(M_this_sprites_address_qZ0Z_2));
    LocalMux I__4549 (
            .O(N__22656),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv4 I__4548 (
            .O(N__22651),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv12 I__4547 (
            .O(N__22646),
            .I(M_this_sprites_address_qZ0Z_2));
    Odrv4 I__4546 (
            .O(N__22639),
            .I(M_this_sprites_address_qZ0Z_2));
    InMux I__4545 (
            .O(N__22626),
            .I(N__22620));
    InMux I__4544 (
            .O(N__22625),
            .I(N__22620));
    LocalMux I__4543 (
            .O(N__22620),
            .I(N__22617));
    Span4Mux_h I__4542 (
            .O(N__22617),
            .I(N__22614));
    Odrv4 I__4541 (
            .O(N__22614),
            .I(un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0));
    InMux I__4540 (
            .O(N__22611),
            .I(un1_M_this_sprites_address_q_cry_1));
    CascadeMux I__4539 (
            .O(N__22608),
            .I(N__22605));
    InMux I__4538 (
            .O(N__22605),
            .I(N__22599));
    CascadeMux I__4537 (
            .O(N__22604),
            .I(N__22596));
    CascadeMux I__4536 (
            .O(N__22603),
            .I(N__22593));
    CascadeMux I__4535 (
            .O(N__22602),
            .I(N__22588));
    LocalMux I__4534 (
            .O(N__22599),
            .I(N__22583));
    InMux I__4533 (
            .O(N__22596),
            .I(N__22580));
    InMux I__4532 (
            .O(N__22593),
            .I(N__22577));
    CascadeMux I__4531 (
            .O(N__22592),
            .I(N__22574));
    CascadeMux I__4530 (
            .O(N__22591),
            .I(N__22571));
    InMux I__4529 (
            .O(N__22588),
            .I(N__22566));
    CascadeMux I__4528 (
            .O(N__22587),
            .I(N__22563));
    CascadeMux I__4527 (
            .O(N__22586),
            .I(N__22560));
    Span4Mux_h I__4526 (
            .O(N__22583),
            .I(N__22549));
    LocalMux I__4525 (
            .O(N__22580),
            .I(N__22549));
    LocalMux I__4524 (
            .O(N__22577),
            .I(N__22546));
    InMux I__4523 (
            .O(N__22574),
            .I(N__22543));
    InMux I__4522 (
            .O(N__22571),
            .I(N__22540));
    CascadeMux I__4521 (
            .O(N__22570),
            .I(N__22537));
    CascadeMux I__4520 (
            .O(N__22569),
            .I(N__22534));
    LocalMux I__4519 (
            .O(N__22566),
            .I(N__22531));
    InMux I__4518 (
            .O(N__22563),
            .I(N__22528));
    InMux I__4517 (
            .O(N__22560),
            .I(N__22525));
    CascadeMux I__4516 (
            .O(N__22559),
            .I(N__22522));
    CascadeMux I__4515 (
            .O(N__22558),
            .I(N__22519));
    CascadeMux I__4514 (
            .O(N__22557),
            .I(N__22516));
    CascadeMux I__4513 (
            .O(N__22556),
            .I(N__22513));
    CascadeMux I__4512 (
            .O(N__22555),
            .I(N__22510));
    CascadeMux I__4511 (
            .O(N__22554),
            .I(N__22507));
    Span4Mux_v I__4510 (
            .O(N__22549),
            .I(N__22500));
    Span4Mux_h I__4509 (
            .O(N__22546),
            .I(N__22500));
    LocalMux I__4508 (
            .O(N__22543),
            .I(N__22500));
    LocalMux I__4507 (
            .O(N__22540),
            .I(N__22497));
    InMux I__4506 (
            .O(N__22537),
            .I(N__22494));
    InMux I__4505 (
            .O(N__22534),
            .I(N__22491));
    Span4Mux_s2_v I__4504 (
            .O(N__22531),
            .I(N__22484));
    LocalMux I__4503 (
            .O(N__22528),
            .I(N__22484));
    LocalMux I__4502 (
            .O(N__22525),
            .I(N__22484));
    InMux I__4501 (
            .O(N__22522),
            .I(N__22481));
    InMux I__4500 (
            .O(N__22519),
            .I(N__22478));
    InMux I__4499 (
            .O(N__22516),
            .I(N__22475));
    InMux I__4498 (
            .O(N__22513),
            .I(N__22472));
    InMux I__4497 (
            .O(N__22510),
            .I(N__22469));
    InMux I__4496 (
            .O(N__22507),
            .I(N__22466));
    Span4Mux_v I__4495 (
            .O(N__22500),
            .I(N__22459));
    Span4Mux_h I__4494 (
            .O(N__22497),
            .I(N__22459));
    LocalMux I__4493 (
            .O(N__22494),
            .I(N__22459));
    LocalMux I__4492 (
            .O(N__22491),
            .I(N__22456));
    Span4Mux_v I__4491 (
            .O(N__22484),
            .I(N__22449));
    LocalMux I__4490 (
            .O(N__22481),
            .I(N__22449));
    LocalMux I__4489 (
            .O(N__22478),
            .I(N__22449));
    LocalMux I__4488 (
            .O(N__22475),
            .I(N__22443));
    LocalMux I__4487 (
            .O(N__22472),
            .I(N__22443));
    LocalMux I__4486 (
            .O(N__22469),
            .I(N__22438));
    LocalMux I__4485 (
            .O(N__22466),
            .I(N__22438));
    Span4Mux_v I__4484 (
            .O(N__22459),
            .I(N__22431));
    Span4Mux_h I__4483 (
            .O(N__22456),
            .I(N__22431));
    Span4Mux_v I__4482 (
            .O(N__22449),
            .I(N__22431));
    InMux I__4481 (
            .O(N__22448),
            .I(N__22428));
    Span4Mux_v I__4480 (
            .O(N__22443),
            .I(N__22423));
    Span4Mux_v I__4479 (
            .O(N__22438),
            .I(N__22423));
    Span4Mux_h I__4478 (
            .O(N__22431),
            .I(N__22415));
    LocalMux I__4477 (
            .O(N__22428),
            .I(N__22415));
    Sp12to4 I__4476 (
            .O(N__22423),
            .I(N__22412));
    InMux I__4475 (
            .O(N__22422),
            .I(N__22407));
    InMux I__4474 (
            .O(N__22421),
            .I(N__22407));
    InMux I__4473 (
            .O(N__22420),
            .I(N__22404));
    Span4Mux_h I__4472 (
            .O(N__22415),
            .I(N__22401));
    Odrv12 I__4471 (
            .O(N__22412),
            .I(M_this_sprites_address_qZ0Z_3));
    LocalMux I__4470 (
            .O(N__22407),
            .I(M_this_sprites_address_qZ0Z_3));
    LocalMux I__4469 (
            .O(N__22404),
            .I(M_this_sprites_address_qZ0Z_3));
    Odrv4 I__4468 (
            .O(N__22401),
            .I(M_this_sprites_address_qZ0Z_3));
    CascadeMux I__4467 (
            .O(N__22392),
            .I(N__22389));
    InMux I__4466 (
            .O(N__22389),
            .I(N__22386));
    LocalMux I__4465 (
            .O(N__22386),
            .I(N__22382));
    InMux I__4464 (
            .O(N__22385),
            .I(N__22379));
    Span4Mux_h I__4463 (
            .O(N__22382),
            .I(N__22376));
    LocalMux I__4462 (
            .O(N__22379),
            .I(un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0));
    Odrv4 I__4461 (
            .O(N__22376),
            .I(un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0));
    InMux I__4460 (
            .O(N__22371),
            .I(un1_M_this_sprites_address_q_cry_2));
    CascadeMux I__4459 (
            .O(N__22368),
            .I(N__22362));
    CascadeMux I__4458 (
            .O(N__22367),
            .I(N__22359));
    CascadeMux I__4457 (
            .O(N__22366),
            .I(N__22353));
    CascadeMux I__4456 (
            .O(N__22365),
            .I(N__22349));
    InMux I__4455 (
            .O(N__22362),
            .I(N__22342));
    InMux I__4454 (
            .O(N__22359),
            .I(N__22339));
    CascadeMux I__4453 (
            .O(N__22358),
            .I(N__22336));
    CascadeMux I__4452 (
            .O(N__22357),
            .I(N__22331));
    CascadeMux I__4451 (
            .O(N__22356),
            .I(N__22328));
    InMux I__4450 (
            .O(N__22353),
            .I(N__22325));
    CascadeMux I__4449 (
            .O(N__22352),
            .I(N__22322));
    InMux I__4448 (
            .O(N__22349),
            .I(N__22319));
    CascadeMux I__4447 (
            .O(N__22348),
            .I(N__22316));
    CascadeMux I__4446 (
            .O(N__22347),
            .I(N__22313));
    CascadeMux I__4445 (
            .O(N__22346),
            .I(N__22310));
    CascadeMux I__4444 (
            .O(N__22345),
            .I(N__22306));
    LocalMux I__4443 (
            .O(N__22342),
            .I(N__22301));
    LocalMux I__4442 (
            .O(N__22339),
            .I(N__22301));
    InMux I__4441 (
            .O(N__22336),
            .I(N__22298));
    CascadeMux I__4440 (
            .O(N__22335),
            .I(N__22295));
    CascadeMux I__4439 (
            .O(N__22334),
            .I(N__22292));
    InMux I__4438 (
            .O(N__22331),
            .I(N__22289));
    InMux I__4437 (
            .O(N__22328),
            .I(N__22286));
    LocalMux I__4436 (
            .O(N__22325),
            .I(N__22283));
    InMux I__4435 (
            .O(N__22322),
            .I(N__22280));
    LocalMux I__4434 (
            .O(N__22319),
            .I(N__22276));
    InMux I__4433 (
            .O(N__22316),
            .I(N__22273));
    InMux I__4432 (
            .O(N__22313),
            .I(N__22270));
    InMux I__4431 (
            .O(N__22310),
            .I(N__22267));
    CascadeMux I__4430 (
            .O(N__22309),
            .I(N__22264));
    InMux I__4429 (
            .O(N__22306),
            .I(N__22261));
    Span4Mux_v I__4428 (
            .O(N__22301),
            .I(N__22256));
    LocalMux I__4427 (
            .O(N__22298),
            .I(N__22256));
    InMux I__4426 (
            .O(N__22295),
            .I(N__22253));
    InMux I__4425 (
            .O(N__22292),
            .I(N__22250));
    LocalMux I__4424 (
            .O(N__22289),
            .I(N__22247));
    LocalMux I__4423 (
            .O(N__22286),
            .I(N__22242));
    Span4Mux_h I__4422 (
            .O(N__22283),
            .I(N__22242));
    LocalMux I__4421 (
            .O(N__22280),
            .I(N__22239));
    CascadeMux I__4420 (
            .O(N__22279),
            .I(N__22236));
    Span4Mux_v I__4419 (
            .O(N__22276),
            .I(N__22231));
    LocalMux I__4418 (
            .O(N__22273),
            .I(N__22231));
    LocalMux I__4417 (
            .O(N__22270),
            .I(N__22226));
    LocalMux I__4416 (
            .O(N__22267),
            .I(N__22226));
    InMux I__4415 (
            .O(N__22264),
            .I(N__22223));
    LocalMux I__4414 (
            .O(N__22261),
            .I(N__22220));
    Span4Mux_h I__4413 (
            .O(N__22256),
            .I(N__22217));
    LocalMux I__4412 (
            .O(N__22253),
            .I(N__22212));
    LocalMux I__4411 (
            .O(N__22250),
            .I(N__22212));
    Span4Mux_v I__4410 (
            .O(N__22247),
            .I(N__22205));
    Span4Mux_v I__4409 (
            .O(N__22242),
            .I(N__22205));
    Span4Mux_h I__4408 (
            .O(N__22239),
            .I(N__22205));
    InMux I__4407 (
            .O(N__22236),
            .I(N__22199));
    Span4Mux_s2_v I__4406 (
            .O(N__22231),
            .I(N__22196));
    Span4Mux_v I__4405 (
            .O(N__22226),
            .I(N__22189));
    LocalMux I__4404 (
            .O(N__22223),
            .I(N__22189));
    Span4Mux_v I__4403 (
            .O(N__22220),
            .I(N__22189));
    Span4Mux_v I__4402 (
            .O(N__22217),
            .I(N__22186));
    Span4Mux_v I__4401 (
            .O(N__22212),
            .I(N__22183));
    Span4Mux_h I__4400 (
            .O(N__22205),
            .I(N__22180));
    InMux I__4399 (
            .O(N__22204),
            .I(N__22177));
    CascadeMux I__4398 (
            .O(N__22203),
            .I(N__22174));
    CascadeMux I__4397 (
            .O(N__22202),
            .I(N__22171));
    LocalMux I__4396 (
            .O(N__22199),
            .I(N__22165));
    Sp12to4 I__4395 (
            .O(N__22196),
            .I(N__22165));
    Span4Mux_h I__4394 (
            .O(N__22189),
            .I(N__22160));
    Span4Mux_v I__4393 (
            .O(N__22186),
            .I(N__22160));
    Span4Mux_h I__4392 (
            .O(N__22183),
            .I(N__22153));
    Span4Mux_h I__4391 (
            .O(N__22180),
            .I(N__22153));
    LocalMux I__4390 (
            .O(N__22177),
            .I(N__22153));
    InMux I__4389 (
            .O(N__22174),
            .I(N__22146));
    InMux I__4388 (
            .O(N__22171),
            .I(N__22146));
    InMux I__4387 (
            .O(N__22170),
            .I(N__22146));
    Span12Mux_h I__4386 (
            .O(N__22165),
            .I(N__22143));
    Span4Mux_h I__4385 (
            .O(N__22160),
            .I(N__22140));
    Span4Mux_h I__4384 (
            .O(N__22153),
            .I(N__22137));
    LocalMux I__4383 (
            .O(N__22146),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv12 I__4382 (
            .O(N__22143),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv4 I__4381 (
            .O(N__22140),
            .I(M_this_sprites_address_qZ0Z_4));
    Odrv4 I__4380 (
            .O(N__22137),
            .I(M_this_sprites_address_qZ0Z_4));
    InMux I__4379 (
            .O(N__22128),
            .I(N__22122));
    InMux I__4378 (
            .O(N__22127),
            .I(N__22122));
    LocalMux I__4377 (
            .O(N__22122),
            .I(N__22119));
    Span4Mux_h I__4376 (
            .O(N__22119),
            .I(N__22116));
    Odrv4 I__4375 (
            .O(N__22116),
            .I(un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0));
    InMux I__4374 (
            .O(N__22113),
            .I(un1_M_this_sprites_address_q_cry_3));
    CascadeMux I__4373 (
            .O(N__22110),
            .I(N__22107));
    InMux I__4372 (
            .O(N__22107),
            .I(N__22103));
    CascadeMux I__4371 (
            .O(N__22106),
            .I(N__22100));
    LocalMux I__4370 (
            .O(N__22103),
            .I(N__22095));
    InMux I__4369 (
            .O(N__22100),
            .I(N__22092));
    CascadeMux I__4368 (
            .O(N__22099),
            .I(N__22089));
    CascadeMux I__4367 (
            .O(N__22098),
            .I(N__22085));
    Span4Mux_h I__4366 (
            .O(N__22095),
            .I(N__22078));
    LocalMux I__4365 (
            .O(N__22092),
            .I(N__22078));
    InMux I__4364 (
            .O(N__22089),
            .I(N__22075));
    CascadeMux I__4363 (
            .O(N__22088),
            .I(N__22072));
    InMux I__4362 (
            .O(N__22085),
            .I(N__22067));
    CascadeMux I__4361 (
            .O(N__22084),
            .I(N__22064));
    CascadeMux I__4360 (
            .O(N__22083),
            .I(N__22061));
    Span4Mux_v I__4359 (
            .O(N__22078),
            .I(N__22054));
    LocalMux I__4358 (
            .O(N__22075),
            .I(N__22054));
    InMux I__4357 (
            .O(N__22072),
            .I(N__22051));
    CascadeMux I__4356 (
            .O(N__22071),
            .I(N__22048));
    CascadeMux I__4355 (
            .O(N__22070),
            .I(N__22043));
    LocalMux I__4354 (
            .O(N__22067),
            .I(N__22038));
    InMux I__4353 (
            .O(N__22064),
            .I(N__22035));
    InMux I__4352 (
            .O(N__22061),
            .I(N__22032));
    CascadeMux I__4351 (
            .O(N__22060),
            .I(N__22029));
    CascadeMux I__4350 (
            .O(N__22059),
            .I(N__22026));
    Span4Mux_h I__4349 (
            .O(N__22054),
            .I(N__22021));
    LocalMux I__4348 (
            .O(N__22051),
            .I(N__22021));
    InMux I__4347 (
            .O(N__22048),
            .I(N__22018));
    CascadeMux I__4346 (
            .O(N__22047),
            .I(N__22015));
    CascadeMux I__4345 (
            .O(N__22046),
            .I(N__22011));
    InMux I__4344 (
            .O(N__22043),
            .I(N__22008));
    CascadeMux I__4343 (
            .O(N__22042),
            .I(N__22005));
    CascadeMux I__4342 (
            .O(N__22041),
            .I(N__22002));
    Span4Mux_s2_v I__4341 (
            .O(N__22038),
            .I(N__21997));
    LocalMux I__4340 (
            .O(N__22035),
            .I(N__21997));
    LocalMux I__4339 (
            .O(N__22032),
            .I(N__21994));
    InMux I__4338 (
            .O(N__22029),
            .I(N__21991));
    InMux I__4337 (
            .O(N__22026),
            .I(N__21988));
    Span4Mux_v I__4336 (
            .O(N__22021),
            .I(N__21983));
    LocalMux I__4335 (
            .O(N__22018),
            .I(N__21983));
    InMux I__4334 (
            .O(N__22015),
            .I(N__21980));
    CascadeMux I__4333 (
            .O(N__22014),
            .I(N__21977));
    InMux I__4332 (
            .O(N__22011),
            .I(N__21974));
    LocalMux I__4331 (
            .O(N__22008),
            .I(N__21971));
    InMux I__4330 (
            .O(N__22005),
            .I(N__21968));
    InMux I__4329 (
            .O(N__22002),
            .I(N__21965));
    Span4Mux_v I__4328 (
            .O(N__21997),
            .I(N__21956));
    Span4Mux_v I__4327 (
            .O(N__21994),
            .I(N__21956));
    LocalMux I__4326 (
            .O(N__21991),
            .I(N__21956));
    LocalMux I__4325 (
            .O(N__21988),
            .I(N__21956));
    Span4Mux_h I__4324 (
            .O(N__21983),
            .I(N__21951));
    LocalMux I__4323 (
            .O(N__21980),
            .I(N__21951));
    InMux I__4322 (
            .O(N__21977),
            .I(N__21948));
    LocalMux I__4321 (
            .O(N__21974),
            .I(N__21944));
    Span4Mux_v I__4320 (
            .O(N__21971),
            .I(N__21937));
    LocalMux I__4319 (
            .O(N__21968),
            .I(N__21937));
    LocalMux I__4318 (
            .O(N__21965),
            .I(N__21937));
    Span4Mux_v I__4317 (
            .O(N__21956),
            .I(N__21928));
    Span4Mux_v I__4316 (
            .O(N__21951),
            .I(N__21928));
    LocalMux I__4315 (
            .O(N__21948),
            .I(N__21928));
    InMux I__4314 (
            .O(N__21947),
            .I(N__21925));
    Span4Mux_v I__4313 (
            .O(N__21944),
            .I(N__21920));
    Span4Mux_v I__4312 (
            .O(N__21937),
            .I(N__21920));
    CascadeMux I__4311 (
            .O(N__21936),
            .I(N__21916));
    InMux I__4310 (
            .O(N__21935),
            .I(N__21913));
    Span4Mux_h I__4309 (
            .O(N__21928),
            .I(N__21908));
    LocalMux I__4308 (
            .O(N__21925),
            .I(N__21908));
    Sp12to4 I__4307 (
            .O(N__21920),
            .I(N__21905));
    InMux I__4306 (
            .O(N__21919),
            .I(N__21902));
    InMux I__4305 (
            .O(N__21916),
            .I(N__21899));
    LocalMux I__4304 (
            .O(N__21913),
            .I(N__21894));
    Span4Mux_h I__4303 (
            .O(N__21908),
            .I(N__21894));
    Odrv12 I__4302 (
            .O(N__21905),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__4301 (
            .O(N__21902),
            .I(M_this_sprites_address_qZ0Z_5));
    LocalMux I__4300 (
            .O(N__21899),
            .I(M_this_sprites_address_qZ0Z_5));
    Odrv4 I__4299 (
            .O(N__21894),
            .I(M_this_sprites_address_qZ0Z_5));
    InMux I__4298 (
            .O(N__21885),
            .I(N__21879));
    InMux I__4297 (
            .O(N__21884),
            .I(N__21879));
    LocalMux I__4296 (
            .O(N__21879),
            .I(un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0));
    InMux I__4295 (
            .O(N__21876),
            .I(un1_M_this_sprites_address_q_cry_4));
    InMux I__4294 (
            .O(N__21873),
            .I(un1_M_this_sprites_address_q_cry_5));
    InMux I__4293 (
            .O(N__21870),
            .I(N__21867));
    LocalMux I__4292 (
            .O(N__21867),
            .I(N__21864));
    Odrv4 I__4291 (
            .O(N__21864),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    InMux I__4290 (
            .O(N__21861),
            .I(N__21858));
    LocalMux I__4289 (
            .O(N__21858),
            .I(N__21855));
    Span4Mux_h I__4288 (
            .O(N__21855),
            .I(N__21852));
    Span4Mux_h I__4287 (
            .O(N__21852),
            .I(N__21849));
    Odrv4 I__4286 (
            .O(N__21849),
            .I(\this_sprites_ram.mem_out_bus6_3 ));
    InMux I__4285 (
            .O(N__21846),
            .I(N__21843));
    LocalMux I__4284 (
            .O(N__21843),
            .I(N__21840));
    Span4Mux_v I__4283 (
            .O(N__21840),
            .I(N__21837));
    Sp12to4 I__4282 (
            .O(N__21837),
            .I(N__21834));
    Odrv12 I__4281 (
            .O(N__21834),
            .I(\this_sprites_ram.mem_out_bus2_3 ));
    InMux I__4280 (
            .O(N__21831),
            .I(N__21828));
    LocalMux I__4279 (
            .O(N__21828),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ));
    CascadeMux I__4278 (
            .O(N__21825),
            .I(\this_vga_signals.N_746_cascade_ ));
    InMux I__4277 (
            .O(N__21822),
            .I(N__21819));
    LocalMux I__4276 (
            .O(N__21819),
            .I(\this_vga_signals.N_505 ));
    CascadeMux I__4275 (
            .O(N__21816),
            .I(N__21813));
    InMux I__4274 (
            .O(N__21813),
            .I(N__21810));
    LocalMux I__4273 (
            .O(N__21810),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_i_a4_2Z0Z_0 ));
    InMux I__4272 (
            .O(N__21807),
            .I(N__21804));
    LocalMux I__4271 (
            .O(N__21804),
            .I(N__21801));
    Span4Mux_h I__4270 (
            .O(N__21801),
            .I(N__21798));
    Span4Mux_h I__4269 (
            .O(N__21798),
            .I(N__21795));
    Sp12to4 I__4268 (
            .O(N__21795),
            .I(N__21792));
    Odrv12 I__4267 (
            .O(N__21792),
            .I(\this_sprites_ram.mem_out_bus4_1 ));
    InMux I__4266 (
            .O(N__21789),
            .I(N__21786));
    LocalMux I__4265 (
            .O(N__21786),
            .I(N__21783));
    Span4Mux_h I__4264 (
            .O(N__21783),
            .I(N__21780));
    Sp12to4 I__4263 (
            .O(N__21780),
            .I(N__21777));
    Span12Mux_v I__4262 (
            .O(N__21777),
            .I(N__21774));
    Odrv12 I__4261 (
            .O(N__21774),
            .I(\this_sprites_ram.mem_out_bus0_1 ));
    CascadeMux I__4260 (
            .O(N__21771),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_ ));
    InMux I__4259 (
            .O(N__21768),
            .I(N__21758));
    InMux I__4258 (
            .O(N__21767),
            .I(N__21758));
    CascadeMux I__4257 (
            .O(N__21766),
            .I(N__21754));
    InMux I__4256 (
            .O(N__21765),
            .I(N__21750));
    InMux I__4255 (
            .O(N__21764),
            .I(N__21745));
    InMux I__4254 (
            .O(N__21763),
            .I(N__21745));
    LocalMux I__4253 (
            .O(N__21758),
            .I(N__21742));
    InMux I__4252 (
            .O(N__21757),
            .I(N__21739));
    InMux I__4251 (
            .O(N__21754),
            .I(N__21734));
    InMux I__4250 (
            .O(N__21753),
            .I(N__21734));
    LocalMux I__4249 (
            .O(N__21750),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    LocalMux I__4248 (
            .O(N__21745),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    Odrv4 I__4247 (
            .O(N__21742),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    LocalMux I__4246 (
            .O(N__21739),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    LocalMux I__4245 (
            .O(N__21734),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    CascadeMux I__4244 (
            .O(N__21723),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ));
    InMux I__4243 (
            .O(N__21720),
            .I(N__21717));
    LocalMux I__4242 (
            .O(N__21717),
            .I(N__21713));
    InMux I__4241 (
            .O(N__21716),
            .I(N__21710));
    Span12Mux_h I__4240 (
            .O(N__21713),
            .I(N__21707));
    LocalMux I__4239 (
            .O(N__21710),
            .I(N__21704));
    Odrv12 I__4238 (
            .O(N__21707),
            .I(M_this_ppu_vram_data_1));
    Odrv4 I__4237 (
            .O(N__21704),
            .I(M_this_ppu_vram_data_1));
    InMux I__4236 (
            .O(N__21699),
            .I(N__21696));
    LocalMux I__4235 (
            .O(N__21696),
            .I(N__21693));
    Span12Mux_h I__4234 (
            .O(N__21693),
            .I(N__21690));
    Span12Mux_v I__4233 (
            .O(N__21690),
            .I(N__21687));
    Odrv12 I__4232 (
            .O(N__21687),
            .I(M_this_oam_ram_read_data_6));
    InMux I__4231 (
            .O(N__21684),
            .I(N__21681));
    LocalMux I__4230 (
            .O(N__21681),
            .I(N__21678));
    Sp12to4 I__4229 (
            .O(N__21678),
            .I(N__21675));
    Span12Mux_v I__4228 (
            .O(N__21675),
            .I(N__21672));
    Span12Mux_h I__4227 (
            .O(N__21672),
            .I(N__21669));
    Odrv12 I__4226 (
            .O(N__21669),
            .I(M_this_map_ram_read_data_6));
    CascadeMux I__4225 (
            .O(N__21666),
            .I(N__21663));
    InMux I__4224 (
            .O(N__21663),
            .I(N__21657));
    InMux I__4223 (
            .O(N__21662),
            .I(N__21654));
    InMux I__4222 (
            .O(N__21661),
            .I(N__21651));
    InMux I__4221 (
            .O(N__21660),
            .I(N__21648));
    LocalMux I__4220 (
            .O(N__21657),
            .I(N__21645));
    LocalMux I__4219 (
            .O(N__21654),
            .I(N__21642));
    LocalMux I__4218 (
            .O(N__21651),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    LocalMux I__4217 (
            .O(N__21648),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__4216 (
            .O(N__21645),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__4215 (
            .O(N__21642),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    InMux I__4214 (
            .O(N__21633),
            .I(N__21630));
    LocalMux I__4213 (
            .O(N__21630),
            .I(N__21627));
    Span4Mux_h I__4212 (
            .O(N__21627),
            .I(N__21624));
    Span4Mux_h I__4211 (
            .O(N__21624),
            .I(N__21621));
    Odrv4 I__4210 (
            .O(N__21621),
            .I(\this_sprites_ram.mem_out_bus6_1 ));
    InMux I__4209 (
            .O(N__21618),
            .I(N__21615));
    LocalMux I__4208 (
            .O(N__21615),
            .I(N__21612));
    Odrv12 I__4207 (
            .O(N__21612),
            .I(\this_sprites_ram.mem_out_bus2_1 ));
    InMux I__4206 (
            .O(N__21609),
            .I(N__21606));
    LocalMux I__4205 (
            .O(N__21606),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ));
    InMux I__4204 (
            .O(N__21603),
            .I(N__21600));
    LocalMux I__4203 (
            .O(N__21600),
            .I(N__21597));
    Span4Mux_h I__4202 (
            .O(N__21597),
            .I(N__21594));
    Span4Mux_h I__4201 (
            .O(N__21594),
            .I(N__21591));
    Span4Mux_v I__4200 (
            .O(N__21591),
            .I(N__21588));
    Odrv4 I__4199 (
            .O(N__21588),
            .I(\this_sprites_ram.mem_out_bus5_1 ));
    InMux I__4198 (
            .O(N__21585),
            .I(N__21582));
    LocalMux I__4197 (
            .O(N__21582),
            .I(N__21579));
    Span4Mux_h I__4196 (
            .O(N__21579),
            .I(N__21576));
    Span4Mux_h I__4195 (
            .O(N__21576),
            .I(N__21573));
    Span4Mux_v I__4194 (
            .O(N__21573),
            .I(N__21570));
    Odrv4 I__4193 (
            .O(N__21570),
            .I(\this_sprites_ram.mem_out_bus1_1 ));
    InMux I__4192 (
            .O(N__21567),
            .I(N__21564));
    LocalMux I__4191 (
            .O(N__21564),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ));
    InMux I__4190 (
            .O(N__21561),
            .I(N__21558));
    LocalMux I__4189 (
            .O(N__21558),
            .I(N__21555));
    Odrv12 I__4188 (
            .O(N__21555),
            .I(\this_sprites_ram.mem_out_bus7_1 ));
    InMux I__4187 (
            .O(N__21552),
            .I(N__21549));
    LocalMux I__4186 (
            .O(N__21549),
            .I(N__21546));
    Span4Mux_h I__4185 (
            .O(N__21546),
            .I(N__21543));
    Span4Mux_h I__4184 (
            .O(N__21543),
            .I(N__21540));
    Span4Mux_h I__4183 (
            .O(N__21540),
            .I(N__21537));
    Odrv4 I__4182 (
            .O(N__21537),
            .I(\this_sprites_ram.mem_out_bus3_1 ));
    InMux I__4181 (
            .O(N__21534),
            .I(N__21531));
    LocalMux I__4180 (
            .O(N__21531),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ));
    InMux I__4179 (
            .O(N__21528),
            .I(N__21525));
    LocalMux I__4178 (
            .O(N__21525),
            .I(N__21520));
    InMux I__4177 (
            .O(N__21524),
            .I(N__21516));
    InMux I__4176 (
            .O(N__21523),
            .I(N__21513));
    Span4Mux_h I__4175 (
            .O(N__21520),
            .I(N__21510));
    InMux I__4174 (
            .O(N__21519),
            .I(N__21507));
    LocalMux I__4173 (
            .O(N__21516),
            .I(N__21504));
    LocalMux I__4172 (
            .O(N__21513),
            .I(\this_ppu.M_count_d_0_sqmuxa ));
    Odrv4 I__4171 (
            .O(N__21510),
            .I(\this_ppu.M_count_d_0_sqmuxa ));
    LocalMux I__4170 (
            .O(N__21507),
            .I(\this_ppu.M_count_d_0_sqmuxa ));
    Odrv12 I__4169 (
            .O(N__21504),
            .I(\this_ppu.M_count_d_0_sqmuxa ));
    SRMux I__4168 (
            .O(N__21495),
            .I(N__21491));
    SRMux I__4167 (
            .O(N__21494),
            .I(N__21488));
    LocalMux I__4166 (
            .O(N__21491),
            .I(N__21485));
    LocalMux I__4165 (
            .O(N__21488),
            .I(N__21481));
    Span4Mux_v I__4164 (
            .O(N__21485),
            .I(N__21478));
    SRMux I__4163 (
            .O(N__21484),
            .I(N__21475));
    Span4Mux_h I__4162 (
            .O(N__21481),
            .I(N__21471));
    Span4Mux_h I__4161 (
            .O(N__21478),
            .I(N__21466));
    LocalMux I__4160 (
            .O(N__21475),
            .I(N__21466));
    SRMux I__4159 (
            .O(N__21474),
            .I(N__21463));
    Span4Mux_h I__4158 (
            .O(N__21471),
            .I(N__21460));
    Span4Mux_h I__4157 (
            .O(N__21466),
            .I(N__21457));
    LocalMux I__4156 (
            .O(N__21463),
            .I(N__21454));
    Odrv4 I__4155 (
            .O(N__21460),
            .I(\this_ppu.M_last_q_RNIQRTEB ));
    Odrv4 I__4154 (
            .O(N__21457),
            .I(\this_ppu.M_last_q_RNIQRTEB ));
    Odrv12 I__4153 (
            .O(N__21454),
            .I(\this_ppu.M_last_q_RNIQRTEB ));
    CascadeMux I__4152 (
            .O(N__21447),
            .I(N__21443));
    CascadeMux I__4151 (
            .O(N__21446),
            .I(N__21440));
    CascadeBuf I__4150 (
            .O(N__21443),
            .I(N__21437));
    InMux I__4149 (
            .O(N__21440),
            .I(N__21434));
    CascadeMux I__4148 (
            .O(N__21437),
            .I(N__21431));
    LocalMux I__4147 (
            .O(N__21434),
            .I(N__21428));
    InMux I__4146 (
            .O(N__21431),
            .I(N__21425));
    Span4Mux_v I__4145 (
            .O(N__21428),
            .I(N__21421));
    LocalMux I__4144 (
            .O(N__21425),
            .I(N__21418));
    InMux I__4143 (
            .O(N__21424),
            .I(N__21413));
    Sp12to4 I__4142 (
            .O(N__21421),
            .I(N__21410));
    Span12Mux_h I__4141 (
            .O(N__21418),
            .I(N__21407));
    InMux I__4140 (
            .O(N__21417),
            .I(N__21404));
    InMux I__4139 (
            .O(N__21416),
            .I(N__21401));
    LocalMux I__4138 (
            .O(N__21413),
            .I(N__21398));
    Span12Mux_h I__4137 (
            .O(N__21410),
            .I(N__21393));
    Span12Mux_v I__4136 (
            .O(N__21407),
            .I(N__21393));
    LocalMux I__4135 (
            .O(N__21404),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__4134 (
            .O(N__21401),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__4133 (
            .O(N__21398),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__4132 (
            .O(N__21393),
            .I(M_this_ppu_map_addr_1));
    InMux I__4131 (
            .O(N__21384),
            .I(N__21378));
    InMux I__4130 (
            .O(N__21383),
            .I(N__21378));
    LocalMux I__4129 (
            .O(N__21378),
            .I(\this_ppu.un1_M_haddress_q_3_c2 ));
    CascadeMux I__4128 (
            .O(N__21375),
            .I(N__21371));
    CascadeMux I__4127 (
            .O(N__21374),
            .I(N__21368));
    InMux I__4126 (
            .O(N__21371),
            .I(N__21365));
    CascadeBuf I__4125 (
            .O(N__21368),
            .I(N__21362));
    LocalMux I__4124 (
            .O(N__21365),
            .I(N__21358));
    CascadeMux I__4123 (
            .O(N__21362),
            .I(N__21355));
    InMux I__4122 (
            .O(N__21361),
            .I(N__21352));
    Span4Mux_h I__4121 (
            .O(N__21358),
            .I(N__21349));
    InMux I__4120 (
            .O(N__21355),
            .I(N__21346));
    LocalMux I__4119 (
            .O(N__21352),
            .I(N__21343));
    Span4Mux_h I__4118 (
            .O(N__21349),
            .I(N__21340));
    LocalMux I__4117 (
            .O(N__21346),
            .I(N__21337));
    Span4Mux_v I__4116 (
            .O(N__21343),
            .I(N__21331));
    Sp12to4 I__4115 (
            .O(N__21340),
            .I(N__21326));
    Span12Mux_h I__4114 (
            .O(N__21337),
            .I(N__21326));
    InMux I__4113 (
            .O(N__21336),
            .I(N__21321));
    InMux I__4112 (
            .O(N__21335),
            .I(N__21321));
    InMux I__4111 (
            .O(N__21334),
            .I(N__21318));
    Span4Mux_v I__4110 (
            .O(N__21331),
            .I(N__21315));
    Span12Mux_v I__4109 (
            .O(N__21326),
            .I(N__21312));
    LocalMux I__4108 (
            .O(N__21321),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__4107 (
            .O(N__21318),
            .I(M_this_ppu_map_addr_0));
    Odrv4 I__4106 (
            .O(N__21315),
            .I(M_this_ppu_map_addr_0));
    Odrv12 I__4105 (
            .O(N__21312),
            .I(M_this_ppu_map_addr_0));
    CascadeMux I__4104 (
            .O(N__21303),
            .I(N__21300));
    CascadeBuf I__4103 (
            .O(N__21300),
            .I(N__21297));
    CascadeMux I__4102 (
            .O(N__21297),
            .I(N__21294));
    InMux I__4101 (
            .O(N__21294),
            .I(N__21291));
    LocalMux I__4100 (
            .O(N__21291),
            .I(N__21287));
    InMux I__4099 (
            .O(N__21290),
            .I(N__21284));
    Span12Mux_h I__4098 (
            .O(N__21287),
            .I(N__21281));
    LocalMux I__4097 (
            .O(N__21284),
            .I(N__21277));
    Span12Mux_h I__4096 (
            .O(N__21281),
            .I(N__21274));
    InMux I__4095 (
            .O(N__21280),
            .I(N__21271));
    Span12Mux_h I__4094 (
            .O(N__21277),
            .I(N__21268));
    Span12Mux_v I__4093 (
            .O(N__21274),
            .I(N__21265));
    LocalMux I__4092 (
            .O(N__21271),
            .I(M_this_ppu_map_addr_4));
    Odrv12 I__4091 (
            .O(N__21268),
            .I(M_this_ppu_map_addr_4));
    Odrv12 I__4090 (
            .O(N__21265),
            .I(M_this_ppu_map_addr_4));
    InMux I__4089 (
            .O(N__21258),
            .I(N__21249));
    InMux I__4088 (
            .O(N__21257),
            .I(N__21249));
    InMux I__4087 (
            .O(N__21256),
            .I(N__21249));
    LocalMux I__4086 (
            .O(N__21249),
            .I(\this_ppu.un1_M_haddress_q_3_c5 ));
    CascadeMux I__4085 (
            .O(N__21246),
            .I(N__21242));
    CascadeMux I__4084 (
            .O(N__21245),
            .I(N__21239));
    CascadeBuf I__4083 (
            .O(N__21242),
            .I(N__21236));
    InMux I__4082 (
            .O(N__21239),
            .I(N__21232));
    CascadeMux I__4081 (
            .O(N__21236),
            .I(N__21229));
    InMux I__4080 (
            .O(N__21235),
            .I(N__21226));
    LocalMux I__4079 (
            .O(N__21232),
            .I(N__21223));
    InMux I__4078 (
            .O(N__21229),
            .I(N__21220));
    LocalMux I__4077 (
            .O(N__21226),
            .I(N__21215));
    Span4Mux_h I__4076 (
            .O(N__21223),
            .I(N__21212));
    LocalMux I__4075 (
            .O(N__21220),
            .I(N__21209));
    CascadeMux I__4074 (
            .O(N__21219),
            .I(N__21206));
    CascadeMux I__4073 (
            .O(N__21218),
            .I(N__21203));
    Span4Mux_v I__4072 (
            .O(N__21215),
            .I(N__21199));
    Sp12to4 I__4071 (
            .O(N__21212),
            .I(N__21194));
    Span12Mux_s11_h I__4070 (
            .O(N__21209),
            .I(N__21194));
    InMux I__4069 (
            .O(N__21206),
            .I(N__21187));
    InMux I__4068 (
            .O(N__21203),
            .I(N__21187));
    InMux I__4067 (
            .O(N__21202),
            .I(N__21187));
    Span4Mux_v I__4066 (
            .O(N__21199),
            .I(N__21184));
    Span12Mux_v I__4065 (
            .O(N__21194),
            .I(N__21181));
    LocalMux I__4064 (
            .O(N__21187),
            .I(M_this_ppu_map_addr_2));
    Odrv4 I__4063 (
            .O(N__21184),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__4062 (
            .O(N__21181),
            .I(M_this_ppu_map_addr_2));
    CascadeMux I__4061 (
            .O(N__21174),
            .I(N__21171));
    CascadeBuf I__4060 (
            .O(N__21171),
            .I(N__21167));
    CascadeMux I__4059 (
            .O(N__21170),
            .I(N__21164));
    CascadeMux I__4058 (
            .O(N__21167),
            .I(N__21161));
    InMux I__4057 (
            .O(N__21164),
            .I(N__21157));
    InMux I__4056 (
            .O(N__21161),
            .I(N__21154));
    InMux I__4055 (
            .O(N__21160),
            .I(N__21151));
    LocalMux I__4054 (
            .O(N__21157),
            .I(N__21148));
    LocalMux I__4053 (
            .O(N__21154),
            .I(N__21145));
    LocalMux I__4052 (
            .O(N__21151),
            .I(N__21142));
    Span4Mux_v I__4051 (
            .O(N__21148),
            .I(N__21139));
    Sp12to4 I__4050 (
            .O(N__21145),
            .I(N__21136));
    Span4Mux_v I__4049 (
            .O(N__21142),
            .I(N__21131));
    Span4Mux_h I__4048 (
            .O(N__21139),
            .I(N__21128));
    Span12Mux_h I__4047 (
            .O(N__21136),
            .I(N__21125));
    InMux I__4046 (
            .O(N__21135),
            .I(N__21120));
    InMux I__4045 (
            .O(N__21134),
            .I(N__21120));
    Span4Mux_v I__4044 (
            .O(N__21131),
            .I(N__21117));
    Span4Mux_h I__4043 (
            .O(N__21128),
            .I(N__21114));
    Span12Mux_v I__4042 (
            .O(N__21125),
            .I(N__21111));
    LocalMux I__4041 (
            .O(N__21120),
            .I(M_this_ppu_map_addr_3));
    Odrv4 I__4040 (
            .O(N__21117),
            .I(M_this_ppu_map_addr_3));
    Odrv4 I__4039 (
            .O(N__21114),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__4038 (
            .O(N__21111),
            .I(M_this_ppu_map_addr_3));
    CEMux I__4037 (
            .O(N__21102),
            .I(N__21099));
    LocalMux I__4036 (
            .O(N__21099),
            .I(N__21096));
    Span4Mux_v I__4035 (
            .O(N__21096),
            .I(N__21093));
    Span4Mux_h I__4034 (
            .O(N__21093),
            .I(N__21089));
    InMux I__4033 (
            .O(N__21092),
            .I(N__21086));
    Span4Mux_h I__4032 (
            .O(N__21089),
            .I(N__21082));
    LocalMux I__4031 (
            .O(N__21086),
            .I(N__21079));
    InMux I__4030 (
            .O(N__21085),
            .I(N__21076));
    Odrv4 I__4029 (
            .O(N__21082),
            .I(M_this_ppu_vram_en_0));
    Odrv4 I__4028 (
            .O(N__21079),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__4027 (
            .O(N__21076),
            .I(M_this_ppu_vram_en_0));
    SRMux I__4026 (
            .O(N__21069),
            .I(N__21064));
    SRMux I__4025 (
            .O(N__21068),
            .I(N__21061));
    SRMux I__4024 (
            .O(N__21067),
            .I(N__21058));
    LocalMux I__4023 (
            .O(N__21064),
            .I(N__21055));
    LocalMux I__4022 (
            .O(N__21061),
            .I(N__21052));
    LocalMux I__4021 (
            .O(N__21058),
            .I(N__21049));
    Span4Mux_v I__4020 (
            .O(N__21055),
            .I(N__21046));
    Span4Mux_v I__4019 (
            .O(N__21052),
            .I(N__21041));
    Span4Mux_h I__4018 (
            .O(N__21049),
            .I(N__21041));
    Odrv4 I__4017 (
            .O(N__21046),
            .I(\this_ppu.M_last_q_RNI3BB75 ));
    Odrv4 I__4016 (
            .O(N__21041),
            .I(\this_ppu.M_last_q_RNI3BB75 ));
    InMux I__4015 (
            .O(N__21036),
            .I(N__21033));
    LocalMux I__4014 (
            .O(N__21033),
            .I(N__21030));
    Span4Mux_v I__4013 (
            .O(N__21030),
            .I(N__21027));
    Span4Mux_h I__4012 (
            .O(N__21027),
            .I(N__21024));
    Sp12to4 I__4011 (
            .O(N__21024),
            .I(N__21021));
    Span12Mux_v I__4010 (
            .O(N__21021),
            .I(N__21018));
    Odrv12 I__4009 (
            .O(N__21018),
            .I(M_this_oam_ram_read_data_1));
    InMux I__4008 (
            .O(N__21015),
            .I(N__21012));
    LocalMux I__4007 (
            .O(N__21012),
            .I(N__21009));
    Span4Mux_v I__4006 (
            .O(N__21009),
            .I(N__21006));
    Sp12to4 I__4005 (
            .O(N__21006),
            .I(N__21003));
    Span12Mux_h I__4004 (
            .O(N__21003),
            .I(N__21000));
    Odrv12 I__4003 (
            .O(N__21000),
            .I(M_this_map_ram_read_data_1));
    CascadeMux I__4002 (
            .O(N__20997),
            .I(N__20989));
    CascadeMux I__4001 (
            .O(N__20996),
            .I(N__20984));
    CascadeMux I__4000 (
            .O(N__20995),
            .I(N__20981));
    CascadeMux I__3999 (
            .O(N__20994),
            .I(N__20977));
    CascadeMux I__3998 (
            .O(N__20993),
            .I(N__20973));
    CascadeMux I__3997 (
            .O(N__20992),
            .I(N__20969));
    InMux I__3996 (
            .O(N__20989),
            .I(N__20966));
    CascadeMux I__3995 (
            .O(N__20988),
            .I(N__20963));
    CascadeMux I__3994 (
            .O(N__20987),
            .I(N__20958));
    InMux I__3993 (
            .O(N__20984),
            .I(N__20953));
    InMux I__3992 (
            .O(N__20981),
            .I(N__20950));
    CascadeMux I__3991 (
            .O(N__20980),
            .I(N__20947));
    InMux I__3990 (
            .O(N__20977),
            .I(N__20944));
    CascadeMux I__3989 (
            .O(N__20976),
            .I(N__20941));
    InMux I__3988 (
            .O(N__20973),
            .I(N__20938));
    CascadeMux I__3987 (
            .O(N__20972),
            .I(N__20935));
    InMux I__3986 (
            .O(N__20969),
            .I(N__20932));
    LocalMux I__3985 (
            .O(N__20966),
            .I(N__20929));
    InMux I__3984 (
            .O(N__20963),
            .I(N__20926));
    CascadeMux I__3983 (
            .O(N__20962),
            .I(N__20923));
    CascadeMux I__3982 (
            .O(N__20961),
            .I(N__20920));
    InMux I__3981 (
            .O(N__20958),
            .I(N__20917));
    CascadeMux I__3980 (
            .O(N__20957),
            .I(N__20913));
    CascadeMux I__3979 (
            .O(N__20956),
            .I(N__20910));
    LocalMux I__3978 (
            .O(N__20953),
            .I(N__20907));
    LocalMux I__3977 (
            .O(N__20950),
            .I(N__20904));
    InMux I__3976 (
            .O(N__20947),
            .I(N__20901));
    LocalMux I__3975 (
            .O(N__20944),
            .I(N__20898));
    InMux I__3974 (
            .O(N__20941),
            .I(N__20895));
    LocalMux I__3973 (
            .O(N__20938),
            .I(N__20892));
    InMux I__3972 (
            .O(N__20935),
            .I(N__20889));
    LocalMux I__3971 (
            .O(N__20932),
            .I(N__20886));
    Span4Mux_h I__3970 (
            .O(N__20929),
            .I(N__20883));
    LocalMux I__3969 (
            .O(N__20926),
            .I(N__20880));
    InMux I__3968 (
            .O(N__20923),
            .I(N__20877));
    InMux I__3967 (
            .O(N__20920),
            .I(N__20874));
    LocalMux I__3966 (
            .O(N__20917),
            .I(N__20871));
    CascadeMux I__3965 (
            .O(N__20916),
            .I(N__20868));
    InMux I__3964 (
            .O(N__20913),
            .I(N__20865));
    InMux I__3963 (
            .O(N__20910),
            .I(N__20862));
    Span4Mux_h I__3962 (
            .O(N__20907),
            .I(N__20859));
    Span4Mux_h I__3961 (
            .O(N__20904),
            .I(N__20856));
    LocalMux I__3960 (
            .O(N__20901),
            .I(N__20853));
    Span4Mux_h I__3959 (
            .O(N__20898),
            .I(N__20850));
    LocalMux I__3958 (
            .O(N__20895),
            .I(N__20847));
    Span4Mux_h I__3957 (
            .O(N__20892),
            .I(N__20844));
    LocalMux I__3956 (
            .O(N__20889),
            .I(N__20841));
    Span4Mux_h I__3955 (
            .O(N__20886),
            .I(N__20836));
    Span4Mux_v I__3954 (
            .O(N__20883),
            .I(N__20836));
    Span4Mux_h I__3953 (
            .O(N__20880),
            .I(N__20833));
    LocalMux I__3952 (
            .O(N__20877),
            .I(N__20830));
    LocalMux I__3951 (
            .O(N__20874),
            .I(N__20827));
    Span4Mux_h I__3950 (
            .O(N__20871),
            .I(N__20824));
    InMux I__3949 (
            .O(N__20868),
            .I(N__20821));
    LocalMux I__3948 (
            .O(N__20865),
            .I(N__20818));
    LocalMux I__3947 (
            .O(N__20862),
            .I(N__20815));
    Span4Mux_h I__3946 (
            .O(N__20859),
            .I(N__20810));
    Span4Mux_h I__3945 (
            .O(N__20856),
            .I(N__20810));
    Span4Mux_h I__3944 (
            .O(N__20853),
            .I(N__20807));
    Span4Mux_h I__3943 (
            .O(N__20850),
            .I(N__20804));
    Span4Mux_h I__3942 (
            .O(N__20847),
            .I(N__20801));
    Span4Mux_h I__3941 (
            .O(N__20844),
            .I(N__20798));
    Span4Mux_h I__3940 (
            .O(N__20841),
            .I(N__20793));
    Span4Mux_v I__3939 (
            .O(N__20836),
            .I(N__20793));
    Span4Mux_h I__3938 (
            .O(N__20833),
            .I(N__20790));
    Span4Mux_h I__3937 (
            .O(N__20830),
            .I(N__20787));
    Span4Mux_h I__3936 (
            .O(N__20827),
            .I(N__20782));
    Span4Mux_v I__3935 (
            .O(N__20824),
            .I(N__20782));
    LocalMux I__3934 (
            .O(N__20821),
            .I(N__20775));
    Span4Mux_v I__3933 (
            .O(N__20818),
            .I(N__20775));
    Span4Mux_v I__3932 (
            .O(N__20815),
            .I(N__20775));
    Span4Mux_h I__3931 (
            .O(N__20810),
            .I(N__20768));
    Span4Mux_h I__3930 (
            .O(N__20807),
            .I(N__20768));
    Span4Mux_h I__3929 (
            .O(N__20804),
            .I(N__20768));
    Span4Mux_h I__3928 (
            .O(N__20801),
            .I(N__20759));
    Span4Mux_h I__3927 (
            .O(N__20798),
            .I(N__20759));
    Span4Mux_h I__3926 (
            .O(N__20793),
            .I(N__20759));
    Span4Mux_h I__3925 (
            .O(N__20790),
            .I(N__20759));
    Span4Mux_h I__3924 (
            .O(N__20787),
            .I(N__20754));
    Span4Mux_h I__3923 (
            .O(N__20782),
            .I(N__20754));
    Sp12to4 I__3922 (
            .O(N__20775),
            .I(N__20751));
    Sp12to4 I__3921 (
            .O(N__20768),
            .I(N__20742));
    Sp12to4 I__3920 (
            .O(N__20759),
            .I(N__20742));
    Sp12to4 I__3919 (
            .O(N__20754),
            .I(N__20742));
    Span12Mux_h I__3918 (
            .O(N__20751),
            .I(N__20742));
    Odrv12 I__3917 (
            .O(N__20742),
            .I(M_this_ppu_sprites_addr_7));
    CascadeMux I__3916 (
            .O(N__20739),
            .I(N__20736));
    InMux I__3915 (
            .O(N__20736),
            .I(N__20732));
    CascadeMux I__3914 (
            .O(N__20735),
            .I(N__20729));
    LocalMux I__3913 (
            .O(N__20732),
            .I(N__20726));
    InMux I__3912 (
            .O(N__20729),
            .I(N__20723));
    Odrv4 I__3911 (
            .O(N__20726),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    LocalMux I__3910 (
            .O(N__20723),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    CascadeMux I__3909 (
            .O(N__20718),
            .I(N__20715));
    InMux I__3908 (
            .O(N__20715),
            .I(N__20711));
    CascadeMux I__3907 (
            .O(N__20714),
            .I(N__20708));
    LocalMux I__3906 (
            .O(N__20711),
            .I(N__20705));
    InMux I__3905 (
            .O(N__20708),
            .I(N__20702));
    Odrv4 I__3904 (
            .O(N__20705),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    LocalMux I__3903 (
            .O(N__20702),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    InMux I__3902 (
            .O(N__20697),
            .I(bfn_19_8_0_));
    InMux I__3901 (
            .O(N__20694),
            .I(N__20691));
    LocalMux I__3900 (
            .O(N__20691),
            .I(N__20688));
    Span4Mux_h I__3899 (
            .O(N__20688),
            .I(N__20683));
    InMux I__3898 (
            .O(N__20687),
            .I(N__20680));
    InMux I__3897 (
            .O(N__20686),
            .I(N__20677));
    Odrv4 I__3896 (
            .O(N__20683),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    LocalMux I__3895 (
            .O(N__20680),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    LocalMux I__3894 (
            .O(N__20677),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    InMux I__3893 (
            .O(N__20670),
            .I(N__20666));
    InMux I__3892 (
            .O(N__20669),
            .I(N__20662));
    LocalMux I__3891 (
            .O(N__20666),
            .I(N__20659));
    InMux I__3890 (
            .O(N__20665),
            .I(N__20656));
    LocalMux I__3889 (
            .O(N__20662),
            .I(N__20651));
    Span4Mux_v I__3888 (
            .O(N__20659),
            .I(N__20651));
    LocalMux I__3887 (
            .O(N__20656),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__3886 (
            .O(N__20651),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    InMux I__3885 (
            .O(N__20646),
            .I(N__20643));
    LocalMux I__3884 (
            .O(N__20643),
            .I(N__20639));
    CascadeMux I__3883 (
            .O(N__20642),
            .I(N__20636));
    Span4Mux_h I__3882 (
            .O(N__20639),
            .I(N__20633));
    InMux I__3881 (
            .O(N__20636),
            .I(N__20630));
    Odrv4 I__3880 (
            .O(N__20633),
            .I(\this_ppu.N_122 ));
    LocalMux I__3879 (
            .O(N__20630),
            .I(\this_ppu.N_122 ));
    InMux I__3878 (
            .O(N__20625),
            .I(N__20622));
    LocalMux I__3877 (
            .O(N__20622),
            .I(N__20617));
    InMux I__3876 (
            .O(N__20621),
            .I(N__20612));
    InMux I__3875 (
            .O(N__20620),
            .I(N__20612));
    Span4Mux_v I__3874 (
            .O(N__20617),
            .I(N__20607));
    LocalMux I__3873 (
            .O(N__20612),
            .I(N__20607));
    Odrv4 I__3872 (
            .O(N__20607),
            .I(\this_ppu.un1_M_vaddress_q_2_c2 ));
    InMux I__3871 (
            .O(N__20604),
            .I(N__20600));
    InMux I__3870 (
            .O(N__20603),
            .I(N__20597));
    LocalMux I__3869 (
            .O(N__20600),
            .I(N__20594));
    LocalMux I__3868 (
            .O(N__20597),
            .I(N__20590));
    Span4Mux_h I__3867 (
            .O(N__20594),
            .I(N__20586));
    InMux I__3866 (
            .O(N__20593),
            .I(N__20582));
    Span4Mux_v I__3865 (
            .O(N__20590),
            .I(N__20579));
    CascadeMux I__3864 (
            .O(N__20589),
            .I(N__20576));
    Sp12to4 I__3863 (
            .O(N__20586),
            .I(N__20573));
    InMux I__3862 (
            .O(N__20585),
            .I(N__20570));
    LocalMux I__3861 (
            .O(N__20582),
            .I(N__20567));
    Sp12to4 I__3860 (
            .O(N__20579),
            .I(N__20564));
    InMux I__3859 (
            .O(N__20576),
            .I(N__20561));
    Span12Mux_v I__3858 (
            .O(N__20573),
            .I(N__20558));
    LocalMux I__3857 (
            .O(N__20570),
            .I(N__20555));
    Span4Mux_v I__3856 (
            .O(N__20567),
            .I(N__20552));
    Span12Mux_s11_h I__3855 (
            .O(N__20564),
            .I(N__20547));
    LocalMux I__3854 (
            .O(N__20561),
            .I(N__20547));
    Odrv12 I__3853 (
            .O(N__20558),
            .I(this_vga_signals_vvisibility));
    Odrv12 I__3852 (
            .O(N__20555),
            .I(this_vga_signals_vvisibility));
    Odrv4 I__3851 (
            .O(N__20552),
            .I(this_vga_signals_vvisibility));
    Odrv12 I__3850 (
            .O(N__20547),
            .I(this_vga_signals_vvisibility));
    InMux I__3849 (
            .O(N__20538),
            .I(bfn_19_6_0_));
    CascadeMux I__3848 (
            .O(N__20535),
            .I(N__20532));
    InMux I__3847 (
            .O(N__20532),
            .I(N__20528));
    CascadeMux I__3846 (
            .O(N__20531),
            .I(N__20525));
    LocalMux I__3845 (
            .O(N__20528),
            .I(N__20522));
    InMux I__3844 (
            .O(N__20525),
            .I(N__20519));
    Odrv4 I__3843 (
            .O(N__20522),
            .I(\this_ppu.M_this_ppu_vram_addr_i_0 ));
    LocalMux I__3842 (
            .O(N__20519),
            .I(\this_ppu.M_this_ppu_vram_addr_i_0 ));
    InMux I__3841 (
            .O(N__20514),
            .I(N__20510));
    CascadeMux I__3840 (
            .O(N__20513),
            .I(N__20507));
    LocalMux I__3839 (
            .O(N__20510),
            .I(N__20504));
    InMux I__3838 (
            .O(N__20507),
            .I(N__20501));
    Odrv4 I__3837 (
            .O(N__20504),
            .I(\this_ppu.M_this_ppu_vram_addr_i_1 ));
    LocalMux I__3836 (
            .O(N__20501),
            .I(\this_ppu.M_this_ppu_vram_addr_i_1 ));
    InMux I__3835 (
            .O(N__20496),
            .I(N__20493));
    LocalMux I__3834 (
            .O(N__20493),
            .I(N__20489));
    InMux I__3833 (
            .O(N__20492),
            .I(N__20486));
    Odrv4 I__3832 (
            .O(N__20489),
            .I(\this_ppu.M_this_ppu_vram_addr_i_2 ));
    LocalMux I__3831 (
            .O(N__20486),
            .I(\this_ppu.M_this_ppu_vram_addr_i_2 ));
    CascadeMux I__3830 (
            .O(N__20481),
            .I(N__20478));
    InMux I__3829 (
            .O(N__20478),
            .I(N__20474));
    CascadeMux I__3828 (
            .O(N__20477),
            .I(N__20471));
    LocalMux I__3827 (
            .O(N__20474),
            .I(N__20468));
    InMux I__3826 (
            .O(N__20471),
            .I(N__20465));
    Odrv4 I__3825 (
            .O(N__20468),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    LocalMux I__3824 (
            .O(N__20465),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    CascadeMux I__3823 (
            .O(N__20460),
            .I(N__20457));
    InMux I__3822 (
            .O(N__20457),
            .I(N__20454));
    LocalMux I__3821 (
            .O(N__20454),
            .I(N__20450));
    InMux I__3820 (
            .O(N__20453),
            .I(N__20447));
    Odrv4 I__3819 (
            .O(N__20450),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    LocalMux I__3818 (
            .O(N__20447),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    CascadeMux I__3817 (
            .O(N__20442),
            .I(N__20439));
    InMux I__3816 (
            .O(N__20439),
            .I(N__20435));
    CascadeMux I__3815 (
            .O(N__20438),
            .I(N__20432));
    LocalMux I__3814 (
            .O(N__20435),
            .I(N__20429));
    InMux I__3813 (
            .O(N__20432),
            .I(N__20426));
    Odrv4 I__3812 (
            .O(N__20429),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    LocalMux I__3811 (
            .O(N__20426),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    InMux I__3810 (
            .O(N__20421),
            .I(N__20418));
    LocalMux I__3809 (
            .O(N__20418),
            .I(N_617));
    InMux I__3808 (
            .O(N__20415),
            .I(N__20412));
    LocalMux I__3807 (
            .O(N__20412),
            .I(M_this_sprites_address_qc_11_0));
    InMux I__3806 (
            .O(N__20409),
            .I(N__20406));
    LocalMux I__3805 (
            .O(N__20406),
            .I(N_896_0));
    InMux I__3804 (
            .O(N__20403),
            .I(N__20400));
    LocalMux I__3803 (
            .O(N__20400),
            .I(N_512_0));
    CascadeMux I__3802 (
            .O(N__20397),
            .I(N__20394));
    InMux I__3801 (
            .O(N__20394),
            .I(N__20391));
    LocalMux I__3800 (
            .O(N__20391),
            .I(N__20388));
    Odrv4 I__3799 (
            .O(N__20388),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_8 ));
    InMux I__3798 (
            .O(N__20385),
            .I(N__20382));
    LocalMux I__3797 (
            .O(N__20382),
            .I(N__20379));
    Span4Mux_v I__3796 (
            .O(N__20379),
            .I(N__20376));
    Odrv4 I__3795 (
            .O(N__20376),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1Z0Z_5 ));
    CascadeMux I__3794 (
            .O(N__20373),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_11_cascade_ ));
    InMux I__3793 (
            .O(N__20370),
            .I(N__20367));
    LocalMux I__3792 (
            .O(N__20367),
            .I(N__20364));
    Odrv4 I__3791 (
            .O(N__20364),
            .I(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_1));
    InMux I__3790 (
            .O(N__20361),
            .I(N__20358));
    LocalMux I__3789 (
            .O(N__20358),
            .I(M_this_sprites_address_qc_10_0));
    CascadeMux I__3788 (
            .O(N__20355),
            .I(N_1286_tz_0_cascade_));
    CascadeMux I__3787 (
            .O(N__20352),
            .I(N_562_cascade_));
    InMux I__3786 (
            .O(N__20349),
            .I(N__20346));
    LocalMux I__3785 (
            .O(N__20346),
            .I(M_this_sprites_address_q_0_0_i_476));
    CascadeMux I__3784 (
            .O(N__20343),
            .I(M_this_sprites_address_q_0_0_i_496_cascade_));
    InMux I__3783 (
            .O(N__20340),
            .I(N__20337));
    LocalMux I__3782 (
            .O(N__20337),
            .I(M_this_sprites_address_qc_0_1));
    CascadeMux I__3781 (
            .O(N__20334),
            .I(N__20331));
    InMux I__3780 (
            .O(N__20331),
            .I(N__20328));
    LocalMux I__3779 (
            .O(N__20328),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_0 ));
    CascadeMux I__3778 (
            .O(N__20325),
            .I(N_773_cascade_));
    InMux I__3777 (
            .O(N__20322),
            .I(N__20319));
    LocalMux I__3776 (
            .O(N__20319),
            .I(M_this_sprites_address_q_0_0_i_492));
    CascadeMux I__3775 (
            .O(N__20316),
            .I(M_this_sprites_address_qc_1_0_cascade_));
    CascadeMux I__3774 (
            .O(N__20313),
            .I(\this_vga_signals.N_419_0_cascade_ ));
    CascadeMux I__3773 (
            .O(N__20310),
            .I(N_440_0_cascade_));
    CascadeMux I__3772 (
            .O(N__20307),
            .I(\this_vga_signals.N_467_0_cascade_ ));
    InMux I__3771 (
            .O(N__20304),
            .I(N__20301));
    LocalMux I__3770 (
            .O(N__20301),
            .I(\this_vga_signals.N_467_0 ));
    CascadeMux I__3769 (
            .O(N__20298),
            .I(N__20295));
    InMux I__3768 (
            .O(N__20295),
            .I(N__20292));
    LocalMux I__3767 (
            .O(N__20292),
            .I(N__20289));
    Span4Mux_v I__3766 (
            .O(N__20289),
            .I(N__20286));
    Odrv4 I__3765 (
            .O(N__20286),
            .I(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_6 ));
    InMux I__3764 (
            .O(N__20283),
            .I(N__20280));
    LocalMux I__3763 (
            .O(N__20280),
            .I(N_510_0));
    InMux I__3762 (
            .O(N__20277),
            .I(N__20274));
    LocalMux I__3761 (
            .O(N__20274),
            .I(N__20271));
    Odrv4 I__3760 (
            .O(N__20271),
            .I(M_this_sprites_address_qc_5_0));
    InMux I__3759 (
            .O(N__20268),
            .I(N__20265));
    LocalMux I__3758 (
            .O(N__20265),
            .I(N__20262));
    Span4Mux_v I__3757 (
            .O(N__20262),
            .I(N__20259));
    Span4Mux_h I__3756 (
            .O(N__20259),
            .I(N__20256));
    Span4Mux_h I__3755 (
            .O(N__20256),
            .I(N__20253));
    Odrv4 I__3754 (
            .O(N__20253),
            .I(\this_sprites_ram.mem_out_bus5_2 ));
    InMux I__3753 (
            .O(N__20250),
            .I(N__20247));
    LocalMux I__3752 (
            .O(N__20247),
            .I(N__20244));
    Span4Mux_h I__3751 (
            .O(N__20244),
            .I(N__20241));
    Span4Mux_h I__3750 (
            .O(N__20241),
            .I(N__20238));
    Odrv4 I__3749 (
            .O(N__20238),
            .I(\this_sprites_ram.mem_out_bus1_2 ));
    InMux I__3748 (
            .O(N__20235),
            .I(N__20232));
    LocalMux I__3747 (
            .O(N__20232),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ));
    IoInMux I__3746 (
            .O(N__20229),
            .I(N__20225));
    IoInMux I__3745 (
            .O(N__20228),
            .I(N__20222));
    LocalMux I__3744 (
            .O(N__20225),
            .I(N__20216));
    LocalMux I__3743 (
            .O(N__20222),
            .I(N__20216));
    IoInMux I__3742 (
            .O(N__20221),
            .I(N__20208));
    IoSpan4Mux I__3741 (
            .O(N__20216),
            .I(N__20205));
    IoInMux I__3740 (
            .O(N__20215),
            .I(N__20202));
    IoInMux I__3739 (
            .O(N__20214),
            .I(N__20199));
    IoInMux I__3738 (
            .O(N__20213),
            .I(N__20196));
    IoInMux I__3737 (
            .O(N__20212),
            .I(N__20193));
    IoInMux I__3736 (
            .O(N__20211),
            .I(N__20189));
    LocalMux I__3735 (
            .O(N__20208),
            .I(N__20184));
    IoSpan4Mux I__3734 (
            .O(N__20205),
            .I(N__20181));
    LocalMux I__3733 (
            .O(N__20202),
            .I(N__20172));
    LocalMux I__3732 (
            .O(N__20199),
            .I(N__20172));
    LocalMux I__3731 (
            .O(N__20196),
            .I(N__20172));
    LocalMux I__3730 (
            .O(N__20193),
            .I(N__20172));
    IoInMux I__3729 (
            .O(N__20192),
            .I(N__20169));
    LocalMux I__3728 (
            .O(N__20189),
            .I(N__20166));
    IoInMux I__3727 (
            .O(N__20188),
            .I(N__20163));
    IoInMux I__3726 (
            .O(N__20187),
            .I(N__20160));
    Span4Mux_s1_h I__3725 (
            .O(N__20184),
            .I(N__20152));
    IoSpan4Mux I__3724 (
            .O(N__20181),
            .I(N__20144));
    IoSpan4Mux I__3723 (
            .O(N__20172),
            .I(N__20144));
    LocalMux I__3722 (
            .O(N__20169),
            .I(N__20144));
    IoSpan4Mux I__3721 (
            .O(N__20166),
            .I(N__20139));
    LocalMux I__3720 (
            .O(N__20163),
            .I(N__20139));
    LocalMux I__3719 (
            .O(N__20160),
            .I(N__20136));
    IoInMux I__3718 (
            .O(N__20159),
            .I(N__20133));
    IoInMux I__3717 (
            .O(N__20158),
            .I(N__20130));
    IoInMux I__3716 (
            .O(N__20157),
            .I(N__20127));
    IoInMux I__3715 (
            .O(N__20156),
            .I(N__20124));
    IoInMux I__3714 (
            .O(N__20155),
            .I(N__20121));
    Span4Mux_h I__3713 (
            .O(N__20152),
            .I(N__20118));
    IoInMux I__3712 (
            .O(N__20151),
            .I(N__20115));
    IoSpan4Mux I__3711 (
            .O(N__20144),
            .I(N__20112));
    IoSpan4Mux I__3710 (
            .O(N__20139),
            .I(N__20105));
    IoSpan4Mux I__3709 (
            .O(N__20136),
            .I(N__20105));
    LocalMux I__3708 (
            .O(N__20133),
            .I(N__20105));
    LocalMux I__3707 (
            .O(N__20130),
            .I(N__20100));
    LocalMux I__3706 (
            .O(N__20127),
            .I(N__20100));
    LocalMux I__3705 (
            .O(N__20124),
            .I(N__20097));
    LocalMux I__3704 (
            .O(N__20121),
            .I(N__20094));
    Sp12to4 I__3703 (
            .O(N__20118),
            .I(N__20091));
    LocalMux I__3702 (
            .O(N__20115),
            .I(N__20088));
    Span4Mux_s0_h I__3701 (
            .O(N__20112),
            .I(N__20085));
    IoSpan4Mux I__3700 (
            .O(N__20105),
            .I(N__20080));
    IoSpan4Mux I__3699 (
            .O(N__20100),
            .I(N__20080));
    Span12Mux_s4_v I__3698 (
            .O(N__20097),
            .I(N__20075));
    Span12Mux_s2_h I__3697 (
            .O(N__20094),
            .I(N__20075));
    Span12Mux_v I__3696 (
            .O(N__20091),
            .I(N__20072));
    Span12Mux_s2_h I__3695 (
            .O(N__20088),
            .I(N__20067));
    Sp12to4 I__3694 (
            .O(N__20085),
            .I(N__20067));
    Span4Mux_s3_v I__3693 (
            .O(N__20080),
            .I(N__20064));
    Span12Mux_h I__3692 (
            .O(N__20075),
            .I(N__20055));
    Span12Mux_h I__3691 (
            .O(N__20072),
            .I(N__20055));
    Span12Mux_h I__3690 (
            .O(N__20067),
            .I(N__20055));
    Sp12to4 I__3689 (
            .O(N__20064),
            .I(N__20055));
    Odrv12 I__3688 (
            .O(N__20055),
            .I(dma_0_i));
    InMux I__3687 (
            .O(N__20052),
            .I(N__20049));
    LocalMux I__3686 (
            .O(N__20049),
            .I(N__20046));
    Span12Mux_h I__3685 (
            .O(N__20046),
            .I(N__20043));
    Span12Mux_v I__3684 (
            .O(N__20043),
            .I(N__20040));
    Odrv12 I__3683 (
            .O(N__20040),
            .I(\this_sprites_ram.mem_out_bus4_3 ));
    InMux I__3682 (
            .O(N__20037),
            .I(N__20034));
    LocalMux I__3681 (
            .O(N__20034),
            .I(N__20031));
    Span4Mux_v I__3680 (
            .O(N__20031),
            .I(N__20028));
    Span4Mux_h I__3679 (
            .O(N__20028),
            .I(N__20025));
    Span4Mux_v I__3678 (
            .O(N__20025),
            .I(N__20022));
    Odrv4 I__3677 (
            .O(N__20022),
            .I(\this_sprites_ram.mem_out_bus0_3 ));
    CascadeMux I__3676 (
            .O(N__20019),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0_cascade_ ));
    CascadeMux I__3675 (
            .O(N__20016),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ));
    InMux I__3674 (
            .O(N__20013),
            .I(N__20010));
    LocalMux I__3673 (
            .O(N__20010),
            .I(N__20007));
    Span4Mux_h I__3672 (
            .O(N__20007),
            .I(N__20003));
    CascadeMux I__3671 (
            .O(N__20006),
            .I(N__20000));
    Span4Mux_h I__3670 (
            .O(N__20003),
            .I(N__19997));
    InMux I__3669 (
            .O(N__20000),
            .I(N__19994));
    Span4Mux_h I__3668 (
            .O(N__19997),
            .I(N__19991));
    LocalMux I__3667 (
            .O(N__19994),
            .I(N__19988));
    Odrv4 I__3666 (
            .O(N__19991),
            .I(M_this_ppu_vram_data_3));
    Odrv4 I__3665 (
            .O(N__19988),
            .I(M_this_ppu_vram_data_3));
    InMux I__3664 (
            .O(N__19983),
            .I(N__19980));
    LocalMux I__3663 (
            .O(N__19980),
            .I(N__19977));
    Span4Mux_h I__3662 (
            .O(N__19977),
            .I(N__19974));
    Span4Mux_v I__3661 (
            .O(N__19974),
            .I(N__19971));
    Span4Mux_h I__3660 (
            .O(N__19971),
            .I(N__19968));
    Odrv4 I__3659 (
            .O(N__19968),
            .I(\this_sprites_ram.mem_out_bus5_3 ));
    InMux I__3658 (
            .O(N__19965),
            .I(N__19962));
    LocalMux I__3657 (
            .O(N__19962),
            .I(N__19959));
    Span4Mux_v I__3656 (
            .O(N__19959),
            .I(N__19956));
    Span4Mux_h I__3655 (
            .O(N__19956),
            .I(N__19953));
    Odrv4 I__3654 (
            .O(N__19953),
            .I(\this_sprites_ram.mem_out_bus1_3 ));
    InMux I__3653 (
            .O(N__19950),
            .I(N__19947));
    LocalMux I__3652 (
            .O(N__19947),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ));
    InMux I__3651 (
            .O(N__19944),
            .I(N__19941));
    LocalMux I__3650 (
            .O(N__19941),
            .I(N__19938));
    Span4Mux_h I__3649 (
            .O(N__19938),
            .I(N__19935));
    Span4Mux_h I__3648 (
            .O(N__19935),
            .I(N__19932));
    Odrv4 I__3647 (
            .O(N__19932),
            .I(\this_sprites_ram.mem_out_bus7_3 ));
    InMux I__3646 (
            .O(N__19929),
            .I(N__19926));
    LocalMux I__3645 (
            .O(N__19926),
            .I(N__19923));
    Span4Mux_v I__3644 (
            .O(N__19923),
            .I(N__19920));
    Span4Mux_v I__3643 (
            .O(N__19920),
            .I(N__19917));
    Sp12to4 I__3642 (
            .O(N__19917),
            .I(N__19914));
    Odrv12 I__3641 (
            .O(N__19914),
            .I(\this_sprites_ram.mem_out_bus3_3 ));
    InMux I__3640 (
            .O(N__19911),
            .I(N__19908));
    LocalMux I__3639 (
            .O(N__19908),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ));
    InMux I__3638 (
            .O(N__19905),
            .I(N__19901));
    InMux I__3637 (
            .O(N__19904),
            .I(N__19898));
    LocalMux I__3636 (
            .O(N__19901),
            .I(N__19891));
    LocalMux I__3635 (
            .O(N__19898),
            .I(N__19891));
    InMux I__3634 (
            .O(N__19897),
            .I(N__19886));
    InMux I__3633 (
            .O(N__19896),
            .I(N__19886));
    Odrv4 I__3632 (
            .O(N__19891),
            .I(M_this_vga_signals_line_clk_0));
    LocalMux I__3631 (
            .O(N__19886),
            .I(M_this_vga_signals_line_clk_0));
    InMux I__3630 (
            .O(N__19881),
            .I(N__19878));
    LocalMux I__3629 (
            .O(N__19878),
            .I(N__19875));
    Span4Mux_v I__3628 (
            .O(N__19875),
            .I(N__19872));
    Sp12to4 I__3627 (
            .O(N__19872),
            .I(N__19869));
    Span12Mux_h I__3626 (
            .O(N__19869),
            .I(N__19866));
    Span12Mux_v I__3625 (
            .O(N__19866),
            .I(N__19863));
    Odrv12 I__3624 (
            .O(N__19863),
            .I(\this_sprites_ram.mem_out_bus4_0 ));
    InMux I__3623 (
            .O(N__19860),
            .I(N__19857));
    LocalMux I__3622 (
            .O(N__19857),
            .I(N__19854));
    Span4Mux_h I__3621 (
            .O(N__19854),
            .I(N__19851));
    Span4Mux_h I__3620 (
            .O(N__19851),
            .I(N__19848));
    Span4Mux_v I__3619 (
            .O(N__19848),
            .I(N__19845));
    Odrv4 I__3618 (
            .O(N__19845),
            .I(\this_sprites_ram.mem_out_bus0_0 ));
    InMux I__3617 (
            .O(N__19842),
            .I(N__19838));
    InMux I__3616 (
            .O(N__19841),
            .I(N__19835));
    LocalMux I__3615 (
            .O(N__19838),
            .I(N__19832));
    LocalMux I__3614 (
            .O(N__19835),
            .I(N__19829));
    Odrv12 I__3613 (
            .O(N__19832),
            .I(\this_ppu.vram_en_i_a2Z0Z_0 ));
    Odrv4 I__3612 (
            .O(N__19829),
            .I(\this_ppu.vram_en_i_a2Z0Z_0 ));
    CascadeMux I__3611 (
            .O(N__19824),
            .I(\this_ppu.vram_en_i_a2Z0Z_0_cascade_ ));
    CascadeMux I__3610 (
            .O(N__19821),
            .I(M_this_ppu_vram_en_0_cascade_));
    CascadeMux I__3609 (
            .O(N__19818),
            .I(\this_ppu.un1_M_haddress_q_3_c2_cascade_ ));
    InMux I__3608 (
            .O(N__19815),
            .I(N__19812));
    LocalMux I__3607 (
            .O(N__19812),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ));
    InMux I__3606 (
            .O(N__19809),
            .I(N__19806));
    LocalMux I__3605 (
            .O(N__19806),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2 ));
    InMux I__3604 (
            .O(N__19803),
            .I(N__19800));
    LocalMux I__3603 (
            .O(N__19800),
            .I(N__19797));
    Span12Mux_h I__3602 (
            .O(N__19797),
            .I(N__19793));
    InMux I__3601 (
            .O(N__19796),
            .I(N__19790));
    Odrv12 I__3600 (
            .O(N__19793),
            .I(M_this_ppu_vram_data_2));
    LocalMux I__3599 (
            .O(N__19790),
            .I(M_this_ppu_vram_data_2));
    InMux I__3598 (
            .O(N__19785),
            .I(N__19782));
    LocalMux I__3597 (
            .O(N__19782),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ));
    InMux I__3596 (
            .O(N__19779),
            .I(N__19776));
    LocalMux I__3595 (
            .O(N__19776),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ));
    InMux I__3594 (
            .O(N__19773),
            .I(N__19770));
    LocalMux I__3593 (
            .O(N__19770),
            .I(N__19767));
    Span4Mux_h I__3592 (
            .O(N__19767),
            .I(N__19764));
    Odrv4 I__3591 (
            .O(N__19764),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ));
    CascadeMux I__3590 (
            .O(N__19761),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_ ));
    InMux I__3589 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__3588 (
            .O(N__19755),
            .I(N__19752));
    Span12Mux_h I__3587 (
            .O(N__19752),
            .I(N__19748));
    InMux I__3586 (
            .O(N__19751),
            .I(N__19745));
    Odrv12 I__3585 (
            .O(N__19748),
            .I(M_this_ppu_vram_data_0));
    LocalMux I__3584 (
            .O(N__19745),
            .I(M_this_ppu_vram_data_0));
    InMux I__3583 (
            .O(N__19740),
            .I(N__19737));
    LocalMux I__3582 (
            .O(N__19737),
            .I(\this_ppu.N_124 ));
    CascadeMux I__3581 (
            .O(N__19734),
            .I(\this_ppu.N_124_cascade_ ));
    CascadeMux I__3580 (
            .O(N__19731),
            .I(\this_ppu.un1_M_vaddress_q_2_c5_cascade_ ));
    InMux I__3579 (
            .O(N__19728),
            .I(N__19724));
    InMux I__3578 (
            .O(N__19727),
            .I(N__19721));
    LocalMux I__3577 (
            .O(N__19724),
            .I(\this_ppu.un1_M_vaddress_q_2_c5 ));
    LocalMux I__3576 (
            .O(N__19721),
            .I(\this_ppu.un1_M_vaddress_q_2_c5 ));
    InMux I__3575 (
            .O(N__19716),
            .I(N__19712));
    InMux I__3574 (
            .O(N__19715),
            .I(N__19706));
    LocalMux I__3573 (
            .O(N__19712),
            .I(N__19703));
    InMux I__3572 (
            .O(N__19711),
            .I(N__19696));
    InMux I__3571 (
            .O(N__19710),
            .I(N__19696));
    InMux I__3570 (
            .O(N__19709),
            .I(N__19696));
    LocalMux I__3569 (
            .O(N__19706),
            .I(\this_ppu.M_last_q ));
    Odrv4 I__3568 (
            .O(N__19703),
            .I(\this_ppu.M_last_q ));
    LocalMux I__3567 (
            .O(N__19696),
            .I(\this_ppu.M_last_q ));
    CascadeMux I__3566 (
            .O(N__19689),
            .I(N__19685));
    CascadeMux I__3565 (
            .O(N__19688),
            .I(N__19680));
    InMux I__3564 (
            .O(N__19685),
            .I(N__19677));
    CascadeMux I__3563 (
            .O(N__19684),
            .I(N__19674));
    InMux I__3562 (
            .O(N__19683),
            .I(N__19665));
    InMux I__3561 (
            .O(N__19680),
            .I(N__19665));
    LocalMux I__3560 (
            .O(N__19677),
            .I(N__19662));
    InMux I__3559 (
            .O(N__19674),
            .I(N__19655));
    InMux I__3558 (
            .O(N__19673),
            .I(N__19655));
    InMux I__3557 (
            .O(N__19672),
            .I(N__19655));
    CascadeMux I__3556 (
            .O(N__19671),
            .I(N__19652));
    InMux I__3555 (
            .O(N__19670),
            .I(N__19649));
    LocalMux I__3554 (
            .O(N__19665),
            .I(N__19642));
    Span4Mux_h I__3553 (
            .O(N__19662),
            .I(N__19642));
    LocalMux I__3552 (
            .O(N__19655),
            .I(N__19642));
    InMux I__3551 (
            .O(N__19652),
            .I(N__19639));
    LocalMux I__3550 (
            .O(N__19649),
            .I(N__19636));
    Span4Mux_h I__3549 (
            .O(N__19642),
            .I(N__19633));
    LocalMux I__3548 (
            .O(N__19639),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv12 I__3547 (
            .O(N__19636),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv4 I__3546 (
            .O(N__19633),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    InMux I__3545 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__3544 (
            .O(N__19623),
            .I(N__19620));
    Odrv4 I__3543 (
            .O(N__19620),
            .I(N_1318_tz_0));
    InMux I__3542 (
            .O(N__19617),
            .I(N__19614));
    LocalMux I__3541 (
            .O(N__19614),
            .I(\this_ppu.M_this_oam_ram_read_data_i_16 ));
    InMux I__3540 (
            .O(N__19611),
            .I(N__19608));
    LocalMux I__3539 (
            .O(N__19608),
            .I(N__19605));
    Odrv4 I__3538 (
            .O(N__19605),
            .I(\this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ));
    InMux I__3537 (
            .O(N__19602),
            .I(\this_ppu.un2_vscroll_cry_0 ));
    InMux I__3536 (
            .O(N__19599),
            .I(\this_ppu.un2_vscroll_cry_1 ));
    InMux I__3535 (
            .O(N__19596),
            .I(N__19593));
    LocalMux I__3534 (
            .O(N__19593),
            .I(\this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ));
    InMux I__3533 (
            .O(N__19590),
            .I(N__19587));
    LocalMux I__3532 (
            .O(N__19587),
            .I(M_this_oam_ram_read_data_i_17));
    CascadeMux I__3531 (
            .O(N__19584),
            .I(N__19581));
    InMux I__3530 (
            .O(N__19581),
            .I(N__19578));
    LocalMux I__3529 (
            .O(N__19578),
            .I(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_5));
    CascadeMux I__3528 (
            .O(N__19575),
            .I(\this_vga_signals.N_659_cascade_ ));
    CascadeMux I__3527 (
            .O(N__19572),
            .I(N_572_cascade_));
    InMux I__3526 (
            .O(N__19569),
            .I(N__19566));
    LocalMux I__3525 (
            .O(N__19566),
            .I(M_this_sprites_address_qc_2_0));
    CascadeMux I__3524 (
            .O(N__19563),
            .I(N__19560));
    InMux I__3523 (
            .O(N__19560),
            .I(N__19557));
    LocalMux I__3522 (
            .O(N__19557),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_2 ));
    InMux I__3521 (
            .O(N__19554),
            .I(N__19551));
    LocalMux I__3520 (
            .O(N__19551),
            .I(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_3));
    InMux I__3519 (
            .O(N__19548),
            .I(N__19545));
    LocalMux I__3518 (
            .O(N__19545),
            .I(M_this_sprites_address_q_0_0_i_484));
    CascadeMux I__3517 (
            .O(N__19542),
            .I(M_this_sprites_address_qc_3_0_cascade_));
    CascadeMux I__3516 (
            .O(N__19539),
            .I(N__19536));
    InMux I__3515 (
            .O(N__19536),
            .I(N__19533));
    LocalMux I__3514 (
            .O(N__19533),
            .I(M_this_substate_q_s_1));
    CascadeMux I__3513 (
            .O(N__19530),
            .I(M_this_sprites_address_q_0_0_i_480_cascade_));
    InMux I__3512 (
            .O(N__19527),
            .I(N__19524));
    LocalMux I__3511 (
            .O(N__19524),
            .I(M_this_sprites_address_qc_4_0));
    InMux I__3510 (
            .O(N__19521),
            .I(N__19518));
    LocalMux I__3509 (
            .O(N__19518),
            .I(N_511_1));
    InMux I__3508 (
            .O(N__19515),
            .I(N__19512));
    LocalMux I__3507 (
            .O(N__19512),
            .I(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_4));
    CascadeMux I__3506 (
            .O(N__19509),
            .I(N__19502));
    InMux I__3505 (
            .O(N__19508),
            .I(N__19492));
    InMux I__3504 (
            .O(N__19507),
            .I(N__19492));
    InMux I__3503 (
            .O(N__19506),
            .I(N__19492));
    InMux I__3502 (
            .O(N__19505),
            .I(N__19492));
    InMux I__3501 (
            .O(N__19502),
            .I(N__19487));
    InMux I__3500 (
            .O(N__19501),
            .I(N__19487));
    LocalMux I__3499 (
            .O(N__19492),
            .I(N__19481));
    LocalMux I__3498 (
            .O(N__19487),
            .I(N__19478));
    InMux I__3497 (
            .O(N__19486),
            .I(N__19475));
    InMux I__3496 (
            .O(N__19485),
            .I(N__19470));
    InMux I__3495 (
            .O(N__19484),
            .I(N__19470));
    Span12Mux_v I__3494 (
            .O(N__19481),
            .I(N__19462));
    Sp12to4 I__3493 (
            .O(N__19478),
            .I(N__19462));
    LocalMux I__3492 (
            .O(N__19475),
            .I(N__19462));
    LocalMux I__3491 (
            .O(N__19470),
            .I(N__19459));
    InMux I__3490 (
            .O(N__19469),
            .I(N__19456));
    Span12Mux_v I__3489 (
            .O(N__19462),
            .I(N__19453));
    Span12Mux_v I__3488 (
            .O(N__19459),
            .I(N__19450));
    LocalMux I__3487 (
            .O(N__19456),
            .I(N__19447));
    Odrv12 I__3486 (
            .O(N__19453),
            .I(rst_n_c));
    Odrv12 I__3485 (
            .O(N__19450),
            .I(rst_n_c));
    Odrv12 I__3484 (
            .O(N__19447),
            .I(rst_n_c));
    InMux I__3483 (
            .O(N__19440),
            .I(N__19437));
    LocalMux I__3482 (
            .O(N__19437),
            .I(\this_reset_cond.M_stage_qZ0Z_4 ));
    InMux I__3481 (
            .O(N__19434),
            .I(N__19431));
    LocalMux I__3480 (
            .O(N__19431),
            .I(\this_reset_cond.M_stage_qZ0Z_5 ));
    InMux I__3479 (
            .O(N__19428),
            .I(N__19425));
    LocalMux I__3478 (
            .O(N__19425),
            .I(N__19422));
    Span4Mux_h I__3477 (
            .O(N__19422),
            .I(N__19419));
    Span4Mux_v I__3476 (
            .O(N__19419),
            .I(N__19416));
    Span4Mux_h I__3475 (
            .O(N__19416),
            .I(N__19413));
    Odrv4 I__3474 (
            .O(N__19413),
            .I(\this_sprites_ram.mem_out_bus6_0 ));
    InMux I__3473 (
            .O(N__19410),
            .I(N__19407));
    LocalMux I__3472 (
            .O(N__19407),
            .I(N__19404));
    Span4Mux_v I__3471 (
            .O(N__19404),
            .I(N__19401));
    Sp12to4 I__3470 (
            .O(N__19401),
            .I(N__19398));
    Odrv12 I__3469 (
            .O(N__19398),
            .I(\this_sprites_ram.mem_out_bus2_0 ));
    InMux I__3468 (
            .O(N__19395),
            .I(N__19392));
    LocalMux I__3467 (
            .O(N__19392),
            .I(N__19389));
    Span4Mux_v I__3466 (
            .O(N__19389),
            .I(N__19386));
    Span4Mux_v I__3465 (
            .O(N__19386),
            .I(N__19383));
    Span4Mux_h I__3464 (
            .O(N__19383),
            .I(N__19380));
    Span4Mux_h I__3463 (
            .O(N__19380),
            .I(N__19377));
    Odrv4 I__3462 (
            .O(N__19377),
            .I(M_this_map_ram_read_data_5));
    CascadeMux I__3461 (
            .O(N__19374),
            .I(N__19371));
    InMux I__3460 (
            .O(N__19371),
            .I(N__19368));
    LocalMux I__3459 (
            .O(N__19368),
            .I(N__19365));
    Span4Mux_v I__3458 (
            .O(N__19365),
            .I(N__19362));
    Sp12to4 I__3457 (
            .O(N__19362),
            .I(N__19359));
    Span12Mux_h I__3456 (
            .O(N__19359),
            .I(N__19356));
    Odrv12 I__3455 (
            .O(N__19356),
            .I(M_this_oam_ram_read_data_5));
    InMux I__3454 (
            .O(N__19353),
            .I(N__19350));
    LocalMux I__3453 (
            .O(N__19350),
            .I(N__19347));
    Span4Mux_h I__3452 (
            .O(N__19347),
            .I(N__19344));
    Sp12to4 I__3451 (
            .O(N__19344),
            .I(N__19341));
    Span12Mux_v I__3450 (
            .O(N__19341),
            .I(N__19338));
    Odrv12 I__3449 (
            .O(N__19338),
            .I(M_this_map_ram_read_data_7));
    CascadeMux I__3448 (
            .O(N__19335),
            .I(N__19332));
    InMux I__3447 (
            .O(N__19332),
            .I(N__19329));
    LocalMux I__3446 (
            .O(N__19329),
            .I(N__19326));
    Span4Mux_v I__3445 (
            .O(N__19326),
            .I(N__19323));
    Span4Mux_h I__3444 (
            .O(N__19323),
            .I(N__19320));
    Sp12to4 I__3443 (
            .O(N__19320),
            .I(N__19317));
    Span12Mux_v I__3442 (
            .O(N__19317),
            .I(N__19314));
    Odrv12 I__3441 (
            .O(N__19314),
            .I(M_this_oam_ram_read_data_7));
    InMux I__3440 (
            .O(N__19311),
            .I(N__19308));
    LocalMux I__3439 (
            .O(N__19308),
            .I(N__19305));
    Sp12to4 I__3438 (
            .O(N__19305),
            .I(N__19302));
    Span12Mux_v I__3437 (
            .O(N__19302),
            .I(N__19299));
    Odrv12 I__3436 (
            .O(N__19299),
            .I(\this_sprites_ram.mem_out_bus4_2 ));
    InMux I__3435 (
            .O(N__19296),
            .I(N__19293));
    LocalMux I__3434 (
            .O(N__19293),
            .I(N__19290));
    Span12Mux_v I__3433 (
            .O(N__19290),
            .I(N__19287));
    Odrv12 I__3432 (
            .O(N__19287),
            .I(\this_sprites_ram.mem_out_bus0_2 ));
    CascadeMux I__3431 (
            .O(N__19284),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ));
    InMux I__3430 (
            .O(N__19281),
            .I(N__19278));
    LocalMux I__3429 (
            .O(N__19278),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ));
    InMux I__3428 (
            .O(N__19275),
            .I(N__19272));
    LocalMux I__3427 (
            .O(N__19272),
            .I(N__19269));
    Span4Mux_v I__3426 (
            .O(N__19269),
            .I(N__19266));
    Span4Mux_h I__3425 (
            .O(N__19266),
            .I(N__19263));
    Span4Mux_h I__3424 (
            .O(N__19263),
            .I(N__19260));
    Span4Mux_v I__3423 (
            .O(N__19260),
            .I(N__19257));
    Span4Mux_v I__3422 (
            .O(N__19257),
            .I(N__19254));
    Odrv4 I__3421 (
            .O(N__19254),
            .I(M_this_oam_ram_read_data_3));
    InMux I__3420 (
            .O(N__19251),
            .I(N__19248));
    LocalMux I__3419 (
            .O(N__19248),
            .I(N__19245));
    Span4Mux_v I__3418 (
            .O(N__19245),
            .I(N__19242));
    Sp12to4 I__3417 (
            .O(N__19242),
            .I(N__19239));
    Span12Mux_h I__3416 (
            .O(N__19239),
            .I(N__19236));
    Odrv12 I__3415 (
            .O(N__19236),
            .I(M_this_map_ram_read_data_3));
    CascadeMux I__3414 (
            .O(N__19233),
            .I(N__19225));
    CascadeMux I__3413 (
            .O(N__19232),
            .I(N__19222));
    CascadeMux I__3412 (
            .O(N__19231),
            .I(N__19219));
    CascadeMux I__3411 (
            .O(N__19230),
            .I(N__19216));
    CascadeMux I__3410 (
            .O(N__19229),
            .I(N__19209));
    CascadeMux I__3409 (
            .O(N__19228),
            .I(N__19206));
    InMux I__3408 (
            .O(N__19225),
            .I(N__19203));
    InMux I__3407 (
            .O(N__19222),
            .I(N__19200));
    InMux I__3406 (
            .O(N__19219),
            .I(N__19197));
    InMux I__3405 (
            .O(N__19216),
            .I(N__19194));
    CascadeMux I__3404 (
            .O(N__19215),
            .I(N__19190));
    CascadeMux I__3403 (
            .O(N__19214),
            .I(N__19187));
    CascadeMux I__3402 (
            .O(N__19213),
            .I(N__19184));
    CascadeMux I__3401 (
            .O(N__19212),
            .I(N__19178));
    InMux I__3400 (
            .O(N__19209),
            .I(N__19175));
    InMux I__3399 (
            .O(N__19206),
            .I(N__19172));
    LocalMux I__3398 (
            .O(N__19203),
            .I(N__19169));
    LocalMux I__3397 (
            .O(N__19200),
            .I(N__19166));
    LocalMux I__3396 (
            .O(N__19197),
            .I(N__19162));
    LocalMux I__3395 (
            .O(N__19194),
            .I(N__19159));
    CascadeMux I__3394 (
            .O(N__19193),
            .I(N__19156));
    InMux I__3393 (
            .O(N__19190),
            .I(N__19153));
    InMux I__3392 (
            .O(N__19187),
            .I(N__19150));
    InMux I__3391 (
            .O(N__19184),
            .I(N__19147));
    CascadeMux I__3390 (
            .O(N__19183),
            .I(N__19143));
    CascadeMux I__3389 (
            .O(N__19182),
            .I(N__19140));
    CascadeMux I__3388 (
            .O(N__19181),
            .I(N__19137));
    InMux I__3387 (
            .O(N__19178),
            .I(N__19134));
    LocalMux I__3386 (
            .O(N__19175),
            .I(N__19127));
    LocalMux I__3385 (
            .O(N__19172),
            .I(N__19127));
    Span4Mux_v I__3384 (
            .O(N__19169),
            .I(N__19127));
    Span4Mux_h I__3383 (
            .O(N__19166),
            .I(N__19124));
    CascadeMux I__3382 (
            .O(N__19165),
            .I(N__19121));
    Span4Mux_h I__3381 (
            .O(N__19162),
            .I(N__19118));
    Span4Mux_h I__3380 (
            .O(N__19159),
            .I(N__19115));
    InMux I__3379 (
            .O(N__19156),
            .I(N__19112));
    LocalMux I__3378 (
            .O(N__19153),
            .I(N__19109));
    LocalMux I__3377 (
            .O(N__19150),
            .I(N__19106));
    LocalMux I__3376 (
            .O(N__19147),
            .I(N__19103));
    CascadeMux I__3375 (
            .O(N__19146),
            .I(N__19100));
    InMux I__3374 (
            .O(N__19143),
            .I(N__19097));
    InMux I__3373 (
            .O(N__19140),
            .I(N__19094));
    InMux I__3372 (
            .O(N__19137),
            .I(N__19091));
    LocalMux I__3371 (
            .O(N__19134),
            .I(N__19088));
    Span4Mux_v I__3370 (
            .O(N__19127),
            .I(N__19085));
    Span4Mux_v I__3369 (
            .O(N__19124),
            .I(N__19082));
    InMux I__3368 (
            .O(N__19121),
            .I(N__19079));
    Span4Mux_h I__3367 (
            .O(N__19118),
            .I(N__19076));
    Span4Mux_h I__3366 (
            .O(N__19115),
            .I(N__19073));
    LocalMux I__3365 (
            .O(N__19112),
            .I(N__19070));
    Span4Mux_h I__3364 (
            .O(N__19109),
            .I(N__19067));
    Span4Mux_h I__3363 (
            .O(N__19106),
            .I(N__19064));
    Span4Mux_h I__3362 (
            .O(N__19103),
            .I(N__19061));
    InMux I__3361 (
            .O(N__19100),
            .I(N__19058));
    LocalMux I__3360 (
            .O(N__19097),
            .I(N__19055));
    LocalMux I__3359 (
            .O(N__19094),
            .I(N__19052));
    LocalMux I__3358 (
            .O(N__19091),
            .I(N__19049));
    Span4Mux_h I__3357 (
            .O(N__19088),
            .I(N__19046));
    Span4Mux_h I__3356 (
            .O(N__19085),
            .I(N__19041));
    Span4Mux_v I__3355 (
            .O(N__19082),
            .I(N__19041));
    LocalMux I__3354 (
            .O(N__19079),
            .I(N__19038));
    Sp12to4 I__3353 (
            .O(N__19076),
            .I(N__19031));
    Sp12to4 I__3352 (
            .O(N__19073),
            .I(N__19031));
    Span12Mux_h I__3351 (
            .O(N__19070),
            .I(N__19031));
    Span4Mux_v I__3350 (
            .O(N__19067),
            .I(N__19028));
    Sp12to4 I__3349 (
            .O(N__19064),
            .I(N__19023));
    Sp12to4 I__3348 (
            .O(N__19061),
            .I(N__19023));
    LocalMux I__3347 (
            .O(N__19058),
            .I(N__19020));
    Span12Mux_h I__3346 (
            .O(N__19055),
            .I(N__19013));
    Span12Mux_h I__3345 (
            .O(N__19052),
            .I(N__19013));
    Span12Mux_h I__3344 (
            .O(N__19049),
            .I(N__19013));
    Span4Mux_h I__3343 (
            .O(N__19046),
            .I(N__19008));
    Span4Mux_h I__3342 (
            .O(N__19041),
            .I(N__19008));
    Sp12to4 I__3341 (
            .O(N__19038),
            .I(N__18999));
    Span12Mux_v I__3340 (
            .O(N__19031),
            .I(N__18999));
    Sp12to4 I__3339 (
            .O(N__19028),
            .I(N__18999));
    Span12Mux_v I__3338 (
            .O(N__19023),
            .I(N__18999));
    Odrv12 I__3337 (
            .O(N__19020),
            .I(M_this_ppu_sprites_addr_9));
    Odrv12 I__3336 (
            .O(N__19013),
            .I(M_this_ppu_sprites_addr_9));
    Odrv4 I__3335 (
            .O(N__19008),
            .I(M_this_ppu_sprites_addr_9));
    Odrv12 I__3334 (
            .O(N__18999),
            .I(M_this_ppu_sprites_addr_9));
    InMux I__3333 (
            .O(N__18990),
            .I(N__18987));
    LocalMux I__3332 (
            .O(N__18987),
            .I(N__18984));
    Span4Mux_v I__3331 (
            .O(N__18984),
            .I(N__18981));
    Span4Mux_h I__3330 (
            .O(N__18981),
            .I(N__18978));
    Odrv4 I__3329 (
            .O(N__18978),
            .I(\this_sprites_ram.mem_out_bus7_2 ));
    InMux I__3328 (
            .O(N__18975),
            .I(N__18972));
    LocalMux I__3327 (
            .O(N__18972),
            .I(N__18969));
    Span4Mux_v I__3326 (
            .O(N__18969),
            .I(N__18966));
    Span4Mux_h I__3325 (
            .O(N__18966),
            .I(N__18963));
    Span4Mux_h I__3324 (
            .O(N__18963),
            .I(N__18960));
    Odrv4 I__3323 (
            .O(N__18960),
            .I(\this_sprites_ram.mem_out_bus3_2 ));
    InMux I__3322 (
            .O(N__18957),
            .I(N__18954));
    LocalMux I__3321 (
            .O(N__18954),
            .I(\this_reset_cond.M_stage_qZ0Z_8 ));
    InMux I__3320 (
            .O(N__18951),
            .I(N__18947));
    InMux I__3319 (
            .O(N__18950),
            .I(N__18941));
    LocalMux I__3318 (
            .O(N__18947),
            .I(N__18938));
    InMux I__3317 (
            .O(N__18946),
            .I(N__18935));
    InMux I__3316 (
            .O(N__18945),
            .I(N__18932));
    InMux I__3315 (
            .O(N__18944),
            .I(N__18929));
    LocalMux I__3314 (
            .O(N__18941),
            .I(N__18922));
    Span4Mux_h I__3313 (
            .O(N__18938),
            .I(N__18922));
    LocalMux I__3312 (
            .O(N__18935),
            .I(N__18922));
    LocalMux I__3311 (
            .O(N__18932),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    LocalMux I__3310 (
            .O(N__18929),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv4 I__3309 (
            .O(N__18922),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    InMux I__3308 (
            .O(N__18915),
            .I(N__18912));
    LocalMux I__3307 (
            .O(N__18912),
            .I(N__18909));
    Odrv4 I__3306 (
            .O(N__18909),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5 ));
    InMux I__3305 (
            .O(N__18906),
            .I(N__18902));
    InMux I__3304 (
            .O(N__18905),
            .I(N__18899));
    LocalMux I__3303 (
            .O(N__18902),
            .I(N__18896));
    LocalMux I__3302 (
            .O(N__18899),
            .I(N__18893));
    Span4Mux_v I__3301 (
            .O(N__18896),
            .I(N__18890));
    Span4Mux_h I__3300 (
            .O(N__18893),
            .I(N__18887));
    Odrv4 I__3299 (
            .O(N__18890),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4 ));
    Odrv4 I__3298 (
            .O(N__18887),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4 ));
    InMux I__3297 (
            .O(N__18882),
            .I(N__18878));
    InMux I__3296 (
            .O(N__18881),
            .I(N__18875));
    LocalMux I__3295 (
            .O(N__18878),
            .I(N__18872));
    LocalMux I__3294 (
            .O(N__18875),
            .I(N__18869));
    Odrv4 I__3293 (
            .O(N__18872),
            .I(\this_ppu.M_count_d_0_sqmuxa_1 ));
    Odrv4 I__3292 (
            .O(N__18869),
            .I(\this_ppu.M_count_d_0_sqmuxa_1 ));
    CascadeMux I__3291 (
            .O(N__18864),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_cascade_ ));
    InMux I__3290 (
            .O(N__18861),
            .I(N__18858));
    LocalMux I__3289 (
            .O(N__18858),
            .I(N__18853));
    InMux I__3288 (
            .O(N__18857),
            .I(N__18850));
    InMux I__3287 (
            .O(N__18856),
            .I(N__18846));
    Span4Mux_h I__3286 (
            .O(N__18853),
            .I(N__18841));
    LocalMux I__3285 (
            .O(N__18850),
            .I(N__18841));
    InMux I__3284 (
            .O(N__18849),
            .I(N__18838));
    LocalMux I__3283 (
            .O(N__18846),
            .I(\this_ppu.M_line_clk_out_0 ));
    Odrv4 I__3282 (
            .O(N__18841),
            .I(\this_ppu.M_line_clk_out_0 ));
    LocalMux I__3281 (
            .O(N__18838),
            .I(\this_ppu.M_line_clk_out_0 ));
    InMux I__3280 (
            .O(N__18831),
            .I(N__18823));
    InMux I__3279 (
            .O(N__18830),
            .I(N__18816));
    InMux I__3278 (
            .O(N__18829),
            .I(N__18816));
    InMux I__3277 (
            .O(N__18828),
            .I(N__18816));
    InMux I__3276 (
            .O(N__18827),
            .I(N__18811));
    InMux I__3275 (
            .O(N__18826),
            .I(N__18811));
    LocalMux I__3274 (
            .O(N__18823),
            .I(\this_ppu.N_1417_0 ));
    LocalMux I__3273 (
            .O(N__18816),
            .I(\this_ppu.N_1417_0 ));
    LocalMux I__3272 (
            .O(N__18811),
            .I(\this_ppu.N_1417_0 ));
    InMux I__3271 (
            .O(N__18804),
            .I(N__18801));
    LocalMux I__3270 (
            .O(N__18801),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ));
    CascadeMux I__3269 (
            .O(N__18798),
            .I(\this_ppu.N_1417_0_cascade_ ));
    CascadeMux I__3268 (
            .O(N__18795),
            .I(N__18791));
    CascadeMux I__3267 (
            .O(N__18794),
            .I(N__18788));
    InMux I__3266 (
            .O(N__18791),
            .I(N__18779));
    InMux I__3265 (
            .O(N__18788),
            .I(N__18779));
    InMux I__3264 (
            .O(N__18787),
            .I(N__18779));
    InMux I__3263 (
            .O(N__18786),
            .I(N__18774));
    LocalMux I__3262 (
            .O(N__18779),
            .I(N__18771));
    InMux I__3261 (
            .O(N__18778),
            .I(N__18766));
    InMux I__3260 (
            .O(N__18777),
            .I(N__18766));
    LocalMux I__3259 (
            .O(N__18774),
            .I(\this_ppu.un13_0 ));
    Odrv4 I__3258 (
            .O(N__18771),
            .I(\this_ppu.un13_0 ));
    LocalMux I__3257 (
            .O(N__18766),
            .I(\this_ppu.un13_0 ));
    CascadeMux I__3256 (
            .O(N__18759),
            .I(N__18755));
    InMux I__3255 (
            .O(N__18758),
            .I(N__18752));
    InMux I__3254 (
            .O(N__18755),
            .I(N__18748));
    LocalMux I__3253 (
            .O(N__18752),
            .I(N__18745));
    InMux I__3252 (
            .O(N__18751),
            .I(N__18742));
    LocalMux I__3251 (
            .O(N__18748),
            .I(N__18739));
    Span4Mux_h I__3250 (
            .O(N__18745),
            .I(N__18736));
    LocalMux I__3249 (
            .O(N__18742),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    Odrv4 I__3248 (
            .O(N__18739),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    Odrv4 I__3247 (
            .O(N__18736),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    InMux I__3246 (
            .O(N__18729),
            .I(N__18726));
    LocalMux I__3245 (
            .O(N__18726),
            .I(N__18723));
    Span4Mux_h I__3244 (
            .O(N__18723),
            .I(N__18720));
    Span4Mux_h I__3243 (
            .O(N__18720),
            .I(N__18717));
    Odrv4 I__3242 (
            .O(N__18717),
            .I(\this_sprites_ram.mem_out_bus6_2 ));
    InMux I__3241 (
            .O(N__18714),
            .I(N__18711));
    LocalMux I__3240 (
            .O(N__18711),
            .I(N__18708));
    Span4Mux_h I__3239 (
            .O(N__18708),
            .I(N__18705));
    Span4Mux_h I__3238 (
            .O(N__18705),
            .I(N__18702));
    Span4Mux_h I__3237 (
            .O(N__18702),
            .I(N__18699));
    Odrv4 I__3236 (
            .O(N__18699),
            .I(\this_sprites_ram.mem_out_bus2_2 ));
    InMux I__3235 (
            .O(N__18696),
            .I(N__18693));
    LocalMux I__3234 (
            .O(N__18693),
            .I(N__18690));
    Odrv12 I__3233 (
            .O(N__18690),
            .I(\this_reset_cond.M_stage_qZ0Z_3 ));
    InMux I__3232 (
            .O(N__18687),
            .I(N__18684));
    LocalMux I__3231 (
            .O(N__18684),
            .I(\this_reset_cond.M_stage_qZ0Z_6 ));
    InMux I__3230 (
            .O(N__18681),
            .I(N__18678));
    LocalMux I__3229 (
            .O(N__18678),
            .I(\this_reset_cond.M_stage_qZ0Z_7 ));
    InMux I__3228 (
            .O(N__18675),
            .I(N__18672));
    LocalMux I__3227 (
            .O(N__18672),
            .I(N__18669));
    Odrv4 I__3226 (
            .O(N__18669),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    CascadeMux I__3225 (
            .O(N__18666),
            .I(\this_ppu.M_state_q_srsts_i_2_1_cascade_ ));
    InMux I__3224 (
            .O(N__18663),
            .I(N__18658));
    InMux I__3223 (
            .O(N__18662),
            .I(N__18655));
    InMux I__3222 (
            .O(N__18661),
            .I(N__18652));
    LocalMux I__3221 (
            .O(N__18658),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__3220 (
            .O(N__18655),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__3219 (
            .O(N__18652),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    CascadeMux I__3218 (
            .O(N__18645),
            .I(N__18641));
    CascadeMux I__3217 (
            .O(N__18644),
            .I(N__18638));
    InMux I__3216 (
            .O(N__18641),
            .I(N__18635));
    InMux I__3215 (
            .O(N__18638),
            .I(N__18632));
    LocalMux I__3214 (
            .O(N__18635),
            .I(N__18629));
    LocalMux I__3213 (
            .O(N__18632),
            .I(N__18626));
    Span4Mux_h I__3212 (
            .O(N__18629),
            .I(N__18623));
    Odrv4 I__3211 (
            .O(N__18626),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    Odrv4 I__3210 (
            .O(N__18623),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    CascadeMux I__3209 (
            .O(N__18618),
            .I(\this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5_cascade_ ));
    CascadeMux I__3208 (
            .O(N__18615),
            .I(N__18612));
    InMux I__3207 (
            .O(N__18612),
            .I(N__18609));
    LocalMux I__3206 (
            .O(N__18609),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ));
    CascadeMux I__3205 (
            .O(N__18606),
            .I(N__18601));
    InMux I__3204 (
            .O(N__18605),
            .I(N__18598));
    InMux I__3203 (
            .O(N__18604),
            .I(N__18595));
    InMux I__3202 (
            .O(N__18601),
            .I(N__18592));
    LocalMux I__3201 (
            .O(N__18598),
            .I(N__18589));
    LocalMux I__3200 (
            .O(N__18595),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    LocalMux I__3199 (
            .O(N__18592),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    Odrv4 I__3198 (
            .O(N__18589),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    InMux I__3197 (
            .O(N__18582),
            .I(N__18577));
    InMux I__3196 (
            .O(N__18581),
            .I(N__18574));
    InMux I__3195 (
            .O(N__18580),
            .I(N__18571));
    LocalMux I__3194 (
            .O(N__18577),
            .I(N__18568));
    LocalMux I__3193 (
            .O(N__18574),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    LocalMux I__3192 (
            .O(N__18571),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    Odrv4 I__3191 (
            .O(N__18568),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    InMux I__3190 (
            .O(N__18561),
            .I(N__18558));
    LocalMux I__3189 (
            .O(N__18558),
            .I(M_this_sprites_address_qc_8_0));
    InMux I__3188 (
            .O(N__18555),
            .I(N__18552));
    LocalMux I__3187 (
            .O(N__18552),
            .I(N__18549));
    Span12Mux_s10_h I__3186 (
            .O(N__18549),
            .I(N__18546));
    Odrv12 I__3185 (
            .O(N__18546),
            .I(M_this_map_ram_write_data_3));
    InMux I__3184 (
            .O(N__18543),
            .I(N__18540));
    LocalMux I__3183 (
            .O(N__18540),
            .I(N__18537));
    Span12Mux_h I__3182 (
            .O(N__18537),
            .I(N__18534));
    Odrv12 I__3181 (
            .O(N__18534),
            .I(M_this_oam_ram_read_data_2));
    CascadeMux I__3180 (
            .O(N__18531),
            .I(N__18528));
    InMux I__3179 (
            .O(N__18528),
            .I(N__18525));
    LocalMux I__3178 (
            .O(N__18525),
            .I(N__18522));
    Span4Mux_v I__3177 (
            .O(N__18522),
            .I(N__18519));
    Sp12to4 I__3176 (
            .O(N__18519),
            .I(N__18516));
    Span12Mux_v I__3175 (
            .O(N__18516),
            .I(N__18513));
    Odrv12 I__3174 (
            .O(N__18513),
            .I(M_this_map_ram_read_data_2));
    CascadeMux I__3173 (
            .O(N__18510),
            .I(N__18507));
    InMux I__3172 (
            .O(N__18507),
            .I(N__18502));
    CascadeMux I__3171 (
            .O(N__18506),
            .I(N__18499));
    CascadeMux I__3170 (
            .O(N__18505),
            .I(N__18496));
    LocalMux I__3169 (
            .O(N__18502),
            .I(N__18488));
    InMux I__3168 (
            .O(N__18499),
            .I(N__18485));
    InMux I__3167 (
            .O(N__18496),
            .I(N__18482));
    CascadeMux I__3166 (
            .O(N__18495),
            .I(N__18477));
    CascadeMux I__3165 (
            .O(N__18494),
            .I(N__18474));
    CascadeMux I__3164 (
            .O(N__18493),
            .I(N__18471));
    CascadeMux I__3163 (
            .O(N__18492),
            .I(N__18468));
    CascadeMux I__3162 (
            .O(N__18491),
            .I(N__18461));
    Span4Mux_v I__3161 (
            .O(N__18488),
            .I(N__18452));
    LocalMux I__3160 (
            .O(N__18485),
            .I(N__18452));
    LocalMux I__3159 (
            .O(N__18482),
            .I(N__18452));
    CascadeMux I__3158 (
            .O(N__18481),
            .I(N__18449));
    CascadeMux I__3157 (
            .O(N__18480),
            .I(N__18446));
    InMux I__3156 (
            .O(N__18477),
            .I(N__18443));
    InMux I__3155 (
            .O(N__18474),
            .I(N__18440));
    InMux I__3154 (
            .O(N__18471),
            .I(N__18437));
    InMux I__3153 (
            .O(N__18468),
            .I(N__18434));
    CascadeMux I__3152 (
            .O(N__18467),
            .I(N__18431));
    CascadeMux I__3151 (
            .O(N__18466),
            .I(N__18428));
    CascadeMux I__3150 (
            .O(N__18465),
            .I(N__18425));
    CascadeMux I__3149 (
            .O(N__18464),
            .I(N__18422));
    InMux I__3148 (
            .O(N__18461),
            .I(N__18419));
    CascadeMux I__3147 (
            .O(N__18460),
            .I(N__18416));
    CascadeMux I__3146 (
            .O(N__18459),
            .I(N__18413));
    Span4Mux_v I__3145 (
            .O(N__18452),
            .I(N__18410));
    InMux I__3144 (
            .O(N__18449),
            .I(N__18407));
    InMux I__3143 (
            .O(N__18446),
            .I(N__18404));
    LocalMux I__3142 (
            .O(N__18443),
            .I(N__18395));
    LocalMux I__3141 (
            .O(N__18440),
            .I(N__18395));
    LocalMux I__3140 (
            .O(N__18437),
            .I(N__18395));
    LocalMux I__3139 (
            .O(N__18434),
            .I(N__18395));
    InMux I__3138 (
            .O(N__18431),
            .I(N__18392));
    InMux I__3137 (
            .O(N__18428),
            .I(N__18389));
    InMux I__3136 (
            .O(N__18425),
            .I(N__18386));
    InMux I__3135 (
            .O(N__18422),
            .I(N__18383));
    LocalMux I__3134 (
            .O(N__18419),
            .I(N__18380));
    InMux I__3133 (
            .O(N__18416),
            .I(N__18377));
    InMux I__3132 (
            .O(N__18413),
            .I(N__18374));
    Sp12to4 I__3131 (
            .O(N__18410),
            .I(N__18369));
    LocalMux I__3130 (
            .O(N__18407),
            .I(N__18369));
    LocalMux I__3129 (
            .O(N__18404),
            .I(N__18366));
    Span12Mux_s9_v I__3128 (
            .O(N__18395),
            .I(N__18351));
    LocalMux I__3127 (
            .O(N__18392),
            .I(N__18351));
    LocalMux I__3126 (
            .O(N__18389),
            .I(N__18351));
    LocalMux I__3125 (
            .O(N__18386),
            .I(N__18351));
    LocalMux I__3124 (
            .O(N__18383),
            .I(N__18351));
    Sp12to4 I__3123 (
            .O(N__18380),
            .I(N__18351));
    LocalMux I__3122 (
            .O(N__18377),
            .I(N__18351));
    LocalMux I__3121 (
            .O(N__18374),
            .I(N__18348));
    Span12Mux_h I__3120 (
            .O(N__18369),
            .I(N__18345));
    Span12Mux_s10_v I__3119 (
            .O(N__18366),
            .I(N__18338));
    Span12Mux_v I__3118 (
            .O(N__18351),
            .I(N__18338));
    Span12Mux_s7_h I__3117 (
            .O(N__18348),
            .I(N__18338));
    Odrv12 I__3116 (
            .O(N__18345),
            .I(M_this_ppu_sprites_addr_8));
    Odrv12 I__3115 (
            .O(N__18338),
            .I(M_this_ppu_sprites_addr_8));
    CascadeMux I__3114 (
            .O(N__18333),
            .I(N__18330));
    InMux I__3113 (
            .O(N__18330),
            .I(N__18323));
    CascadeMux I__3112 (
            .O(N__18329),
            .I(N__18320));
    CascadeMux I__3111 (
            .O(N__18328),
            .I(N__18317));
    CascadeMux I__3110 (
            .O(N__18327),
            .I(N__18313));
    CascadeMux I__3109 (
            .O(N__18326),
            .I(N__18309));
    LocalMux I__3108 (
            .O(N__18323),
            .I(N__18304));
    InMux I__3107 (
            .O(N__18320),
            .I(N__18301));
    InMux I__3106 (
            .O(N__18317),
            .I(N__18298));
    CascadeMux I__3105 (
            .O(N__18316),
            .I(N__18295));
    InMux I__3104 (
            .O(N__18313),
            .I(N__18292));
    CascadeMux I__3103 (
            .O(N__18312),
            .I(N__18289));
    InMux I__3102 (
            .O(N__18309),
            .I(N__18285));
    CascadeMux I__3101 (
            .O(N__18308),
            .I(N__18282));
    CascadeMux I__3100 (
            .O(N__18307),
            .I(N__18276));
    Span4Mux_v I__3099 (
            .O(N__18304),
            .I(N__18267));
    LocalMux I__3098 (
            .O(N__18301),
            .I(N__18267));
    LocalMux I__3097 (
            .O(N__18298),
            .I(N__18267));
    InMux I__3096 (
            .O(N__18295),
            .I(N__18264));
    LocalMux I__3095 (
            .O(N__18292),
            .I(N__18261));
    InMux I__3094 (
            .O(N__18289),
            .I(N__18258));
    CascadeMux I__3093 (
            .O(N__18288),
            .I(N__18255));
    LocalMux I__3092 (
            .O(N__18285),
            .I(N__18252));
    InMux I__3091 (
            .O(N__18282),
            .I(N__18249));
    CascadeMux I__3090 (
            .O(N__18281),
            .I(N__18246));
    CascadeMux I__3089 (
            .O(N__18280),
            .I(N__18243));
    CascadeMux I__3088 (
            .O(N__18279),
            .I(N__18240));
    InMux I__3087 (
            .O(N__18276),
            .I(N__18237));
    CascadeMux I__3086 (
            .O(N__18275),
            .I(N__18234));
    CascadeMux I__3085 (
            .O(N__18274),
            .I(N__18231));
    Span4Mux_v I__3084 (
            .O(N__18267),
            .I(N__18226));
    LocalMux I__3083 (
            .O(N__18264),
            .I(N__18226));
    Span4Mux_v I__3082 (
            .O(N__18261),
            .I(N__18221));
    LocalMux I__3081 (
            .O(N__18258),
            .I(N__18221));
    InMux I__3080 (
            .O(N__18255),
            .I(N__18218));
    Span4Mux_v I__3079 (
            .O(N__18252),
            .I(N__18213));
    LocalMux I__3078 (
            .O(N__18249),
            .I(N__18213));
    InMux I__3077 (
            .O(N__18246),
            .I(N__18210));
    InMux I__3076 (
            .O(N__18243),
            .I(N__18207));
    InMux I__3075 (
            .O(N__18240),
            .I(N__18204));
    LocalMux I__3074 (
            .O(N__18237),
            .I(N__18201));
    InMux I__3073 (
            .O(N__18234),
            .I(N__18198));
    InMux I__3072 (
            .O(N__18231),
            .I(N__18195));
    Span4Mux_v I__3071 (
            .O(N__18226),
            .I(N__18191));
    Span4Mux_v I__3070 (
            .O(N__18221),
            .I(N__18188));
    LocalMux I__3069 (
            .O(N__18218),
            .I(N__18185));
    Span4Mux_v I__3068 (
            .O(N__18213),
            .I(N__18178));
    LocalMux I__3067 (
            .O(N__18210),
            .I(N__18178));
    LocalMux I__3066 (
            .O(N__18207),
            .I(N__18178));
    LocalMux I__3065 (
            .O(N__18204),
            .I(N__18175));
    Span4Mux_v I__3064 (
            .O(N__18201),
            .I(N__18168));
    LocalMux I__3063 (
            .O(N__18198),
            .I(N__18168));
    LocalMux I__3062 (
            .O(N__18195),
            .I(N__18168));
    CascadeMux I__3061 (
            .O(N__18194),
            .I(N__18165));
    Span4Mux_v I__3060 (
            .O(N__18191),
            .I(N__18162));
    Sp12to4 I__3059 (
            .O(N__18188),
            .I(N__18155));
    Span12Mux_h I__3058 (
            .O(N__18185),
            .I(N__18155));
    Sp12to4 I__3057 (
            .O(N__18178),
            .I(N__18155));
    Span4Mux_v I__3056 (
            .O(N__18175),
            .I(N__18150));
    Span4Mux_v I__3055 (
            .O(N__18168),
            .I(N__18150));
    InMux I__3054 (
            .O(N__18165),
            .I(N__18147));
    Sp12to4 I__3053 (
            .O(N__18162),
            .I(N__18144));
    Span12Mux_v I__3052 (
            .O(N__18155),
            .I(N__18137));
    Sp12to4 I__3051 (
            .O(N__18150),
            .I(N__18137));
    LocalMux I__3050 (
            .O(N__18147),
            .I(N__18137));
    Odrv12 I__3049 (
            .O(N__18144),
            .I(M_this_ppu_sprites_addr_5));
    Odrv12 I__3048 (
            .O(N__18137),
            .I(M_this_ppu_sprites_addr_5));
    InMux I__3047 (
            .O(N__18132),
            .I(N__18129));
    LocalMux I__3046 (
            .O(N__18129),
            .I(N__18126));
    Odrv4 I__3045 (
            .O(N__18126),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__3044 (
            .O(N__18123),
            .I(N__18120));
    LocalMux I__3043 (
            .O(N__18120),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    CascadeMux I__3042 (
            .O(N__18117),
            .I(N__18107));
    CascadeMux I__3041 (
            .O(N__18116),
            .I(N__18103));
    CascadeMux I__3040 (
            .O(N__18115),
            .I(N__18095));
    CascadeMux I__3039 (
            .O(N__18114),
            .I(N__18091));
    CascadeMux I__3038 (
            .O(N__18113),
            .I(N__18088));
    CascadeMux I__3037 (
            .O(N__18112),
            .I(N__18085));
    CascadeMux I__3036 (
            .O(N__18111),
            .I(N__18082));
    CascadeMux I__3035 (
            .O(N__18110),
            .I(N__18079));
    InMux I__3034 (
            .O(N__18107),
            .I(N__18076));
    CascadeMux I__3033 (
            .O(N__18106),
            .I(N__18073));
    InMux I__3032 (
            .O(N__18103),
            .I(N__18070));
    CascadeMux I__3031 (
            .O(N__18102),
            .I(N__18067));
    CascadeMux I__3030 (
            .O(N__18101),
            .I(N__18064));
    CascadeMux I__3029 (
            .O(N__18100),
            .I(N__18061));
    CascadeMux I__3028 (
            .O(N__18099),
            .I(N__18058));
    CascadeMux I__3027 (
            .O(N__18098),
            .I(N__18055));
    InMux I__3026 (
            .O(N__18095),
            .I(N__18052));
    CascadeMux I__3025 (
            .O(N__18094),
            .I(N__18049));
    InMux I__3024 (
            .O(N__18091),
            .I(N__18046));
    InMux I__3023 (
            .O(N__18088),
            .I(N__18043));
    InMux I__3022 (
            .O(N__18085),
            .I(N__18040));
    InMux I__3021 (
            .O(N__18082),
            .I(N__18037));
    InMux I__3020 (
            .O(N__18079),
            .I(N__18034));
    LocalMux I__3019 (
            .O(N__18076),
            .I(N__18031));
    InMux I__3018 (
            .O(N__18073),
            .I(N__18028));
    LocalMux I__3017 (
            .O(N__18070),
            .I(N__18025));
    InMux I__3016 (
            .O(N__18067),
            .I(N__18021));
    InMux I__3015 (
            .O(N__18064),
            .I(N__18018));
    InMux I__3014 (
            .O(N__18061),
            .I(N__18015));
    InMux I__3013 (
            .O(N__18058),
            .I(N__18012));
    InMux I__3012 (
            .O(N__18055),
            .I(N__18009));
    LocalMux I__3011 (
            .O(N__18052),
            .I(N__18006));
    InMux I__3010 (
            .O(N__18049),
            .I(N__18003));
    LocalMux I__3009 (
            .O(N__18046),
            .I(N__17998));
    LocalMux I__3008 (
            .O(N__18043),
            .I(N__17998));
    LocalMux I__3007 (
            .O(N__18040),
            .I(N__17995));
    LocalMux I__3006 (
            .O(N__18037),
            .I(N__17992));
    LocalMux I__3005 (
            .O(N__18034),
            .I(N__17985));
    Span4Mux_v I__3004 (
            .O(N__18031),
            .I(N__17985));
    LocalMux I__3003 (
            .O(N__18028),
            .I(N__17985));
    Span4Mux_v I__3002 (
            .O(N__18025),
            .I(N__17982));
    CascadeMux I__3001 (
            .O(N__18024),
            .I(N__17979));
    LocalMux I__3000 (
            .O(N__18021),
            .I(N__17976));
    LocalMux I__2999 (
            .O(N__18018),
            .I(N__17973));
    LocalMux I__2998 (
            .O(N__18015),
            .I(N__17970));
    LocalMux I__2997 (
            .O(N__18012),
            .I(N__17967));
    LocalMux I__2996 (
            .O(N__18009),
            .I(N__17960));
    Span4Mux_v I__2995 (
            .O(N__18006),
            .I(N__17960));
    LocalMux I__2994 (
            .O(N__18003),
            .I(N__17960));
    Span4Mux_v I__2993 (
            .O(N__17998),
            .I(N__17957));
    Span4Mux_v I__2992 (
            .O(N__17995),
            .I(N__17954));
    Span4Mux_h I__2991 (
            .O(N__17992),
            .I(N__17949));
    Span4Mux_v I__2990 (
            .O(N__17985),
            .I(N__17949));
    Span4Mux_h I__2989 (
            .O(N__17982),
            .I(N__17946));
    InMux I__2988 (
            .O(N__17979),
            .I(N__17943));
    Span4Mux_v I__2987 (
            .O(N__17976),
            .I(N__17940));
    Span4Mux_h I__2986 (
            .O(N__17973),
            .I(N__17935));
    Span4Mux_v I__2985 (
            .O(N__17970),
            .I(N__17935));
    Span4Mux_h I__2984 (
            .O(N__17967),
            .I(N__17930));
    Span4Mux_v I__2983 (
            .O(N__17960),
            .I(N__17930));
    Span4Mux_h I__2982 (
            .O(N__17957),
            .I(N__17927));
    Span4Mux_h I__2981 (
            .O(N__17954),
            .I(N__17924));
    Span4Mux_h I__2980 (
            .O(N__17949),
            .I(N__17921));
    Span4Mux_h I__2979 (
            .O(N__17946),
            .I(N__17918));
    LocalMux I__2978 (
            .O(N__17943),
            .I(N__17915));
    Span4Mux_h I__2977 (
            .O(N__17940),
            .I(N__17912));
    Span4Mux_h I__2976 (
            .O(N__17935),
            .I(N__17909));
    Span4Mux_h I__2975 (
            .O(N__17930),
            .I(N__17906));
    Span4Mux_h I__2974 (
            .O(N__17927),
            .I(N__17897));
    Span4Mux_h I__2973 (
            .O(N__17924),
            .I(N__17897));
    Span4Mux_h I__2972 (
            .O(N__17921),
            .I(N__17897));
    Span4Mux_v I__2971 (
            .O(N__17918),
            .I(N__17897));
    Span12Mux_s8_h I__2970 (
            .O(N__17915),
            .I(N__17894));
    Span4Mux_h I__2969 (
            .O(N__17912),
            .I(N__17887));
    Span4Mux_h I__2968 (
            .O(N__17909),
            .I(N__17887));
    Span4Mux_h I__2967 (
            .O(N__17906),
            .I(N__17887));
    Sp12to4 I__2966 (
            .O(N__17897),
            .I(N__17884));
    Odrv12 I__2965 (
            .O(N__17894),
            .I(M_this_ppu_sprites_addr_4));
    Odrv4 I__2964 (
            .O(N__17887),
            .I(M_this_ppu_sprites_addr_4));
    Odrv12 I__2963 (
            .O(N__17884),
            .I(M_this_ppu_sprites_addr_4));
    CascadeMux I__2962 (
            .O(N__17877),
            .I(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_7_cascade_ ));
    CascadeMux I__2961 (
            .O(N__17874),
            .I(N_597_cascade_));
    InMux I__2960 (
            .O(N__17871),
            .I(N__17868));
    LocalMux I__2959 (
            .O(N__17868),
            .I(M_this_sprites_address_qc_7_0));
    InMux I__2958 (
            .O(N__17865),
            .I(N__17862));
    LocalMux I__2957 (
            .O(N__17862),
            .I(N_1298_tz_0));
    InMux I__2956 (
            .O(N__17859),
            .I(N__17856));
    LocalMux I__2955 (
            .O(N__17856),
            .I(N__17853));
    Odrv4 I__2954 (
            .O(N__17853),
            .I(N_1294_tz_0));
    CascadeMux I__2953 (
            .O(N__17850),
            .I(N_602_cascade_));
    InMux I__2952 (
            .O(N__17847),
            .I(N__17844));
    LocalMux I__2951 (
            .O(N__17844),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_7 ));
    InMux I__2950 (
            .O(N__17841),
            .I(N__17838));
    LocalMux I__2949 (
            .O(N__17838),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ));
    InMux I__2948 (
            .O(N__17835),
            .I(N__17830));
    InMux I__2947 (
            .O(N__17834),
            .I(N__17827));
    InMux I__2946 (
            .O(N__17833),
            .I(N__17824));
    LocalMux I__2945 (
            .O(N__17830),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__2944 (
            .O(N__17827),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__2943 (
            .O(N__17824),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    InMux I__2942 (
            .O(N__17817),
            .I(N__17814));
    LocalMux I__2941 (
            .O(N__17814),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ));
    CascadeMux I__2940 (
            .O(N__17811),
            .I(N__17806));
    InMux I__2939 (
            .O(N__17810),
            .I(N__17803));
    InMux I__2938 (
            .O(N__17809),
            .I(N__17800));
    InMux I__2937 (
            .O(N__17806),
            .I(N__17797));
    LocalMux I__2936 (
            .O(N__17803),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__2935 (
            .O(N__17800),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__2934 (
            .O(N__17797),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    CascadeMux I__2933 (
            .O(N__17790),
            .I(N__17787));
    InMux I__2932 (
            .O(N__17787),
            .I(N__17784));
    LocalMux I__2931 (
            .O(N__17784),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ));
    CascadeMux I__2930 (
            .O(N__17781),
            .I(N__17777));
    InMux I__2929 (
            .O(N__17780),
            .I(N__17773));
    InMux I__2928 (
            .O(N__17777),
            .I(N__17770));
    InMux I__2927 (
            .O(N__17776),
            .I(N__17767));
    LocalMux I__2926 (
            .O(N__17773),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__2925 (
            .O(N__17770),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__2924 (
            .O(N__17767),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    CascadeMux I__2923 (
            .O(N__17760),
            .I(N__17753));
    CascadeMux I__2922 (
            .O(N__17759),
            .I(N__17750));
    CascadeMux I__2921 (
            .O(N__17758),
            .I(N__17745));
    InMux I__2920 (
            .O(N__17757),
            .I(N__17742));
    InMux I__2919 (
            .O(N__17756),
            .I(N__17739));
    InMux I__2918 (
            .O(N__17753),
            .I(N__17736));
    InMux I__2917 (
            .O(N__17750),
            .I(N__17733));
    CascadeMux I__2916 (
            .O(N__17749),
            .I(N__17729));
    InMux I__2915 (
            .O(N__17748),
            .I(N__17726));
    InMux I__2914 (
            .O(N__17745),
            .I(N__17723));
    LocalMux I__2913 (
            .O(N__17742),
            .I(N__17716));
    LocalMux I__2912 (
            .O(N__17739),
            .I(N__17716));
    LocalMux I__2911 (
            .O(N__17736),
            .I(N__17716));
    LocalMux I__2910 (
            .O(N__17733),
            .I(N__17713));
    InMux I__2909 (
            .O(N__17732),
            .I(N__17710));
    InMux I__2908 (
            .O(N__17729),
            .I(N__17707));
    LocalMux I__2907 (
            .O(N__17726),
            .I(N__17704));
    LocalMux I__2906 (
            .O(N__17723),
            .I(N__17697));
    Span4Mux_v I__2905 (
            .O(N__17716),
            .I(N__17697));
    Span4Mux_v I__2904 (
            .O(N__17713),
            .I(N__17697));
    LocalMux I__2903 (
            .O(N__17710),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2902 (
            .O(N__17707),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv12 I__2901 (
            .O(N__17704),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2900 (
            .O(N__17697),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    CEMux I__2899 (
            .O(N__17688),
            .I(N__17678));
    InMux I__2898 (
            .O(N__17687),
            .I(N__17664));
    InMux I__2897 (
            .O(N__17686),
            .I(N__17664));
    InMux I__2896 (
            .O(N__17685),
            .I(N__17659));
    InMux I__2895 (
            .O(N__17684),
            .I(N__17659));
    InMux I__2894 (
            .O(N__17683),
            .I(N__17654));
    InMux I__2893 (
            .O(N__17682),
            .I(N__17654));
    InMux I__2892 (
            .O(N__17681),
            .I(N__17651));
    LocalMux I__2891 (
            .O(N__17678),
            .I(N__17648));
    InMux I__2890 (
            .O(N__17677),
            .I(N__17639));
    InMux I__2889 (
            .O(N__17676),
            .I(N__17639));
    InMux I__2888 (
            .O(N__17675),
            .I(N__17639));
    InMux I__2887 (
            .O(N__17674),
            .I(N__17639));
    InMux I__2886 (
            .O(N__17673),
            .I(N__17632));
    InMux I__2885 (
            .O(N__17672),
            .I(N__17632));
    InMux I__2884 (
            .O(N__17671),
            .I(N__17632));
    InMux I__2883 (
            .O(N__17670),
            .I(N__17629));
    CEMux I__2882 (
            .O(N__17669),
            .I(N__17624));
    LocalMux I__2881 (
            .O(N__17664),
            .I(N__17621));
    LocalMux I__2880 (
            .O(N__17659),
            .I(N__17616));
    LocalMux I__2879 (
            .O(N__17654),
            .I(N__17616));
    LocalMux I__2878 (
            .O(N__17651),
            .I(N__17611));
    Span4Mux_v I__2877 (
            .O(N__17648),
            .I(N__17608));
    LocalMux I__2876 (
            .O(N__17639),
            .I(N__17601));
    LocalMux I__2875 (
            .O(N__17632),
            .I(N__17601));
    LocalMux I__2874 (
            .O(N__17629),
            .I(N__17601));
    InMux I__2873 (
            .O(N__17628),
            .I(N__17596));
    InMux I__2872 (
            .O(N__17627),
            .I(N__17596));
    LocalMux I__2871 (
            .O(N__17624),
            .I(N__17589));
    Span4Mux_h I__2870 (
            .O(N__17621),
            .I(N__17589));
    Span4Mux_v I__2869 (
            .O(N__17616),
            .I(N__17589));
    InMux I__2868 (
            .O(N__17615),
            .I(N__17586));
    InMux I__2867 (
            .O(N__17614),
            .I(N__17583));
    Span4Mux_v I__2866 (
            .O(N__17611),
            .I(N__17574));
    Span4Mux_v I__2865 (
            .O(N__17608),
            .I(N__17574));
    Span4Mux_v I__2864 (
            .O(N__17601),
            .I(N__17574));
    LocalMux I__2863 (
            .O(N__17596),
            .I(N__17574));
    Odrv4 I__2862 (
            .O(N__17589),
            .I(\this_vga_signals.GZ0Z_394 ));
    LocalMux I__2861 (
            .O(N__17586),
            .I(\this_vga_signals.GZ0Z_394 ));
    LocalMux I__2860 (
            .O(N__17583),
            .I(\this_vga_signals.GZ0Z_394 ));
    Odrv4 I__2859 (
            .O(N__17574),
            .I(\this_vga_signals.GZ0Z_394 ));
    CascadeMux I__2858 (
            .O(N__17565),
            .I(N__17562));
    InMux I__2857 (
            .O(N__17562),
            .I(N__17557));
    InMux I__2856 (
            .O(N__17561),
            .I(N__17552));
    InMux I__2855 (
            .O(N__17560),
            .I(N__17549));
    LocalMux I__2854 (
            .O(N__17557),
            .I(N__17545));
    InMux I__2853 (
            .O(N__17556),
            .I(N__17540));
    InMux I__2852 (
            .O(N__17555),
            .I(N__17540));
    LocalMux I__2851 (
            .O(N__17552),
            .I(N__17537));
    LocalMux I__2850 (
            .O(N__17549),
            .I(N__17534));
    InMux I__2849 (
            .O(N__17548),
            .I(N__17531));
    Span4Mux_v I__2848 (
            .O(N__17545),
            .I(N__17522));
    LocalMux I__2847 (
            .O(N__17540),
            .I(N__17522));
    Span4Mux_h I__2846 (
            .O(N__17537),
            .I(N__17522));
    Span4Mux_v I__2845 (
            .O(N__17534),
            .I(N__17522));
    LocalMux I__2844 (
            .O(N__17531),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv4 I__2843 (
            .O(N__17522),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    SRMux I__2842 (
            .O(N__17517),
            .I(N__17512));
    SRMux I__2841 (
            .O(N__17516),
            .I(N__17509));
    SRMux I__2840 (
            .O(N__17515),
            .I(N__17506));
    LocalMux I__2839 (
            .O(N__17512),
            .I(N__17501));
    LocalMux I__2838 (
            .O(N__17509),
            .I(N__17501));
    LocalMux I__2837 (
            .O(N__17506),
            .I(N__17498));
    Span4Mux_v I__2836 (
            .O(N__17501),
            .I(N__17494));
    Span4Mux_h I__2835 (
            .O(N__17498),
            .I(N__17491));
    InMux I__2834 (
            .O(N__17497),
            .I(N__17488));
    Span4Mux_h I__2833 (
            .O(N__17494),
            .I(N__17484));
    Span4Mux_h I__2832 (
            .O(N__17491),
            .I(N__17481));
    LocalMux I__2831 (
            .O(N__17488),
            .I(N__17478));
    InMux I__2830 (
            .O(N__17487),
            .I(N__17475));
    Odrv4 I__2829 (
            .O(N__17484),
            .I(\this_vga_signals.M_vcounter_q_501_0 ));
    Odrv4 I__2828 (
            .O(N__17481),
            .I(\this_vga_signals.M_vcounter_q_501_0 ));
    Odrv4 I__2827 (
            .O(N__17478),
            .I(\this_vga_signals.M_vcounter_q_501_0 ));
    LocalMux I__2826 (
            .O(N__17475),
            .I(\this_vga_signals.M_vcounter_q_501_0 ));
    InMux I__2825 (
            .O(N__17466),
            .I(N__17463));
    LocalMux I__2824 (
            .O(N__17463),
            .I(N__17460));
    Odrv12 I__2823 (
            .O(N__17460),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__2822 (
            .O(N__17457),
            .I(N__17454));
    LocalMux I__2821 (
            .O(N__17454),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    CEMux I__2820 (
            .O(N__17451),
            .I(N__17447));
    CEMux I__2819 (
            .O(N__17450),
            .I(N__17444));
    LocalMux I__2818 (
            .O(N__17447),
            .I(N__17439));
    LocalMux I__2817 (
            .O(N__17444),
            .I(N__17439));
    Span4Mux_v I__2816 (
            .O(N__17439),
            .I(N__17436));
    Span4Mux_h I__2815 (
            .O(N__17436),
            .I(N__17433));
    Span4Mux_h I__2814 (
            .O(N__17433),
            .I(N__17430));
    Odrv4 I__2813 (
            .O(N__17430),
            .I(\this_sprites_ram.mem_WE_10 ));
    InMux I__2812 (
            .O(N__17427),
            .I(N__17424));
    LocalMux I__2811 (
            .O(N__17424),
            .I(N__17418));
    InMux I__2810 (
            .O(N__17423),
            .I(N__17413));
    InMux I__2809 (
            .O(N__17422),
            .I(N__17413));
    InMux I__2808 (
            .O(N__17421),
            .I(N__17408));
    Span4Mux_v I__2807 (
            .O(N__17418),
            .I(N__17401));
    LocalMux I__2806 (
            .O(N__17413),
            .I(N__17401));
    InMux I__2805 (
            .O(N__17412),
            .I(N__17396));
    InMux I__2804 (
            .O(N__17411),
            .I(N__17396));
    LocalMux I__2803 (
            .O(N__17408),
            .I(N__17392));
    InMux I__2802 (
            .O(N__17407),
            .I(N__17389));
    InMux I__2801 (
            .O(N__17406),
            .I(N__17386));
    Span4Mux_h I__2800 (
            .O(N__17401),
            .I(N__17383));
    LocalMux I__2799 (
            .O(N__17396),
            .I(N__17380));
    InMux I__2798 (
            .O(N__17395),
            .I(N__17377));
    Odrv4 I__2797 (
            .O(N__17392),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2796 (
            .O(N__17389),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2795 (
            .O(N__17386),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2794 (
            .O(N__17383),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2793 (
            .O(N__17380),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2792 (
            .O(N__17377),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    CascadeMux I__2791 (
            .O(N__17364),
            .I(M_this_vga_signals_line_clk_0_cascade_));
    InMux I__2790 (
            .O(N__17361),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1 ));
    InMux I__2789 (
            .O(N__17358),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1 ));
    InMux I__2788 (
            .O(N__17355),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1 ));
    InMux I__2787 (
            .O(N__17352),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1 ));
    InMux I__2786 (
            .O(N__17349),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1 ));
    InMux I__2785 (
            .O(N__17346),
            .I(N__17343));
    LocalMux I__2784 (
            .O(N__17343),
            .I(N__17340));
    Odrv12 I__2783 (
            .O(N__17340),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ));
    InMux I__2782 (
            .O(N__17337),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1 ));
    InMux I__2781 (
            .O(N__17334),
            .I(\this_ppu.un1_M_count_q_1_cry_6_s1 ));
    InMux I__2780 (
            .O(N__17331),
            .I(N__17328));
    LocalMux I__2779 (
            .O(N__17328),
            .I(N__17319));
    CascadeMux I__2778 (
            .O(N__17327),
            .I(N__17316));
    InMux I__2777 (
            .O(N__17326),
            .I(N__17299));
    InMux I__2776 (
            .O(N__17325),
            .I(N__17294));
    InMux I__2775 (
            .O(N__17324),
            .I(N__17294));
    InMux I__2774 (
            .O(N__17323),
            .I(N__17289));
    InMux I__2773 (
            .O(N__17322),
            .I(N__17289));
    Span4Mux_v I__2772 (
            .O(N__17319),
            .I(N__17286));
    InMux I__2771 (
            .O(N__17316),
            .I(N__17283));
    InMux I__2770 (
            .O(N__17315),
            .I(N__17277));
    InMux I__2769 (
            .O(N__17314),
            .I(N__17272));
    InMux I__2768 (
            .O(N__17313),
            .I(N__17272));
    InMux I__2767 (
            .O(N__17312),
            .I(N__17265));
    InMux I__2766 (
            .O(N__17311),
            .I(N__17265));
    InMux I__2765 (
            .O(N__17310),
            .I(N__17265));
    InMux I__2764 (
            .O(N__17309),
            .I(N__17260));
    InMux I__2763 (
            .O(N__17308),
            .I(N__17260));
    InMux I__2762 (
            .O(N__17307),
            .I(N__17250));
    InMux I__2761 (
            .O(N__17306),
            .I(N__17250));
    InMux I__2760 (
            .O(N__17305),
            .I(N__17250));
    InMux I__2759 (
            .O(N__17304),
            .I(N__17250));
    InMux I__2758 (
            .O(N__17303),
            .I(N__17245));
    InMux I__2757 (
            .O(N__17302),
            .I(N__17245));
    LocalMux I__2756 (
            .O(N__17299),
            .I(N__17229));
    LocalMux I__2755 (
            .O(N__17294),
            .I(N__17229));
    LocalMux I__2754 (
            .O(N__17289),
            .I(N__17229));
    Span4Mux_h I__2753 (
            .O(N__17286),
            .I(N__17229));
    LocalMux I__2752 (
            .O(N__17283),
            .I(N__17229));
    InMux I__2751 (
            .O(N__17282),
            .I(N__17222));
    InMux I__2750 (
            .O(N__17281),
            .I(N__17222));
    InMux I__2749 (
            .O(N__17280),
            .I(N__17222));
    LocalMux I__2748 (
            .O(N__17277),
            .I(N__17219));
    LocalMux I__2747 (
            .O(N__17272),
            .I(N__17212));
    LocalMux I__2746 (
            .O(N__17265),
            .I(N__17212));
    LocalMux I__2745 (
            .O(N__17260),
            .I(N__17212));
    InMux I__2744 (
            .O(N__17259),
            .I(N__17209));
    LocalMux I__2743 (
            .O(N__17250),
            .I(N__17206));
    LocalMux I__2742 (
            .O(N__17245),
            .I(N__17203));
    InMux I__2741 (
            .O(N__17244),
            .I(N__17192));
    InMux I__2740 (
            .O(N__17243),
            .I(N__17192));
    InMux I__2739 (
            .O(N__17242),
            .I(N__17192));
    InMux I__2738 (
            .O(N__17241),
            .I(N__17192));
    InMux I__2737 (
            .O(N__17240),
            .I(N__17192));
    Span4Mux_v I__2736 (
            .O(N__17229),
            .I(N__17189));
    LocalMux I__2735 (
            .O(N__17222),
            .I(N__17186));
    Span4Mux_v I__2734 (
            .O(N__17219),
            .I(N__17181));
    Span4Mux_v I__2733 (
            .O(N__17212),
            .I(N__17181));
    LocalMux I__2732 (
            .O(N__17209),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__2731 (
            .O(N__17206),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__2730 (
            .O(N__17203),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__2729 (
            .O(N__17192),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__2728 (
            .O(N__17189),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__2727 (
            .O(N__17186),
            .I(\this_vga_signals.vaddress_5 ));
    Odrv4 I__2726 (
            .O(N__17181),
            .I(\this_vga_signals.vaddress_5 ));
    InMux I__2725 (
            .O(N__17166),
            .I(N__17157));
    InMux I__2724 (
            .O(N__17165),
            .I(N__17154));
    InMux I__2723 (
            .O(N__17164),
            .I(N__17144));
    InMux I__2722 (
            .O(N__17163),
            .I(N__17144));
    InMux I__2721 (
            .O(N__17162),
            .I(N__17144));
    InMux I__2720 (
            .O(N__17161),
            .I(N__17144));
    InMux I__2719 (
            .O(N__17160),
            .I(N__17135));
    LocalMux I__2718 (
            .O(N__17157),
            .I(N__17130));
    LocalMux I__2717 (
            .O(N__17154),
            .I(N__17130));
    InMux I__2716 (
            .O(N__17153),
            .I(N__17127));
    LocalMux I__2715 (
            .O(N__17144),
            .I(N__17124));
    InMux I__2714 (
            .O(N__17143),
            .I(N__17119));
    InMux I__2713 (
            .O(N__17142),
            .I(N__17119));
    CascadeMux I__2712 (
            .O(N__17141),
            .I(N__17115));
    InMux I__2711 (
            .O(N__17140),
            .I(N__17109));
    InMux I__2710 (
            .O(N__17139),
            .I(N__17109));
    InMux I__2709 (
            .O(N__17138),
            .I(N__17106));
    LocalMux I__2708 (
            .O(N__17135),
            .I(N__17101));
    Span4Mux_v I__2707 (
            .O(N__17130),
            .I(N__17101));
    LocalMux I__2706 (
            .O(N__17127),
            .I(N__17094));
    Span4Mux_v I__2705 (
            .O(N__17124),
            .I(N__17094));
    LocalMux I__2704 (
            .O(N__17119),
            .I(N__17094));
    InMux I__2703 (
            .O(N__17118),
            .I(N__17091));
    InMux I__2702 (
            .O(N__17115),
            .I(N__17086));
    InMux I__2701 (
            .O(N__17114),
            .I(N__17086));
    LocalMux I__2700 (
            .O(N__17109),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2699 (
            .O(N__17106),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__2698 (
            .O(N__17101),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__2697 (
            .O(N__17094),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2696 (
            .O(N__17091),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2695 (
            .O(N__17086),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__2694 (
            .O(N__17073),
            .I(N__17070));
    InMux I__2693 (
            .O(N__17070),
            .I(N__17067));
    LocalMux I__2692 (
            .O(N__17067),
            .I(\this_vga_signals.vaddress_0_0_6 ));
    InMux I__2691 (
            .O(N__17064),
            .I(N__17059));
    InMux I__2690 (
            .O(N__17063),
            .I(N__17053));
    InMux I__2689 (
            .O(N__17062),
            .I(N__17053));
    LocalMux I__2688 (
            .O(N__17059),
            .I(N__17050));
    InMux I__2687 (
            .O(N__17058),
            .I(N__17046));
    LocalMux I__2686 (
            .O(N__17053),
            .I(N__17042));
    Span4Mux_h I__2685 (
            .O(N__17050),
            .I(N__17039));
    InMux I__2684 (
            .O(N__17049),
            .I(N__17036));
    LocalMux I__2683 (
            .O(N__17046),
            .I(N__17033));
    InMux I__2682 (
            .O(N__17045),
            .I(N__17030));
    Span4Mux_v I__2681 (
            .O(N__17042),
            .I(N__17023));
    Span4Mux_h I__2680 (
            .O(N__17039),
            .I(N__17020));
    LocalMux I__2679 (
            .O(N__17036),
            .I(N__17017));
    Span4Mux_v I__2678 (
            .O(N__17033),
            .I(N__17012));
    LocalMux I__2677 (
            .O(N__17030),
            .I(N__17012));
    InMux I__2676 (
            .O(N__17029),
            .I(N__17009));
    InMux I__2675 (
            .O(N__17028),
            .I(N__17004));
    InMux I__2674 (
            .O(N__17027),
            .I(N__17004));
    InMux I__2673 (
            .O(N__17026),
            .I(N__17001));
    Odrv4 I__2672 (
            .O(N__17023),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__2671 (
            .O(N__17020),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__2670 (
            .O(N__17017),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__2669 (
            .O(N__17012),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__2668 (
            .O(N__17009),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__2667 (
            .O(N__17004),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__2666 (
            .O(N__17001),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    InMux I__2665 (
            .O(N__16986),
            .I(N__16977));
    InMux I__2664 (
            .O(N__16985),
            .I(N__16974));
    CascadeMux I__2663 (
            .O(N__16984),
            .I(N__16966));
    CascadeMux I__2662 (
            .O(N__16983),
            .I(N__16963));
    CascadeMux I__2661 (
            .O(N__16982),
            .I(N__16958));
    CascadeMux I__2660 (
            .O(N__16981),
            .I(N__16954));
    CascadeMux I__2659 (
            .O(N__16980),
            .I(N__16949));
    LocalMux I__2658 (
            .O(N__16977),
            .I(N__16942));
    LocalMux I__2657 (
            .O(N__16974),
            .I(N__16942));
    InMux I__2656 (
            .O(N__16973),
            .I(N__16939));
    InMux I__2655 (
            .O(N__16972),
            .I(N__16936));
    InMux I__2654 (
            .O(N__16971),
            .I(N__16933));
    InMux I__2653 (
            .O(N__16970),
            .I(N__16924));
    InMux I__2652 (
            .O(N__16969),
            .I(N__16924));
    InMux I__2651 (
            .O(N__16966),
            .I(N__16924));
    InMux I__2650 (
            .O(N__16963),
            .I(N__16919));
    InMux I__2649 (
            .O(N__16962),
            .I(N__16919));
    InMux I__2648 (
            .O(N__16961),
            .I(N__16914));
    InMux I__2647 (
            .O(N__16958),
            .I(N__16914));
    InMux I__2646 (
            .O(N__16957),
            .I(N__16911));
    InMux I__2645 (
            .O(N__16954),
            .I(N__16903));
    InMux I__2644 (
            .O(N__16953),
            .I(N__16903));
    InMux I__2643 (
            .O(N__16952),
            .I(N__16898));
    InMux I__2642 (
            .O(N__16949),
            .I(N__16898));
    InMux I__2641 (
            .O(N__16948),
            .I(N__16895));
    InMux I__2640 (
            .O(N__16947),
            .I(N__16892));
    Span4Mux_v I__2639 (
            .O(N__16942),
            .I(N__16889));
    LocalMux I__2638 (
            .O(N__16939),
            .I(N__16882));
    LocalMux I__2637 (
            .O(N__16936),
            .I(N__16882));
    LocalMux I__2636 (
            .O(N__16933),
            .I(N__16882));
    InMux I__2635 (
            .O(N__16932),
            .I(N__16879));
    InMux I__2634 (
            .O(N__16931),
            .I(N__16876));
    LocalMux I__2633 (
            .O(N__16924),
            .I(N__16871));
    LocalMux I__2632 (
            .O(N__16919),
            .I(N__16871));
    LocalMux I__2631 (
            .O(N__16914),
            .I(N__16866));
    LocalMux I__2630 (
            .O(N__16911),
            .I(N__16866));
    InMux I__2629 (
            .O(N__16910),
            .I(N__16863));
    InMux I__2628 (
            .O(N__16909),
            .I(N__16860));
    InMux I__2627 (
            .O(N__16908),
            .I(N__16857));
    LocalMux I__2626 (
            .O(N__16903),
            .I(N__16848));
    LocalMux I__2625 (
            .O(N__16898),
            .I(N__16848));
    LocalMux I__2624 (
            .O(N__16895),
            .I(N__16848));
    LocalMux I__2623 (
            .O(N__16892),
            .I(N__16848));
    Span4Mux_h I__2622 (
            .O(N__16889),
            .I(N__16843));
    Span4Mux_v I__2621 (
            .O(N__16882),
            .I(N__16843));
    LocalMux I__2620 (
            .O(N__16879),
            .I(N__16832));
    LocalMux I__2619 (
            .O(N__16876),
            .I(N__16832));
    Span4Mux_v I__2618 (
            .O(N__16871),
            .I(N__16832));
    Span4Mux_h I__2617 (
            .O(N__16866),
            .I(N__16832));
    LocalMux I__2616 (
            .O(N__16863),
            .I(N__16832));
    LocalMux I__2615 (
            .O(N__16860),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2614 (
            .O(N__16857),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv12 I__2613 (
            .O(N__16848),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2612 (
            .O(N__16843),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2611 (
            .O(N__16832),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    CascadeMux I__2610 (
            .O(N__16821),
            .I(N__16815));
    CascadeMux I__2609 (
            .O(N__16820),
            .I(N__16812));
    CascadeMux I__2608 (
            .O(N__16819),
            .I(N__16806));
    InMux I__2607 (
            .O(N__16818),
            .I(N__16799));
    InMux I__2606 (
            .O(N__16815),
            .I(N__16799));
    InMux I__2605 (
            .O(N__16812),
            .I(N__16799));
    CascadeMux I__2604 (
            .O(N__16811),
            .I(N__16796));
    CascadeMux I__2603 (
            .O(N__16810),
            .I(N__16785));
    CascadeMux I__2602 (
            .O(N__16809),
            .I(N__16780));
    InMux I__2601 (
            .O(N__16806),
            .I(N__16775));
    LocalMux I__2600 (
            .O(N__16799),
            .I(N__16772));
    InMux I__2599 (
            .O(N__16796),
            .I(N__16767));
    InMux I__2598 (
            .O(N__16795),
            .I(N__16767));
    InMux I__2597 (
            .O(N__16794),
            .I(N__16761));
    CascadeMux I__2596 (
            .O(N__16793),
            .I(N__16758));
    CascadeMux I__2595 (
            .O(N__16792),
            .I(N__16751));
    InMux I__2594 (
            .O(N__16791),
            .I(N__16747));
    InMux I__2593 (
            .O(N__16790),
            .I(N__16744));
    InMux I__2592 (
            .O(N__16789),
            .I(N__16741));
    InMux I__2591 (
            .O(N__16788),
            .I(N__16738));
    InMux I__2590 (
            .O(N__16785),
            .I(N__16733));
    InMux I__2589 (
            .O(N__16784),
            .I(N__16733));
    InMux I__2588 (
            .O(N__16783),
            .I(N__16729));
    InMux I__2587 (
            .O(N__16780),
            .I(N__16722));
    InMux I__2586 (
            .O(N__16779),
            .I(N__16722));
    InMux I__2585 (
            .O(N__16778),
            .I(N__16722));
    LocalMux I__2584 (
            .O(N__16775),
            .I(N__16711));
    Span4Mux_h I__2583 (
            .O(N__16772),
            .I(N__16711));
    LocalMux I__2582 (
            .O(N__16767),
            .I(N__16711));
    InMux I__2581 (
            .O(N__16766),
            .I(N__16708));
    InMux I__2580 (
            .O(N__16765),
            .I(N__16703));
    InMux I__2579 (
            .O(N__16764),
            .I(N__16703));
    LocalMux I__2578 (
            .O(N__16761),
            .I(N__16700));
    InMux I__2577 (
            .O(N__16758),
            .I(N__16697));
    InMux I__2576 (
            .O(N__16757),
            .I(N__16690));
    InMux I__2575 (
            .O(N__16756),
            .I(N__16690));
    InMux I__2574 (
            .O(N__16755),
            .I(N__16690));
    InMux I__2573 (
            .O(N__16754),
            .I(N__16683));
    InMux I__2572 (
            .O(N__16751),
            .I(N__16683));
    InMux I__2571 (
            .O(N__16750),
            .I(N__16683));
    LocalMux I__2570 (
            .O(N__16747),
            .I(N__16676));
    LocalMux I__2569 (
            .O(N__16744),
            .I(N__16676));
    LocalMux I__2568 (
            .O(N__16741),
            .I(N__16676));
    LocalMux I__2567 (
            .O(N__16738),
            .I(N__16671));
    LocalMux I__2566 (
            .O(N__16733),
            .I(N__16671));
    InMux I__2565 (
            .O(N__16732),
            .I(N__16668));
    LocalMux I__2564 (
            .O(N__16729),
            .I(N__16665));
    LocalMux I__2563 (
            .O(N__16722),
            .I(N__16662));
    InMux I__2562 (
            .O(N__16721),
            .I(N__16655));
    InMux I__2561 (
            .O(N__16720),
            .I(N__16655));
    InMux I__2560 (
            .O(N__16719),
            .I(N__16655));
    InMux I__2559 (
            .O(N__16718),
            .I(N__16652));
    Span4Mux_v I__2558 (
            .O(N__16711),
            .I(N__16649));
    LocalMux I__2557 (
            .O(N__16708),
            .I(N__16640));
    LocalMux I__2556 (
            .O(N__16703),
            .I(N__16640));
    Span4Mux_v I__2555 (
            .O(N__16700),
            .I(N__16640));
    LocalMux I__2554 (
            .O(N__16697),
            .I(N__16640));
    LocalMux I__2553 (
            .O(N__16690),
            .I(N__16635));
    LocalMux I__2552 (
            .O(N__16683),
            .I(N__16635));
    Span4Mux_v I__2551 (
            .O(N__16676),
            .I(N__16632));
    Span4Mux_v I__2550 (
            .O(N__16671),
            .I(N__16629));
    LocalMux I__2549 (
            .O(N__16668),
            .I(N__16626));
    Span4Mux_h I__2548 (
            .O(N__16665),
            .I(N__16619));
    Span4Mux_h I__2547 (
            .O(N__16662),
            .I(N__16619));
    LocalMux I__2546 (
            .O(N__16655),
            .I(N__16619));
    LocalMux I__2545 (
            .O(N__16652),
            .I(N__16608));
    Span4Mux_h I__2544 (
            .O(N__16649),
            .I(N__16608));
    Span4Mux_v I__2543 (
            .O(N__16640),
            .I(N__16608));
    Span4Mux_v I__2542 (
            .O(N__16635),
            .I(N__16608));
    Span4Mux_h I__2541 (
            .O(N__16632),
            .I(N__16608));
    Odrv4 I__2540 (
            .O(N__16629),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__2539 (
            .O(N__16626),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2538 (
            .O(N__16619),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2537 (
            .O(N__16608),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    CascadeMux I__2536 (
            .O(N__16599),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_1_cascade_ ));
    CascadeMux I__2535 (
            .O(N__16596),
            .I(N__16593));
    InMux I__2534 (
            .O(N__16593),
            .I(N__16586));
    CascadeMux I__2533 (
            .O(N__16592),
            .I(N__16583));
    CascadeMux I__2532 (
            .O(N__16591),
            .I(N__16579));
    InMux I__2531 (
            .O(N__16590),
            .I(N__16576));
    InMux I__2530 (
            .O(N__16589),
            .I(N__16573));
    LocalMux I__2529 (
            .O(N__16586),
            .I(N__16570));
    InMux I__2528 (
            .O(N__16583),
            .I(N__16563));
    InMux I__2527 (
            .O(N__16582),
            .I(N__16563));
    InMux I__2526 (
            .O(N__16579),
            .I(N__16563));
    LocalMux I__2525 (
            .O(N__16576),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__2524 (
            .O(N__16573),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    Odrv4 I__2523 (
            .O(N__16570),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    LocalMux I__2522 (
            .O(N__16563),
            .I(\this_vga_signals.mult1_un54_sum_c3_1 ));
    InMux I__2521 (
            .O(N__16554),
            .I(N__16551));
    LocalMux I__2520 (
            .O(N__16551),
            .I(N__16548));
    Span4Mux_h I__2519 (
            .O(N__16548),
            .I(N__16545));
    Odrv4 I__2518 (
            .O(N__16545),
            .I(\this_vga_signals.g0_0_0 ));
    CascadeMux I__2517 (
            .O(N__16542),
            .I(\this_ppu.un13_0_cascade_ ));
    CascadeMux I__2516 (
            .O(N__16539),
            .I(\this_ppu.M_line_clk_out_0_cascade_ ));
    InMux I__2515 (
            .O(N__16536),
            .I(N__16532));
    InMux I__2514 (
            .O(N__16535),
            .I(N__16529));
    LocalMux I__2513 (
            .O(N__16532),
            .I(N__16525));
    LocalMux I__2512 (
            .O(N__16529),
            .I(N__16522));
    InMux I__2511 (
            .O(N__16528),
            .I(N__16519));
    Span4Mux_v I__2510 (
            .O(N__16525),
            .I(N__16516));
    Span4Mux_h I__2509 (
            .O(N__16522),
            .I(N__16513));
    LocalMux I__2508 (
            .O(N__16519),
            .I(\this_vga_signals.M_vcounter_d7lt9_1 ));
    Odrv4 I__2507 (
            .O(N__16516),
            .I(\this_vga_signals.M_vcounter_d7lt9_1 ));
    Odrv4 I__2506 (
            .O(N__16513),
            .I(\this_vga_signals.M_vcounter_d7lt9_1 ));
    CascadeMux I__2505 (
            .O(N__16506),
            .I(N__16502));
    CascadeMux I__2504 (
            .O(N__16505),
            .I(N__16496));
    InMux I__2503 (
            .O(N__16502),
            .I(N__16491));
    InMux I__2502 (
            .O(N__16501),
            .I(N__16488));
    InMux I__2501 (
            .O(N__16500),
            .I(N__16485));
    InMux I__2500 (
            .O(N__16499),
            .I(N__16482));
    InMux I__2499 (
            .O(N__16496),
            .I(N__16479));
    InMux I__2498 (
            .O(N__16495),
            .I(N__16473));
    CascadeMux I__2497 (
            .O(N__16494),
            .I(N__16469));
    LocalMux I__2496 (
            .O(N__16491),
            .I(N__16461));
    LocalMux I__2495 (
            .O(N__16488),
            .I(N__16461));
    LocalMux I__2494 (
            .O(N__16485),
            .I(N__16456));
    LocalMux I__2493 (
            .O(N__16482),
            .I(N__16456));
    LocalMux I__2492 (
            .O(N__16479),
            .I(N__16453));
    InMux I__2491 (
            .O(N__16478),
            .I(N__16448));
    InMux I__2490 (
            .O(N__16477),
            .I(N__16448));
    CascadeMux I__2489 (
            .O(N__16476),
            .I(N__16443));
    LocalMux I__2488 (
            .O(N__16473),
            .I(N__16440));
    CascadeMux I__2487 (
            .O(N__16472),
            .I(N__16437));
    InMux I__2486 (
            .O(N__16469),
            .I(N__16432));
    InMux I__2485 (
            .O(N__16468),
            .I(N__16432));
    InMux I__2484 (
            .O(N__16467),
            .I(N__16427));
    InMux I__2483 (
            .O(N__16466),
            .I(N__16427));
    Span4Mux_v I__2482 (
            .O(N__16461),
            .I(N__16418));
    Span4Mux_v I__2481 (
            .O(N__16456),
            .I(N__16418));
    Span4Mux_h I__2480 (
            .O(N__16453),
            .I(N__16418));
    LocalMux I__2479 (
            .O(N__16448),
            .I(N__16418));
    InMux I__2478 (
            .O(N__16447),
            .I(N__16411));
    InMux I__2477 (
            .O(N__16446),
            .I(N__16411));
    InMux I__2476 (
            .O(N__16443),
            .I(N__16411));
    Span4Mux_v I__2475 (
            .O(N__16440),
            .I(N__16407));
    InMux I__2474 (
            .O(N__16437),
            .I(N__16404));
    LocalMux I__2473 (
            .O(N__16432),
            .I(N__16401));
    LocalMux I__2472 (
            .O(N__16427),
            .I(N__16396));
    Span4Mux_h I__2471 (
            .O(N__16418),
            .I(N__16396));
    LocalMux I__2470 (
            .O(N__16411),
            .I(N__16393));
    InMux I__2469 (
            .O(N__16410),
            .I(N__16390));
    Odrv4 I__2468 (
            .O(N__16407),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2467 (
            .O(N__16404),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2466 (
            .O(N__16401),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2465 (
            .O(N__16396),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv12 I__2464 (
            .O(N__16393),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2463 (
            .O(N__16390),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    CascadeMux I__2462 (
            .O(N__16377),
            .I(N__16372));
    CascadeMux I__2461 (
            .O(N__16376),
            .I(N__16369));
    InMux I__2460 (
            .O(N__16375),
            .I(N__16357));
    InMux I__2459 (
            .O(N__16372),
            .I(N__16354));
    InMux I__2458 (
            .O(N__16369),
            .I(N__16351));
    InMux I__2457 (
            .O(N__16368),
            .I(N__16347));
    InMux I__2456 (
            .O(N__16367),
            .I(N__16344));
    InMux I__2455 (
            .O(N__16366),
            .I(N__16339));
    InMux I__2454 (
            .O(N__16365),
            .I(N__16339));
    InMux I__2453 (
            .O(N__16364),
            .I(N__16336));
    InMux I__2452 (
            .O(N__16363),
            .I(N__16332));
    InMux I__2451 (
            .O(N__16362),
            .I(N__16327));
    InMux I__2450 (
            .O(N__16361),
            .I(N__16327));
    InMux I__2449 (
            .O(N__16360),
            .I(N__16324));
    LocalMux I__2448 (
            .O(N__16357),
            .I(N__16321));
    LocalMux I__2447 (
            .O(N__16354),
            .I(N__16318));
    LocalMux I__2446 (
            .O(N__16351),
            .I(N__16315));
    InMux I__2445 (
            .O(N__16350),
            .I(N__16312));
    LocalMux I__2444 (
            .O(N__16347),
            .I(N__16303));
    LocalMux I__2443 (
            .O(N__16344),
            .I(N__16303));
    LocalMux I__2442 (
            .O(N__16339),
            .I(N__16303));
    LocalMux I__2441 (
            .O(N__16336),
            .I(N__16303));
    CascadeMux I__2440 (
            .O(N__16335),
            .I(N__16298));
    LocalMux I__2439 (
            .O(N__16332),
            .I(N__16291));
    LocalMux I__2438 (
            .O(N__16327),
            .I(N__16291));
    LocalMux I__2437 (
            .O(N__16324),
            .I(N__16291));
    Span4Mux_v I__2436 (
            .O(N__16321),
            .I(N__16284));
    Span4Mux_h I__2435 (
            .O(N__16318),
            .I(N__16284));
    Span4Mux_v I__2434 (
            .O(N__16315),
            .I(N__16284));
    LocalMux I__2433 (
            .O(N__16312),
            .I(N__16279));
    Span4Mux_v I__2432 (
            .O(N__16303),
            .I(N__16279));
    InMux I__2431 (
            .O(N__16302),
            .I(N__16274));
    InMux I__2430 (
            .O(N__16301),
            .I(N__16274));
    InMux I__2429 (
            .O(N__16298),
            .I(N__16271));
    Odrv4 I__2428 (
            .O(N__16291),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2427 (
            .O(N__16284),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2426 (
            .O(N__16279),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2425 (
            .O(N__16274),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2424 (
            .O(N__16271),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    CascadeMux I__2423 (
            .O(N__16260),
            .I(N__16257));
    InMux I__2422 (
            .O(N__16257),
            .I(N__16254));
    LocalMux I__2421 (
            .O(N__16254),
            .I(\this_vga_signals.un4_lvisibility_1 ));
    InMux I__2420 (
            .O(N__16251),
            .I(N__16245));
    InMux I__2419 (
            .O(N__16250),
            .I(N__16245));
    LocalMux I__2418 (
            .O(N__16245),
            .I(N__16242));
    Span4Mux_h I__2417 (
            .O(N__16242),
            .I(N__16239));
    Odrv4 I__2416 (
            .O(N__16239),
            .I(\this_vga_signals.line_clk_1 ));
    InMux I__2415 (
            .O(N__16236),
            .I(N__16230));
    InMux I__2414 (
            .O(N__16235),
            .I(N__16225));
    InMux I__2413 (
            .O(N__16234),
            .I(N__16225));
    InMux I__2412 (
            .O(N__16233),
            .I(N__16219));
    LocalMux I__2411 (
            .O(N__16230),
            .I(N__16214));
    LocalMux I__2410 (
            .O(N__16225),
            .I(N__16211));
    InMux I__2409 (
            .O(N__16224),
            .I(N__16206));
    InMux I__2408 (
            .O(N__16223),
            .I(N__16206));
    CascadeMux I__2407 (
            .O(N__16222),
            .I(N__16203));
    LocalMux I__2406 (
            .O(N__16219),
            .I(N__16200));
    InMux I__2405 (
            .O(N__16218),
            .I(N__16197));
    InMux I__2404 (
            .O(N__16217),
            .I(N__16194));
    Span4Mux_v I__2403 (
            .O(N__16214),
            .I(N__16189));
    Span4Mux_v I__2402 (
            .O(N__16211),
            .I(N__16189));
    LocalMux I__2401 (
            .O(N__16206),
            .I(N__16186));
    InMux I__2400 (
            .O(N__16203),
            .I(N__16183));
    Odrv4 I__2399 (
            .O(N__16200),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2398 (
            .O(N__16197),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2397 (
            .O(N__16194),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2396 (
            .O(N__16189),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2395 (
            .O(N__16186),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2394 (
            .O(N__16183),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    CascadeMux I__2393 (
            .O(N__16170),
            .I(\this_vga_signals.un4_lvisibility_1_cascade_ ));
    InMux I__2392 (
            .O(N__16167),
            .I(N__16162));
    InMux I__2391 (
            .O(N__16166),
            .I(N__16158));
    InMux I__2390 (
            .O(N__16165),
            .I(N__16155));
    LocalMux I__2389 (
            .O(N__16162),
            .I(N__16152));
    InMux I__2388 (
            .O(N__16161),
            .I(N__16149));
    LocalMux I__2387 (
            .O(N__16158),
            .I(N__16143));
    LocalMux I__2386 (
            .O(N__16155),
            .I(N__16143));
    Span4Mux_v I__2385 (
            .O(N__16152),
            .I(N__16138));
    LocalMux I__2384 (
            .O(N__16149),
            .I(N__16138));
    InMux I__2383 (
            .O(N__16148),
            .I(N__16135));
    Span4Mux_h I__2382 (
            .O(N__16143),
            .I(N__16132));
    Odrv4 I__2381 (
            .O(N__16138),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__2380 (
            .O(N__16135),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    Odrv4 I__2379 (
            .O(N__16132),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    InMux I__2378 (
            .O(N__16125),
            .I(N__16116));
    InMux I__2377 (
            .O(N__16124),
            .I(N__16116));
    InMux I__2376 (
            .O(N__16123),
            .I(N__16111));
    InMux I__2375 (
            .O(N__16122),
            .I(N__16104));
    InMux I__2374 (
            .O(N__16121),
            .I(N__16101));
    LocalMux I__2373 (
            .O(N__16116),
            .I(N__16098));
    InMux I__2372 (
            .O(N__16115),
            .I(N__16095));
    InMux I__2371 (
            .O(N__16114),
            .I(N__16088));
    LocalMux I__2370 (
            .O(N__16111),
            .I(N__16085));
    InMux I__2369 (
            .O(N__16110),
            .I(N__16080));
    InMux I__2368 (
            .O(N__16109),
            .I(N__16080));
    InMux I__2367 (
            .O(N__16108),
            .I(N__16075));
    InMux I__2366 (
            .O(N__16107),
            .I(N__16075));
    LocalMux I__2365 (
            .O(N__16104),
            .I(N__16068));
    LocalMux I__2364 (
            .O(N__16101),
            .I(N__16068));
    Span4Mux_h I__2363 (
            .O(N__16098),
            .I(N__16068));
    LocalMux I__2362 (
            .O(N__16095),
            .I(N__16065));
    InMux I__2361 (
            .O(N__16094),
            .I(N__16060));
    InMux I__2360 (
            .O(N__16093),
            .I(N__16060));
    InMux I__2359 (
            .O(N__16092),
            .I(N__16055));
    InMux I__2358 (
            .O(N__16091),
            .I(N__16055));
    LocalMux I__2357 (
            .O(N__16088),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    Odrv4 I__2356 (
            .O(N__16085),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__2355 (
            .O(N__16080),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__2354 (
            .O(N__16075),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    Odrv4 I__2353 (
            .O(N__16068),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    Odrv4 I__2352 (
            .O(N__16065),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__2351 (
            .O(N__16060),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__2350 (
            .O(N__16055),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    CascadeMux I__2349 (
            .O(N__16038),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_cascade_ ));
    InMux I__2348 (
            .O(N__16035),
            .I(N__16032));
    LocalMux I__2347 (
            .O(N__16032),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ));
    InMux I__2346 (
            .O(N__16029),
            .I(N__16023));
    InMux I__2345 (
            .O(N__16028),
            .I(N__16018));
    InMux I__2344 (
            .O(N__16027),
            .I(N__16018));
    InMux I__2343 (
            .O(N__16026),
            .I(N__16015));
    LocalMux I__2342 (
            .O(N__16023),
            .I(N__16012));
    LocalMux I__2341 (
            .O(N__16018),
            .I(N__16009));
    LocalMux I__2340 (
            .O(N__16015),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    Odrv4 I__2339 (
            .O(N__16012),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    Odrv12 I__2338 (
            .O(N__16009),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    CascadeMux I__2337 (
            .O(N__16002),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_cascade_ ));
    InMux I__2336 (
            .O(N__15999),
            .I(N__15996));
    LocalMux I__2335 (
            .O(N__15996),
            .I(N__15989));
    InMux I__2334 (
            .O(N__15995),
            .I(N__15978));
    InMux I__2333 (
            .O(N__15994),
            .I(N__15978));
    InMux I__2332 (
            .O(N__15993),
            .I(N__15978));
    InMux I__2331 (
            .O(N__15992),
            .I(N__15975));
    Span4Mux_h I__2330 (
            .O(N__15989),
            .I(N__15972));
    InMux I__2329 (
            .O(N__15988),
            .I(N__15969));
    InMux I__2328 (
            .O(N__15987),
            .I(N__15962));
    InMux I__2327 (
            .O(N__15986),
            .I(N__15962));
    InMux I__2326 (
            .O(N__15985),
            .I(N__15962));
    LocalMux I__2325 (
            .O(N__15978),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_ns ));
    LocalMux I__2324 (
            .O(N__15975),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_ns ));
    Odrv4 I__2323 (
            .O(N__15972),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_ns ));
    LocalMux I__2322 (
            .O(N__15969),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_ns ));
    LocalMux I__2321 (
            .O(N__15962),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_ns ));
    InMux I__2320 (
            .O(N__15951),
            .I(N__15948));
    LocalMux I__2319 (
            .O(N__15948),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ));
    CascadeMux I__2318 (
            .O(N__15945),
            .I(N__15942));
    InMux I__2317 (
            .O(N__15942),
            .I(N__15939));
    LocalMux I__2316 (
            .O(N__15939),
            .I(N__15936));
    Odrv4 I__2315 (
            .O(N__15936),
            .I(\this_vga_signals.g0_i_i_a5_1_0_0_0 ));
    InMux I__2314 (
            .O(N__15933),
            .I(N__15930));
    LocalMux I__2313 (
            .O(N__15930),
            .I(\this_vga_signals.g0_i_i_0_0_0 ));
    CascadeMux I__2312 (
            .O(N__15927),
            .I(\this_vga_signals.vaddress_2_6_cascade_ ));
    InMux I__2311 (
            .O(N__15924),
            .I(N__15921));
    LocalMux I__2310 (
            .O(N__15921),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_0 ));
    CascadeMux I__2309 (
            .O(N__15918),
            .I(N__15915));
    InMux I__2308 (
            .O(N__15915),
            .I(N__15912));
    LocalMux I__2307 (
            .O(N__15912),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_0 ));
    InMux I__2306 (
            .O(N__15909),
            .I(N__15903));
    CascadeMux I__2305 (
            .O(N__15908),
            .I(N__15900));
    CascadeMux I__2304 (
            .O(N__15907),
            .I(N__15896));
    InMux I__2303 (
            .O(N__15906),
            .I(N__15893));
    LocalMux I__2302 (
            .O(N__15903),
            .I(N__15890));
    InMux I__2301 (
            .O(N__15900),
            .I(N__15887));
    InMux I__2300 (
            .O(N__15899),
            .I(N__15882));
    InMux I__2299 (
            .O(N__15896),
            .I(N__15882));
    LocalMux I__2298 (
            .O(N__15893),
            .I(N__15877));
    Span4Mux_v I__2297 (
            .O(N__15890),
            .I(N__15877));
    LocalMux I__2296 (
            .O(N__15887),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__2295 (
            .O(N__15882),
            .I(\this_vga_signals.vaddress_6 ));
    Odrv4 I__2294 (
            .O(N__15877),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__2293 (
            .O(N__15870),
            .I(N__15867));
    LocalMux I__2292 (
            .O(N__15867),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    InMux I__2291 (
            .O(N__15864),
            .I(N__15861));
    LocalMux I__2290 (
            .O(N__15861),
            .I(N__15856));
    InMux I__2289 (
            .O(N__15860),
            .I(N__15851));
    InMux I__2288 (
            .O(N__15859),
            .I(N__15851));
    Odrv12 I__2287 (
            .O(N__15856),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_0_0 ));
    LocalMux I__2286 (
            .O(N__15851),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_0_0 ));
    InMux I__2285 (
            .O(N__15846),
            .I(N__15843));
    LocalMux I__2284 (
            .O(N__15843),
            .I(N__15840));
    Span4Mux_v I__2283 (
            .O(N__15840),
            .I(N__15837));
    Odrv4 I__2282 (
            .O(N__15837),
            .I(\this_vga_signals.N_7_1_0 ));
    InMux I__2281 (
            .O(N__15834),
            .I(bfn_15_21_0_));
    InMux I__2280 (
            .O(N__15831),
            .I(N__15828));
    LocalMux I__2279 (
            .O(N__15828),
            .I(N__15822));
    InMux I__2278 (
            .O(N__15827),
            .I(N__15819));
    InMux I__2277 (
            .O(N__15826),
            .I(N__15815));
    InMux I__2276 (
            .O(N__15825),
            .I(N__15811));
    Span4Mux_v I__2275 (
            .O(N__15822),
            .I(N__15805));
    LocalMux I__2274 (
            .O(N__15819),
            .I(N__15805));
    InMux I__2273 (
            .O(N__15818),
            .I(N__15802));
    LocalMux I__2272 (
            .O(N__15815),
            .I(N__15799));
    CascadeMux I__2271 (
            .O(N__15814),
            .I(N__15795));
    LocalMux I__2270 (
            .O(N__15811),
            .I(N__15791));
    InMux I__2269 (
            .O(N__15810),
            .I(N__15788));
    Span4Mux_h I__2268 (
            .O(N__15805),
            .I(N__15785));
    LocalMux I__2267 (
            .O(N__15802),
            .I(N__15780));
    Span4Mux_h I__2266 (
            .O(N__15799),
            .I(N__15780));
    InMux I__2265 (
            .O(N__15798),
            .I(N__15775));
    InMux I__2264 (
            .O(N__15795),
            .I(N__15775));
    InMux I__2263 (
            .O(N__15794),
            .I(N__15772));
    Odrv12 I__2262 (
            .O(N__15791),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2261 (
            .O(N__15788),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__2260 (
            .O(N__15785),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__2259 (
            .O(N__15780),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2258 (
            .O(N__15775),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2257 (
            .O(N__15772),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    CEMux I__2256 (
            .O(N__15759),
            .I(N__15756));
    LocalMux I__2255 (
            .O(N__15756),
            .I(\this_vga_signals.N_966_1 ));
    CEMux I__2254 (
            .O(N__15753),
            .I(N__15749));
    CEMux I__2253 (
            .O(N__15752),
            .I(N__15746));
    LocalMux I__2252 (
            .O(N__15749),
            .I(N__15743));
    LocalMux I__2251 (
            .O(N__15746),
            .I(N__15740));
    Span4Mux_h I__2250 (
            .O(N__15743),
            .I(N__15737));
    Span4Mux_v I__2249 (
            .O(N__15740),
            .I(N__15734));
    Span4Mux_h I__2248 (
            .O(N__15737),
            .I(N__15731));
    Span4Mux_h I__2247 (
            .O(N__15734),
            .I(N__15728));
    Odrv4 I__2246 (
            .O(N__15731),
            .I(\this_sprites_ram.mem_WE_8 ));
    Odrv4 I__2245 (
            .O(N__15728),
            .I(\this_sprites_ram.mem_WE_8 ));
    InMux I__2244 (
            .O(N__15723),
            .I(N__15720));
    LocalMux I__2243 (
            .O(N__15720),
            .I(N__15717));
    Odrv12 I__2242 (
            .O(N__15717),
            .I(M_this_map_ram_write_data_2));
    InMux I__2241 (
            .O(N__15714),
            .I(N__15711));
    LocalMux I__2240 (
            .O(N__15711),
            .I(N__15707));
    InMux I__2239 (
            .O(N__15710),
            .I(N__15704));
    Span4Mux_h I__2238 (
            .O(N__15707),
            .I(N__15698));
    LocalMux I__2237 (
            .O(N__15704),
            .I(N__15698));
    InMux I__2236 (
            .O(N__15703),
            .I(N__15695));
    Odrv4 I__2235 (
            .O(N__15698),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__2234 (
            .O(N__15695),
            .I(\this_vga_signals.vaddress_c2 ));
    InMux I__2233 (
            .O(N__15690),
            .I(N__15687));
    LocalMux I__2232 (
            .O(N__15687),
            .I(N__15684));
    Span4Mux_h I__2231 (
            .O(N__15684),
            .I(N__15681));
    Odrv4 I__2230 (
            .O(N__15681),
            .I(\this_vga_signals.g0_0_0_0 ));
    InMux I__2229 (
            .O(N__15678),
            .I(N__15674));
    InMux I__2228 (
            .O(N__15677),
            .I(N__15669));
    LocalMux I__2227 (
            .O(N__15674),
            .I(N__15666));
    InMux I__2226 (
            .O(N__15673),
            .I(N__15663));
    InMux I__2225 (
            .O(N__15672),
            .I(N__15660));
    LocalMux I__2224 (
            .O(N__15669),
            .I(N__15657));
    Span4Mux_v I__2223 (
            .O(N__15666),
            .I(N__15649));
    LocalMux I__2222 (
            .O(N__15663),
            .I(N__15649));
    LocalMux I__2221 (
            .O(N__15660),
            .I(N__15646));
    Span4Mux_h I__2220 (
            .O(N__15657),
            .I(N__15643));
    InMux I__2219 (
            .O(N__15656),
            .I(N__15640));
    CascadeMux I__2218 (
            .O(N__15655),
            .I(N__15637));
    InMux I__2217 (
            .O(N__15654),
            .I(N__15632));
    Span4Mux_h I__2216 (
            .O(N__15649),
            .I(N__15629));
    Span4Mux_h I__2215 (
            .O(N__15646),
            .I(N__15622));
    Span4Mux_v I__2214 (
            .O(N__15643),
            .I(N__15622));
    LocalMux I__2213 (
            .O(N__15640),
            .I(N__15622));
    InMux I__2212 (
            .O(N__15637),
            .I(N__15617));
    InMux I__2211 (
            .O(N__15636),
            .I(N__15617));
    InMux I__2210 (
            .O(N__15635),
            .I(N__15614));
    LocalMux I__2209 (
            .O(N__15632),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2208 (
            .O(N__15629),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2207 (
            .O(N__15622),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2206 (
            .O(N__15617),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2205 (
            .O(N__15614),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    CascadeMux I__2204 (
            .O(N__15603),
            .I(\this_vga_signals.g2_0_0_cascade_ ));
    InMux I__2203 (
            .O(N__15600),
            .I(N__15594));
    InMux I__2202 (
            .O(N__15599),
            .I(N__15591));
    InMux I__2201 (
            .O(N__15598),
            .I(N__15588));
    InMux I__2200 (
            .O(N__15597),
            .I(N__15585));
    LocalMux I__2199 (
            .O(N__15594),
            .I(N__15582));
    LocalMux I__2198 (
            .O(N__15591),
            .I(N__15575));
    LocalMux I__2197 (
            .O(N__15588),
            .I(N__15575));
    LocalMux I__2196 (
            .O(N__15585),
            .I(N__15572));
    Span4Mux_h I__2195 (
            .O(N__15582),
            .I(N__15569));
    InMux I__2194 (
            .O(N__15581),
            .I(N__15563));
    InMux I__2193 (
            .O(N__15580),
            .I(N__15560));
    Span4Mux_h I__2192 (
            .O(N__15575),
            .I(N__15557));
    Span4Mux_h I__2191 (
            .O(N__15572),
            .I(N__15552));
    Span4Mux_v I__2190 (
            .O(N__15569),
            .I(N__15552));
    InMux I__2189 (
            .O(N__15568),
            .I(N__15549));
    InMux I__2188 (
            .O(N__15567),
            .I(N__15544));
    InMux I__2187 (
            .O(N__15566),
            .I(N__15544));
    LocalMux I__2186 (
            .O(N__15563),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2185 (
            .O(N__15560),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__2184 (
            .O(N__15557),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__2183 (
            .O(N__15552),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2182 (
            .O(N__15549),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2181 (
            .O(N__15544),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__2180 (
            .O(N__15531),
            .I(N__15528));
    LocalMux I__2179 (
            .O(N__15528),
            .I(N__15525));
    Span12Mux_h I__2178 (
            .O(N__15525),
            .I(N__15522));
    Odrv12 I__2177 (
            .O(N__15522),
            .I(\this_vga_signals.g0_2_0 ));
    InMux I__2176 (
            .O(N__15519),
            .I(N__15513));
    InMux I__2175 (
            .O(N__15518),
            .I(N__15508));
    InMux I__2174 (
            .O(N__15517),
            .I(N__15508));
    InMux I__2173 (
            .O(N__15516),
            .I(N__15505));
    LocalMux I__2172 (
            .O(N__15513),
            .I(\this_vga_signals.mult1_un40_sum_axb1_0 ));
    LocalMux I__2171 (
            .O(N__15508),
            .I(\this_vga_signals.mult1_un40_sum_axb1_0 ));
    LocalMux I__2170 (
            .O(N__15505),
            .I(\this_vga_signals.mult1_un40_sum_axb1_0 ));
    InMux I__2169 (
            .O(N__15498),
            .I(N__15495));
    LocalMux I__2168 (
            .O(N__15495),
            .I(N__15491));
    InMux I__2167 (
            .O(N__15494),
            .I(N__15486));
    Span4Mux_v I__2166 (
            .O(N__15491),
            .I(N__15483));
    InMux I__2165 (
            .O(N__15490),
            .I(N__15480));
    InMux I__2164 (
            .O(N__15489),
            .I(N__15477));
    LocalMux I__2163 (
            .O(N__15486),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    Odrv4 I__2162 (
            .O(N__15483),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    LocalMux I__2161 (
            .O(N__15480),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    LocalMux I__2160 (
            .O(N__15477),
            .I(\this_vga_signals.SUM_2_i_1_0_3 ));
    CascadeMux I__2159 (
            .O(N__15468),
            .I(N__15465));
    InMux I__2158 (
            .O(N__15465),
            .I(N__15461));
    CascadeMux I__2157 (
            .O(N__15464),
            .I(N__15457));
    LocalMux I__2156 (
            .O(N__15461),
            .I(N__15454));
    CascadeMux I__2155 (
            .O(N__15460),
            .I(N__15451));
    InMux I__2154 (
            .O(N__15457),
            .I(N__15448));
    Span4Mux_h I__2153 (
            .O(N__15454),
            .I(N__15445));
    InMux I__2152 (
            .O(N__15451),
            .I(N__15442));
    LocalMux I__2151 (
            .O(N__15448),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    Odrv4 I__2150 (
            .O(N__15445),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    LocalMux I__2149 (
            .O(N__15442),
            .I(\this_vga_signals.SUM_2_i_1_2_3 ));
    InMux I__2148 (
            .O(N__15435),
            .I(N__15432));
    LocalMux I__2147 (
            .O(N__15432),
            .I(N__15429));
    Span4Mux_h I__2146 (
            .O(N__15429),
            .I(N__15423));
    InMux I__2145 (
            .O(N__15428),
            .I(N__15418));
    InMux I__2144 (
            .O(N__15427),
            .I(N__15418));
    InMux I__2143 (
            .O(N__15426),
            .I(N__15415));
    Odrv4 I__2142 (
            .O(N__15423),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ));
    LocalMux I__2141 (
            .O(N__15418),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ));
    LocalMux I__2140 (
            .O(N__15415),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ));
    InMux I__2139 (
            .O(N__15408),
            .I(N__15398));
    InMux I__2138 (
            .O(N__15407),
            .I(N__15398));
    InMux I__2137 (
            .O(N__15406),
            .I(N__15398));
    InMux I__2136 (
            .O(N__15405),
            .I(N__15395));
    LocalMux I__2135 (
            .O(N__15398),
            .I(N__15390));
    LocalMux I__2134 (
            .O(N__15395),
            .I(N__15387));
    CascadeMux I__2133 (
            .O(N__15394),
            .I(N__15381));
    InMux I__2132 (
            .O(N__15393),
            .I(N__15378));
    Span4Mux_v I__2131 (
            .O(N__15390),
            .I(N__15375));
    Span4Mux_h I__2130 (
            .O(N__15387),
            .I(N__15372));
    InMux I__2129 (
            .O(N__15386),
            .I(N__15369));
    InMux I__2128 (
            .O(N__15385),
            .I(N__15362));
    InMux I__2127 (
            .O(N__15384),
            .I(N__15362));
    InMux I__2126 (
            .O(N__15381),
            .I(N__15362));
    LocalMux I__2125 (
            .O(N__15378),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__2124 (
            .O(N__15375),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__2123 (
            .O(N__15372),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2122 (
            .O(N__15369),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2121 (
            .O(N__15362),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    CascadeMux I__2120 (
            .O(N__15351),
            .I(\this_vga_signals.vaddress_0_0_6_cascade_ ));
    InMux I__2119 (
            .O(N__15348),
            .I(N__15345));
    LocalMux I__2118 (
            .O(N__15345),
            .I(N__15342));
    Span4Mux_v I__2117 (
            .O(N__15342),
            .I(N__15339));
    Odrv4 I__2116 (
            .O(N__15339),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_0_0 ));
    CascadeMux I__2115 (
            .O(N__15336),
            .I(N__15333));
    InMux I__2114 (
            .O(N__15333),
            .I(N__15328));
    InMux I__2113 (
            .O(N__15332),
            .I(N__15322));
    InMux I__2112 (
            .O(N__15331),
            .I(N__15319));
    LocalMux I__2111 (
            .O(N__15328),
            .I(N__15313));
    InMux I__2110 (
            .O(N__15327),
            .I(N__15310));
    InMux I__2109 (
            .O(N__15326),
            .I(N__15307));
    InMux I__2108 (
            .O(N__15325),
            .I(N__15304));
    LocalMux I__2107 (
            .O(N__15322),
            .I(N__15299));
    LocalMux I__2106 (
            .O(N__15319),
            .I(N__15299));
    InMux I__2105 (
            .O(N__15318),
            .I(N__15294));
    InMux I__2104 (
            .O(N__15317),
            .I(N__15294));
    InMux I__2103 (
            .O(N__15316),
            .I(N__15291));
    Odrv4 I__2102 (
            .O(N__15313),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2101 (
            .O(N__15310),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2100 (
            .O(N__15307),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2099 (
            .O(N__15304),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__2098 (
            .O(N__15299),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2097 (
            .O(N__15294),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2096 (
            .O(N__15291),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__2095 (
            .O(N__15276),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__2094 (
            .O(N__15273),
            .I(N__15269));
    CascadeMux I__2093 (
            .O(N__15272),
            .I(N__15266));
    LocalMux I__2092 (
            .O(N__15269),
            .I(N__15260));
    InMux I__2091 (
            .O(N__15266),
            .I(N__15257));
    CascadeMux I__2090 (
            .O(N__15265),
            .I(N__15250));
    CascadeMux I__2089 (
            .O(N__15264),
            .I(N__15247));
    CascadeMux I__2088 (
            .O(N__15263),
            .I(N__15244));
    Span4Mux_v I__2087 (
            .O(N__15260),
            .I(N__15239));
    LocalMux I__2086 (
            .O(N__15257),
            .I(N__15239));
    InMux I__2085 (
            .O(N__15256),
            .I(N__15236));
    InMux I__2084 (
            .O(N__15255),
            .I(N__15232));
    InMux I__2083 (
            .O(N__15254),
            .I(N__15229));
    InMux I__2082 (
            .O(N__15253),
            .I(N__15220));
    InMux I__2081 (
            .O(N__15250),
            .I(N__15220));
    InMux I__2080 (
            .O(N__15247),
            .I(N__15220));
    InMux I__2079 (
            .O(N__15244),
            .I(N__15220));
    Span4Mux_h I__2078 (
            .O(N__15239),
            .I(N__15215));
    LocalMux I__2077 (
            .O(N__15236),
            .I(N__15215));
    InMux I__2076 (
            .O(N__15235),
            .I(N__15212));
    LocalMux I__2075 (
            .O(N__15232),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2074 (
            .O(N__15229),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2073 (
            .O(N__15220),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__2072 (
            .O(N__15215),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2071 (
            .O(N__15212),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__2070 (
            .O(N__15201),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__2069 (
            .O(N__15198),
            .I(N__15192));
    InMux I__2068 (
            .O(N__15197),
            .I(N__15187));
    InMux I__2067 (
            .O(N__15196),
            .I(N__15182));
    InMux I__2066 (
            .O(N__15195),
            .I(N__15182));
    LocalMux I__2065 (
            .O(N__15192),
            .I(N__15174));
    InMux I__2064 (
            .O(N__15191),
            .I(N__15171));
    InMux I__2063 (
            .O(N__15190),
            .I(N__15168));
    LocalMux I__2062 (
            .O(N__15187),
            .I(N__15165));
    LocalMux I__2061 (
            .O(N__15182),
            .I(N__15162));
    InMux I__2060 (
            .O(N__15181),
            .I(N__15157));
    InMux I__2059 (
            .O(N__15180),
            .I(N__15157));
    InMux I__2058 (
            .O(N__15179),
            .I(N__15154));
    InMux I__2057 (
            .O(N__15178),
            .I(N__15151));
    InMux I__2056 (
            .O(N__15177),
            .I(N__15148));
    Odrv4 I__2055 (
            .O(N__15174),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2054 (
            .O(N__15171),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2053 (
            .O(N__15168),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__2052 (
            .O(N__15165),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__2051 (
            .O(N__15162),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2050 (
            .O(N__15157),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2049 (
            .O(N__15154),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2048 (
            .O(N__15151),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2047 (
            .O(N__15148),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__2046 (
            .O(N__15129),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__2045 (
            .O(N__15126),
            .I(N__15121));
    CascadeMux I__2044 (
            .O(N__15125),
            .I(N__15116));
    InMux I__2043 (
            .O(N__15124),
            .I(N__15107));
    LocalMux I__2042 (
            .O(N__15121),
            .I(N__15104));
    InMux I__2041 (
            .O(N__15120),
            .I(N__15097));
    InMux I__2040 (
            .O(N__15119),
            .I(N__15097));
    InMux I__2039 (
            .O(N__15116),
            .I(N__15097));
    InMux I__2038 (
            .O(N__15115),
            .I(N__15092));
    InMux I__2037 (
            .O(N__15114),
            .I(N__15092));
    InMux I__2036 (
            .O(N__15113),
            .I(N__15083));
    InMux I__2035 (
            .O(N__15112),
            .I(N__15083));
    InMux I__2034 (
            .O(N__15111),
            .I(N__15083));
    InMux I__2033 (
            .O(N__15110),
            .I(N__15083));
    LocalMux I__2032 (
            .O(N__15107),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2031 (
            .O(N__15104),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2030 (
            .O(N__15097),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2029 (
            .O(N__15092),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2028 (
            .O(N__15083),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    InMux I__2027 (
            .O(N__15072),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__2026 (
            .O(N__15069),
            .I(N__15066));
    LocalMux I__2025 (
            .O(N__15066),
            .I(N__15060));
    CascadeMux I__2024 (
            .O(N__15065),
            .I(N__15051));
    CascadeMux I__2023 (
            .O(N__15064),
            .I(N__15048));
    InMux I__2022 (
            .O(N__15063),
            .I(N__15045));
    Span4Mux_h I__2021 (
            .O(N__15060),
            .I(N__15042));
    InMux I__2020 (
            .O(N__15059),
            .I(N__15037));
    InMux I__2019 (
            .O(N__15058),
            .I(N__15037));
    InMux I__2018 (
            .O(N__15057),
            .I(N__15028));
    InMux I__2017 (
            .O(N__15056),
            .I(N__15028));
    InMux I__2016 (
            .O(N__15055),
            .I(N__15028));
    InMux I__2015 (
            .O(N__15054),
            .I(N__15028));
    InMux I__2014 (
            .O(N__15051),
            .I(N__15023));
    InMux I__2013 (
            .O(N__15048),
            .I(N__15023));
    LocalMux I__2012 (
            .O(N__15045),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__2011 (
            .O(N__15042),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2010 (
            .O(N__15037),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2009 (
            .O(N__15028),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2008 (
            .O(N__15023),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__2007 (
            .O(N__15012),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__2006 (
            .O(N__15009),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__2005 (
            .O(N__15006),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__2004 (
            .O(N__15003),
            .I(N__15000));
    LocalMux I__2003 (
            .O(N__15000),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_0 ));
    CascadeMux I__2002 (
            .O(N__14997),
            .I(\this_vga_signals.mult1_un54_sum_c3_1_0_cascade_ ));
    InMux I__2001 (
            .O(N__14994),
            .I(N__14991));
    LocalMux I__2000 (
            .O(N__14991),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1 ));
    InMux I__1999 (
            .O(N__14988),
            .I(N__14982));
    CascadeMux I__1998 (
            .O(N__14987),
            .I(N__14977));
    CascadeMux I__1997 (
            .O(N__14986),
            .I(N__14974));
    InMux I__1996 (
            .O(N__14985),
            .I(N__14969));
    LocalMux I__1995 (
            .O(N__14982),
            .I(N__14966));
    InMux I__1994 (
            .O(N__14981),
            .I(N__14963));
    InMux I__1993 (
            .O(N__14980),
            .I(N__14960));
    InMux I__1992 (
            .O(N__14977),
            .I(N__14955));
    InMux I__1991 (
            .O(N__14974),
            .I(N__14955));
    CascadeMux I__1990 (
            .O(N__14973),
            .I(N__14952));
    InMux I__1989 (
            .O(N__14972),
            .I(N__14949));
    LocalMux I__1988 (
            .O(N__14969),
            .I(N__14939));
    Span4Mux_h I__1987 (
            .O(N__14966),
            .I(N__14939));
    LocalMux I__1986 (
            .O(N__14963),
            .I(N__14932));
    LocalMux I__1985 (
            .O(N__14960),
            .I(N__14932));
    LocalMux I__1984 (
            .O(N__14955),
            .I(N__14932));
    InMux I__1983 (
            .O(N__14952),
            .I(N__14929));
    LocalMux I__1982 (
            .O(N__14949),
            .I(N__14926));
    InMux I__1981 (
            .O(N__14948),
            .I(N__14923));
    InMux I__1980 (
            .O(N__14947),
            .I(N__14920));
    InMux I__1979 (
            .O(N__14946),
            .I(N__14915));
    InMux I__1978 (
            .O(N__14945),
            .I(N__14915));
    InMux I__1977 (
            .O(N__14944),
            .I(N__14912));
    Span4Mux_v I__1976 (
            .O(N__14939),
            .I(N__14909));
    Span4Mux_v I__1975 (
            .O(N__14932),
            .I(N__14906));
    LocalMux I__1974 (
            .O(N__14929),
            .I(N__14901));
    Span4Mux_h I__1973 (
            .O(N__14926),
            .I(N__14901));
    LocalMux I__1972 (
            .O(N__14923),
            .I(N__14896));
    LocalMux I__1971 (
            .O(N__14920),
            .I(N__14896));
    LocalMux I__1970 (
            .O(N__14915),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1969 (
            .O(N__14912),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1968 (
            .O(N__14909),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1967 (
            .O(N__14906),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1966 (
            .O(N__14901),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv12 I__1965 (
            .O(N__14896),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__1964 (
            .O(N__14883),
            .I(N__14880));
    LocalMux I__1963 (
            .O(N__14880),
            .I(N__14877));
    Span4Mux_h I__1962 (
            .O(N__14877),
            .I(N__14869));
    InMux I__1961 (
            .O(N__14876),
            .I(N__14864));
    InMux I__1960 (
            .O(N__14875),
            .I(N__14864));
    InMux I__1959 (
            .O(N__14874),
            .I(N__14861));
    InMux I__1958 (
            .O(N__14873),
            .I(N__14858));
    InMux I__1957 (
            .O(N__14872),
            .I(N__14855));
    Span4Mux_v I__1956 (
            .O(N__14869),
            .I(N__14852));
    LocalMux I__1955 (
            .O(N__14864),
            .I(N__14847));
    LocalMux I__1954 (
            .O(N__14861),
            .I(N__14847));
    LocalMux I__1953 (
            .O(N__14858),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__1952 (
            .O(N__14855),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__1951 (
            .O(N__14852),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv12 I__1950 (
            .O(N__14847),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    InMux I__1949 (
            .O(N__14838),
            .I(N__14835));
    LocalMux I__1948 (
            .O(N__14835),
            .I(\this_vga_signals.mult1_un68_sum_axb1 ));
    InMux I__1947 (
            .O(N__14832),
            .I(N__14829));
    LocalMux I__1946 (
            .O(N__14829),
            .I(\this_vga_signals.if_m5_s ));
    CascadeMux I__1945 (
            .O(N__14826),
            .I(N__14822));
    CascadeMux I__1944 (
            .O(N__14825),
            .I(N__14819));
    InMux I__1943 (
            .O(N__14822),
            .I(N__14816));
    InMux I__1942 (
            .O(N__14819),
            .I(N__14813));
    LocalMux I__1941 (
            .O(N__14816),
            .I(N__14810));
    LocalMux I__1940 (
            .O(N__14813),
            .I(N__14805));
    Span4Mux_v I__1939 (
            .O(N__14810),
            .I(N__14805));
    Span4Mux_h I__1938 (
            .O(N__14805),
            .I(N__14802));
    Odrv4 I__1937 (
            .O(N__14802),
            .I(\this_vga_signals.M_vcounter_d7lto8_1 ));
    InMux I__1936 (
            .O(N__14799),
            .I(N__14794));
    InMux I__1935 (
            .O(N__14798),
            .I(N__14787));
    CascadeMux I__1934 (
            .O(N__14797),
            .I(N__14784));
    LocalMux I__1933 (
            .O(N__14794),
            .I(N__14780));
    InMux I__1932 (
            .O(N__14793),
            .I(N__14777));
    InMux I__1931 (
            .O(N__14792),
            .I(N__14772));
    InMux I__1930 (
            .O(N__14791),
            .I(N__14772));
    InMux I__1929 (
            .O(N__14790),
            .I(N__14767));
    LocalMux I__1928 (
            .O(N__14787),
            .I(N__14764));
    InMux I__1927 (
            .O(N__14784),
            .I(N__14759));
    InMux I__1926 (
            .O(N__14783),
            .I(N__14759));
    Span4Mux_v I__1925 (
            .O(N__14780),
            .I(N__14754));
    LocalMux I__1924 (
            .O(N__14777),
            .I(N__14754));
    LocalMux I__1923 (
            .O(N__14772),
            .I(N__14749));
    InMux I__1922 (
            .O(N__14771),
            .I(N__14746));
    CascadeMux I__1921 (
            .O(N__14770),
            .I(N__14743));
    LocalMux I__1920 (
            .O(N__14767),
            .I(N__14732));
    Span4Mux_v I__1919 (
            .O(N__14764),
            .I(N__14732));
    LocalMux I__1918 (
            .O(N__14759),
            .I(N__14732));
    Span4Mux_v I__1917 (
            .O(N__14754),
            .I(N__14732));
    InMux I__1916 (
            .O(N__14753),
            .I(N__14729));
    InMux I__1915 (
            .O(N__14752),
            .I(N__14726));
    Span4Mux_v I__1914 (
            .O(N__14749),
            .I(N__14721));
    LocalMux I__1913 (
            .O(N__14746),
            .I(N__14721));
    InMux I__1912 (
            .O(N__14743),
            .I(N__14718));
    InMux I__1911 (
            .O(N__14742),
            .I(N__14713));
    InMux I__1910 (
            .O(N__14741),
            .I(N__14713));
    Odrv4 I__1909 (
            .O(N__14732),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1908 (
            .O(N__14729),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1907 (
            .O(N__14726),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__1906 (
            .O(N__14721),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1905 (
            .O(N__14718),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__1904 (
            .O(N__14713),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    IoInMux I__1903 (
            .O(N__14700),
            .I(N__14697));
    LocalMux I__1902 (
            .O(N__14697),
            .I(N__14694));
    IoSpan4Mux I__1901 (
            .O(N__14694),
            .I(N__14691));
    Span4Mux_s3_v I__1900 (
            .O(N__14691),
            .I(N__14688));
    Sp12to4 I__1899 (
            .O(N__14688),
            .I(N__14684));
    InMux I__1898 (
            .O(N__14687),
            .I(N__14681));
    Span12Mux_v I__1897 (
            .O(N__14684),
            .I(N__14678));
    LocalMux I__1896 (
            .O(N__14681),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ));
    Odrv12 I__1895 (
            .O(N__14678),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ));
    InMux I__1894 (
            .O(N__14673),
            .I(N__14670));
    LocalMux I__1893 (
            .O(N__14670),
            .I(\this_vga_signals.M_hcounter_d7lto4_0 ));
    InMux I__1892 (
            .O(N__14667),
            .I(N__14664));
    LocalMux I__1891 (
            .O(N__14664),
            .I(N__14661));
    Span4Mux_v I__1890 (
            .O(N__14661),
            .I(N__14658));
    Sp12to4 I__1889 (
            .O(N__14658),
            .I(N__14655));
    Odrv12 I__1888 (
            .O(N__14655),
            .I(\this_sprites_ram.mem_out_bus7_0 ));
    InMux I__1887 (
            .O(N__14652),
            .I(N__14649));
    LocalMux I__1886 (
            .O(N__14649),
            .I(N__14646));
    Span4Mux_h I__1885 (
            .O(N__14646),
            .I(N__14643));
    Span4Mux_v I__1884 (
            .O(N__14643),
            .I(N__14640));
    Span4Mux_h I__1883 (
            .O(N__14640),
            .I(N__14637));
    Odrv4 I__1882 (
            .O(N__14637),
            .I(\this_sprites_ram.mem_out_bus3_0 ));
    CascadeMux I__1881 (
            .O(N__14634),
            .I(N__14631));
    InMux I__1880 (
            .O(N__14631),
            .I(N__14627));
    InMux I__1879 (
            .O(N__14630),
            .I(N__14621));
    LocalMux I__1878 (
            .O(N__14627),
            .I(N__14618));
    InMux I__1877 (
            .O(N__14626),
            .I(N__14615));
    InMux I__1876 (
            .O(N__14625),
            .I(N__14610));
    InMux I__1875 (
            .O(N__14624),
            .I(N__14610));
    LocalMux I__1874 (
            .O(N__14621),
            .I(N__14605));
    Span4Mux_h I__1873 (
            .O(N__14618),
            .I(N__14605));
    LocalMux I__1872 (
            .O(N__14615),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1871 (
            .O(N__14610),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    Odrv4 I__1870 (
            .O(N__14605),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    CascadeMux I__1869 (
            .O(N__14598),
            .I(N__14595));
    InMux I__1868 (
            .O(N__14595),
            .I(N__14592));
    LocalMux I__1867 (
            .O(N__14592),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_x0 ));
    InMux I__1866 (
            .O(N__14589),
            .I(N__14586));
    LocalMux I__1865 (
            .O(N__14586),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_x1 ));
    CascadeMux I__1864 (
            .O(N__14583),
            .I(\this_vga_signals.mult1_un68_sum_axb1_654_ns_cascade_ ));
    InMux I__1863 (
            .O(N__14580),
            .I(N__14577));
    LocalMux I__1862 (
            .O(N__14577),
            .I(\this_vga_signals.if_m1_3 ));
    CascadeMux I__1861 (
            .O(N__14574),
            .I(\this_vga_signals.if_m1_3_cascade_ ));
    CascadeMux I__1860 (
            .O(N__14571),
            .I(N__14568));
    InMux I__1859 (
            .O(N__14568),
            .I(N__14565));
    LocalMux I__1858 (
            .O(N__14565),
            .I(N__14562));
    Odrv4 I__1857 (
            .O(N__14562),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1 ));
    CascadeMux I__1856 (
            .O(N__14559),
            .I(N__14556));
    InMux I__1855 (
            .O(N__14556),
            .I(N__14553));
    LocalMux I__1854 (
            .O(N__14553),
            .I(N__14550));
    Span4Mux_h I__1853 (
            .O(N__14550),
            .I(N__14547));
    Odrv4 I__1852 (
            .O(N__14547),
            .I(\this_vga_signals.vaddress_0_6 ));
    InMux I__1851 (
            .O(N__14544),
            .I(N__14541));
    LocalMux I__1850 (
            .O(N__14541),
            .I(\this_vga_signals.mult1_un47_sum_c3_1_0 ));
    CascadeMux I__1849 (
            .O(N__14538),
            .I(N__14533));
    InMux I__1848 (
            .O(N__14537),
            .I(N__14529));
    InMux I__1847 (
            .O(N__14536),
            .I(N__14526));
    InMux I__1846 (
            .O(N__14533),
            .I(N__14523));
    InMux I__1845 (
            .O(N__14532),
            .I(N__14520));
    LocalMux I__1844 (
            .O(N__14529),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3 ));
    LocalMux I__1843 (
            .O(N__14526),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3 ));
    LocalMux I__1842 (
            .O(N__14523),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3 ));
    LocalMux I__1841 (
            .O(N__14520),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3 ));
    InMux I__1840 (
            .O(N__14511),
            .I(N__14508));
    LocalMux I__1839 (
            .O(N__14508),
            .I(\this_vga_signals.g1 ));
    InMux I__1838 (
            .O(N__14505),
            .I(N__14502));
    LocalMux I__1837 (
            .O(N__14502),
            .I(N__14489));
    InMux I__1836 (
            .O(N__14501),
            .I(N__14484));
    InMux I__1835 (
            .O(N__14500),
            .I(N__14481));
    InMux I__1834 (
            .O(N__14499),
            .I(N__14474));
    InMux I__1833 (
            .O(N__14498),
            .I(N__14474));
    InMux I__1832 (
            .O(N__14497),
            .I(N__14474));
    InMux I__1831 (
            .O(N__14496),
            .I(N__14467));
    InMux I__1830 (
            .O(N__14495),
            .I(N__14467));
    InMux I__1829 (
            .O(N__14494),
            .I(N__14467));
    InMux I__1828 (
            .O(N__14493),
            .I(N__14462));
    InMux I__1827 (
            .O(N__14492),
            .I(N__14462));
    Span4Mux_v I__1826 (
            .O(N__14489),
            .I(N__14459));
    InMux I__1825 (
            .O(N__14488),
            .I(N__14454));
    InMux I__1824 (
            .O(N__14487),
            .I(N__14454));
    LocalMux I__1823 (
            .O(N__14484),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1822 (
            .O(N__14481),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1821 (
            .O(N__14474),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1820 (
            .O(N__14467),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1819 (
            .O(N__14462),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    Odrv4 I__1818 (
            .O(N__14459),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1817 (
            .O(N__14454),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    CascadeMux I__1816 (
            .O(N__14439),
            .I(\this_vga_signals.g0_2_cascade_ ));
    InMux I__1815 (
            .O(N__14436),
            .I(N__14433));
    LocalMux I__1814 (
            .O(N__14433),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0_1 ));
    InMux I__1813 (
            .O(N__14430),
            .I(N__14427));
    LocalMux I__1812 (
            .O(N__14427),
            .I(\this_vga_signals.N_3_1_0 ));
    CascadeMux I__1811 (
            .O(N__14424),
            .I(\this_vga_signals.N_11_0_0_cascade_ ));
    InMux I__1810 (
            .O(N__14421),
            .I(N__14418));
    LocalMux I__1809 (
            .O(N__14418),
            .I(\this_vga_signals.N_4_1_0_0 ));
    InMux I__1808 (
            .O(N__14415),
            .I(N__14412));
    LocalMux I__1807 (
            .O(N__14412),
            .I(N__14409));
    Odrv4 I__1806 (
            .O(N__14409),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_2 ));
    CascadeMux I__1805 (
            .O(N__14406),
            .I(N__14403));
    InMux I__1804 (
            .O(N__14403),
            .I(N__14400));
    LocalMux I__1803 (
            .O(N__14400),
            .I(N__14397));
    Span4Mux_h I__1802 (
            .O(N__14397),
            .I(N__14393));
    InMux I__1801 (
            .O(N__14396),
            .I(N__14390));
    Odrv4 I__1800 (
            .O(N__14393),
            .I(\this_vga_signals.vaddress_3_6 ));
    LocalMux I__1799 (
            .O(N__14390),
            .I(\this_vga_signals.vaddress_3_6 ));
    CascadeMux I__1798 (
            .O(N__14385),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i_2_cascade_ ));
    InMux I__1797 (
            .O(N__14382),
            .I(N__14379));
    LocalMux I__1796 (
            .O(N__14379),
            .I(\this_vga_signals.mult1_un47_sum_c3_2 ));
    CascadeMux I__1795 (
            .O(N__14376),
            .I(\this_vga_signals.mult1_un47_sum_c3_2_cascade_ ));
    InMux I__1794 (
            .O(N__14373),
            .I(N__14370));
    LocalMux I__1793 (
            .O(N__14370),
            .I(\this_vga_signals.g0_1 ));
    InMux I__1792 (
            .O(N__14367),
            .I(N__14361));
    InMux I__1791 (
            .O(N__14366),
            .I(N__14356));
    InMux I__1790 (
            .O(N__14365),
            .I(N__14356));
    CascadeMux I__1789 (
            .O(N__14364),
            .I(N__14350));
    LocalMux I__1788 (
            .O(N__14361),
            .I(N__14345));
    LocalMux I__1787 (
            .O(N__14356),
            .I(N__14345));
    InMux I__1786 (
            .O(N__14355),
            .I(N__14342));
    InMux I__1785 (
            .O(N__14354),
            .I(N__14339));
    InMux I__1784 (
            .O(N__14353),
            .I(N__14334));
    InMux I__1783 (
            .O(N__14350),
            .I(N__14334));
    Span4Mux_h I__1782 (
            .O(N__14345),
            .I(N__14331));
    LocalMux I__1781 (
            .O(N__14342),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1780 (
            .O(N__14339),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1779 (
            .O(N__14334),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__1778 (
            .O(N__14331),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    CascadeMux I__1777 (
            .O(N__14322),
            .I(\this_vga_signals.vaddress_6_cascade_ ));
    CascadeMux I__1776 (
            .O(N__14319),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ));
    InMux I__1775 (
            .O(N__14316),
            .I(N__14313));
    LocalMux I__1774 (
            .O(N__14313),
            .I(N__14310));
    Odrv4 I__1773 (
            .O(N__14310),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_i ));
    InMux I__1772 (
            .O(N__14307),
            .I(N__14304));
    LocalMux I__1771 (
            .O(N__14304),
            .I(N__14301));
    Span4Mux_h I__1770 (
            .O(N__14301),
            .I(N__14296));
    InMux I__1769 (
            .O(N__14300),
            .I(N__14293));
    InMux I__1768 (
            .O(N__14299),
            .I(N__14290));
    Odrv4 I__1767 (
            .O(N__14296),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    LocalMux I__1766 (
            .O(N__14293),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    LocalMux I__1765 (
            .O(N__14290),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3 ));
    InMux I__1764 (
            .O(N__14283),
            .I(N__14280));
    LocalMux I__1763 (
            .O(N__14280),
            .I(N__14277));
    Span4Mux_v I__1762 (
            .O(N__14277),
            .I(N__14274));
    Span4Mux_h I__1761 (
            .O(N__14274),
            .I(N__14270));
    InMux I__1760 (
            .O(N__14273),
            .I(N__14267));
    Odrv4 I__1759 (
            .O(N__14270),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    LocalMux I__1758 (
            .O(N__14267),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__1757 (
            .O(N__14262),
            .I(N__14259));
    LocalMux I__1756 (
            .O(N__14259),
            .I(N__14256));
    Span4Mux_v I__1755 (
            .O(N__14256),
            .I(N__14251));
    InMux I__1754 (
            .O(N__14255),
            .I(N__14246));
    InMux I__1753 (
            .O(N__14254),
            .I(N__14246));
    Odrv4 I__1752 (
            .O(N__14251),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    LocalMux I__1751 (
            .O(N__14246),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    CascadeMux I__1750 (
            .O(N__14241),
            .I(N__14234));
    InMux I__1749 (
            .O(N__14240),
            .I(N__14229));
    InMux I__1748 (
            .O(N__14239),
            .I(N__14229));
    InMux I__1747 (
            .O(N__14238),
            .I(N__14226));
    InMux I__1746 (
            .O(N__14237),
            .I(N__14221));
    InMux I__1745 (
            .O(N__14234),
            .I(N__14221));
    LocalMux I__1744 (
            .O(N__14229),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1743 (
            .O(N__14226),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1742 (
            .O(N__14221),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    CascadeMux I__1741 (
            .O(N__14214),
            .I(N__14210));
    CascadeMux I__1740 (
            .O(N__14213),
            .I(N__14207));
    InMux I__1739 (
            .O(N__14210),
            .I(N__14200));
    InMux I__1738 (
            .O(N__14207),
            .I(N__14200));
    CascadeMux I__1737 (
            .O(N__14206),
            .I(N__14197));
    InMux I__1736 (
            .O(N__14205),
            .I(N__14193));
    LocalMux I__1735 (
            .O(N__14200),
            .I(N__14190));
    InMux I__1734 (
            .O(N__14197),
            .I(N__14185));
    InMux I__1733 (
            .O(N__14196),
            .I(N__14185));
    LocalMux I__1732 (
            .O(N__14193),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    Odrv4 I__1731 (
            .O(N__14190),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1730 (
            .O(N__14185),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    InMux I__1729 (
            .O(N__14178),
            .I(N__14172));
    InMux I__1728 (
            .O(N__14177),
            .I(N__14172));
    LocalMux I__1727 (
            .O(N__14172),
            .I(N__14169));
    Span4Mux_h I__1726 (
            .O(N__14169),
            .I(N__14165));
    InMux I__1725 (
            .O(N__14168),
            .I(N__14162));
    Odrv4 I__1724 (
            .O(N__14165),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__1723 (
            .O(N__14162),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    CEMux I__1722 (
            .O(N__14157),
            .I(N__14151));
    CEMux I__1721 (
            .O(N__14156),
            .I(N__14147));
    CEMux I__1720 (
            .O(N__14155),
            .I(N__14144));
    CEMux I__1719 (
            .O(N__14154),
            .I(N__14141));
    LocalMux I__1718 (
            .O(N__14151),
            .I(N__14138));
    CEMux I__1717 (
            .O(N__14150),
            .I(N__14135));
    LocalMux I__1716 (
            .O(N__14147),
            .I(N__14132));
    LocalMux I__1715 (
            .O(N__14144),
            .I(N__14129));
    LocalMux I__1714 (
            .O(N__14141),
            .I(N__14122));
    Span4Mux_h I__1713 (
            .O(N__14138),
            .I(N__14122));
    LocalMux I__1712 (
            .O(N__14135),
            .I(N__14122));
    Span4Mux_v I__1711 (
            .O(N__14132),
            .I(N__14119));
    Span4Mux_v I__1710 (
            .O(N__14129),
            .I(N__14114));
    Span4Mux_v I__1709 (
            .O(N__14122),
            .I(N__14114));
    Odrv4 I__1708 (
            .O(N__14119),
            .I(\this_vga_signals.N_966_0 ));
    Odrv4 I__1707 (
            .O(N__14114),
            .I(\this_vga_signals.N_966_0 ));
    SRMux I__1706 (
            .O(N__14109),
            .I(N__14091));
    SRMux I__1705 (
            .O(N__14108),
            .I(N__14091));
    SRMux I__1704 (
            .O(N__14107),
            .I(N__14091));
    SRMux I__1703 (
            .O(N__14106),
            .I(N__14091));
    SRMux I__1702 (
            .O(N__14105),
            .I(N__14091));
    SRMux I__1701 (
            .O(N__14104),
            .I(N__14091));
    GlobalMux I__1700 (
            .O(N__14091),
            .I(N__14088));
    gio2CtrlBuf I__1699 (
            .O(N__14088),
            .I(\this_vga_signals.N_1332_g ));
    InMux I__1698 (
            .O(N__14085),
            .I(N__14082));
    LocalMux I__1697 (
            .O(N__14082),
            .I(N__14079));
    Span4Mux_h I__1696 (
            .O(N__14079),
            .I(N__14076));
    Odrv4 I__1695 (
            .O(N__14076),
            .I(\this_vga_signals.g1_0_0_0_0 ));
    InMux I__1694 (
            .O(N__14073),
            .I(N__14070));
    LocalMux I__1693 (
            .O(N__14070),
            .I(N__14067));
    Span4Mux_h I__1692 (
            .O(N__14067),
            .I(N__14064));
    Odrv4 I__1691 (
            .O(N__14064),
            .I(\this_vga_signals.g0_2_2_1 ));
    CascadeMux I__1690 (
            .O(N__14061),
            .I(\this_vga_signals.N_473_0_cascade_ ));
    InMux I__1689 (
            .O(N__14058),
            .I(N__14055));
    LocalMux I__1688 (
            .O(N__14055),
            .I(\this_vga_signals.N_554 ));
    InMux I__1687 (
            .O(N__14052),
            .I(N__14048));
    InMux I__1686 (
            .O(N__14051),
            .I(N__14045));
    LocalMux I__1685 (
            .O(N__14048),
            .I(\this_vga_signals.SUM_3_i_1_0 ));
    LocalMux I__1684 (
            .O(N__14045),
            .I(\this_vga_signals.SUM_3_i_1_0 ));
    CascadeMux I__1683 (
            .O(N__14040),
            .I(\this_vga_signals.N_735_0_cascade_ ));
    CascadeMux I__1682 (
            .O(N__14037),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_2_cascade_ ));
    InMux I__1681 (
            .O(N__14034),
            .I(N__14027));
    InMux I__1680 (
            .O(N__14033),
            .I(N__14027));
    InMux I__1679 (
            .O(N__14032),
            .I(N__14024));
    LocalMux I__1678 (
            .O(N__14027),
            .I(\this_vga_signals.N_735_0 ));
    LocalMux I__1677 (
            .O(N__14024),
            .I(\this_vga_signals.N_735_0 ));
    InMux I__1676 (
            .O(N__14019),
            .I(N__14016));
    LocalMux I__1675 (
            .O(N__14016),
            .I(N__14012));
    InMux I__1674 (
            .O(N__14015),
            .I(N__14009));
    Span4Mux_h I__1673 (
            .O(N__14012),
            .I(N__14003));
    LocalMux I__1672 (
            .O(N__14009),
            .I(N__14000));
    InMux I__1671 (
            .O(N__14008),
            .I(N__13997));
    InMux I__1670 (
            .O(N__14007),
            .I(N__13992));
    InMux I__1669 (
            .O(N__14006),
            .I(N__13992));
    Odrv4 I__1668 (
            .O(N__14003),
            .I(\this_vga_signals.mult1_un61_sum_0_3 ));
    Odrv4 I__1667 (
            .O(N__14000),
            .I(\this_vga_signals.mult1_un61_sum_0_3 ));
    LocalMux I__1666 (
            .O(N__13997),
            .I(\this_vga_signals.mult1_un61_sum_0_3 ));
    LocalMux I__1665 (
            .O(N__13992),
            .I(\this_vga_signals.mult1_un61_sum_0_3 ));
    InMux I__1664 (
            .O(N__13983),
            .I(N__13980));
    LocalMux I__1663 (
            .O(N__13980),
            .I(\this_vga_signals.hsync_1_i_0_1 ));
    CascadeMux I__1662 (
            .O(N__13977),
            .I(N__13974));
    InMux I__1661 (
            .O(N__13974),
            .I(N__13971));
    LocalMux I__1660 (
            .O(N__13971),
            .I(\this_vga_signals.N_507_0 ));
    InMux I__1659 (
            .O(N__13968),
            .I(N__13965));
    LocalMux I__1658 (
            .O(N__13965),
            .I(N__13962));
    Odrv12 I__1657 (
            .O(N__13962),
            .I(M_this_map_ram_write_data_6));
    InMux I__1656 (
            .O(N__13959),
            .I(N__13956));
    LocalMux I__1655 (
            .O(N__13956),
            .I(N__13953));
    Span4Mux_v I__1654 (
            .O(N__13953),
            .I(N__13948));
    InMux I__1653 (
            .O(N__13952),
            .I(N__13943));
    InMux I__1652 (
            .O(N__13951),
            .I(N__13943));
    Odrv4 I__1651 (
            .O(N__13948),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    LocalMux I__1650 (
            .O(N__13943),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    CascadeMux I__1649 (
            .O(N__13938),
            .I(N__13935));
    InMux I__1648 (
            .O(N__13935),
            .I(N__13932));
    LocalMux I__1647 (
            .O(N__13932),
            .I(N__13929));
    Span4Mux_v I__1646 (
            .O(N__13929),
            .I(N__13926));
    Odrv4 I__1645 (
            .O(N__13926),
            .I(\this_vga_signals.M_lcounter_d_0_sqmuxa ));
    CascadeMux I__1644 (
            .O(N__13923),
            .I(N__13918));
    InMux I__1643 (
            .O(N__13922),
            .I(N__13915));
    InMux I__1642 (
            .O(N__13921),
            .I(N__13912));
    InMux I__1641 (
            .O(N__13918),
            .I(N__13909));
    LocalMux I__1640 (
            .O(N__13915),
            .I(N__13905));
    LocalMux I__1639 (
            .O(N__13912),
            .I(N__13900));
    LocalMux I__1638 (
            .O(N__13909),
            .I(N__13900));
    InMux I__1637 (
            .O(N__13908),
            .I(N__13893));
    Span4Mux_v I__1636 (
            .O(N__13905),
            .I(N__13890));
    Span4Mux_v I__1635 (
            .O(N__13900),
            .I(N__13887));
    InMux I__1634 (
            .O(N__13899),
            .I(N__13880));
    InMux I__1633 (
            .O(N__13898),
            .I(N__13880));
    InMux I__1632 (
            .O(N__13897),
            .I(N__13880));
    InMux I__1631 (
            .O(N__13896),
            .I(N__13877));
    LocalMux I__1630 (
            .O(N__13893),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__1629 (
            .O(N__13890),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__1628 (
            .O(N__13887),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    LocalMux I__1627 (
            .O(N__13880),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    LocalMux I__1626 (
            .O(N__13877),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    InMux I__1625 (
            .O(N__13866),
            .I(N__13860));
    InMux I__1624 (
            .O(N__13865),
            .I(N__13860));
    LocalMux I__1623 (
            .O(N__13860),
            .I(N__13856));
    InMux I__1622 (
            .O(N__13859),
            .I(N__13853));
    Span4Mux_v I__1621 (
            .O(N__13856),
            .I(N__13850));
    LocalMux I__1620 (
            .O(N__13853),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    Odrv4 I__1619 (
            .O(N__13850),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    CascadeMux I__1618 (
            .O(N__13845),
            .I(\this_vga_signals.SUM_3_i_1_0_cascade_ ));
    InMux I__1617 (
            .O(N__13842),
            .I(N__13839));
    LocalMux I__1616 (
            .O(N__13839),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_1 ));
    CascadeMux I__1615 (
            .O(N__13836),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_1_cascade_ ));
    InMux I__1614 (
            .O(N__13833),
            .I(N__13830));
    LocalMux I__1613 (
            .O(N__13830),
            .I(\this_vga_signals.if_N_8_i_0 ));
    InMux I__1612 (
            .O(N__13827),
            .I(N__13824));
    LocalMux I__1611 (
            .O(N__13824),
            .I(N__13821));
    Odrv4 I__1610 (
            .O(N__13821),
            .I(\this_vga_signals.M_hcounter_d7lto7_0 ));
    InMux I__1609 (
            .O(N__13818),
            .I(N__13815));
    LocalMux I__1608 (
            .O(N__13815),
            .I(N__13812));
    Span4Mux_h I__1607 (
            .O(N__13812),
            .I(N__13807));
    InMux I__1606 (
            .O(N__13811),
            .I(N__13804));
    InMux I__1605 (
            .O(N__13810),
            .I(N__13801));
    Odrv4 I__1604 (
            .O(N__13807),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1603 (
            .O(N__13804),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1602 (
            .O(N__13801),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    CascadeMux I__1601 (
            .O(N__13794),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    InMux I__1600 (
            .O(N__13791),
            .I(N__13788));
    LocalMux I__1599 (
            .O(N__13788),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1 ));
    CascadeMux I__1598 (
            .O(N__13785),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ));
    InMux I__1597 (
            .O(N__13782),
            .I(N__13779));
    LocalMux I__1596 (
            .O(N__13779),
            .I(N__13775));
    InMux I__1595 (
            .O(N__13778),
            .I(N__13772));
    Span4Mux_h I__1594 (
            .O(N__13775),
            .I(N__13765));
    LocalMux I__1593 (
            .O(N__13772),
            .I(N__13762));
    InMux I__1592 (
            .O(N__13771),
            .I(N__13757));
    InMux I__1591 (
            .O(N__13770),
            .I(N__13757));
    InMux I__1590 (
            .O(N__13769),
            .I(N__13752));
    InMux I__1589 (
            .O(N__13768),
            .I(N__13752));
    Odrv4 I__1588 (
            .O(N__13765),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    Odrv4 I__1587 (
            .O(N__13762),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__1586 (
            .O(N__13757),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    LocalMux I__1585 (
            .O(N__13752),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    IoInMux I__1584 (
            .O(N__13743),
            .I(N__13740));
    LocalMux I__1583 (
            .O(N__13740),
            .I(N__13737));
    Span12Mux_s11_v I__1582 (
            .O(N__13737),
            .I(N__13734));
    Span12Mux_h I__1581 (
            .O(N__13734),
            .I(N__13731));
    Odrv12 I__1580 (
            .O(N__13731),
            .I(M_hcounter_q_esr_RNIR18F4_9));
    CascadeMux I__1579 (
            .O(N__13728),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_1_1_cascade_ ));
    InMux I__1578 (
            .O(N__13725),
            .I(N__13719));
    InMux I__1577 (
            .O(N__13724),
            .I(N__13719));
    LocalMux I__1576 (
            .O(N__13719),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1 ));
    InMux I__1575 (
            .O(N__13716),
            .I(N__13713));
    LocalMux I__1574 (
            .O(N__13713),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    InMux I__1573 (
            .O(N__13710),
            .I(N__13707));
    LocalMux I__1572 (
            .O(N__13707),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    CascadeMux I__1571 (
            .O(N__13704),
            .I(\this_vga_signals.mult1_un75_sum_c2_0_cascade_ ));
    InMux I__1570 (
            .O(N__13701),
            .I(N__13698));
    LocalMux I__1569 (
            .O(N__13698),
            .I(\this_vga_signals.if_N_9_1 ));
    InMux I__1568 (
            .O(N__13695),
            .I(N__13690));
    InMux I__1567 (
            .O(N__13694),
            .I(N__13685));
    InMux I__1566 (
            .O(N__13693),
            .I(N__13685));
    LocalMux I__1565 (
            .O(N__13690),
            .I(\this_vga_signals.if_m7_0_x4_0 ));
    LocalMux I__1564 (
            .O(N__13685),
            .I(\this_vga_signals.if_m7_0_x4_0 ));
    InMux I__1563 (
            .O(N__13680),
            .I(N__13676));
    InMux I__1562 (
            .O(N__13679),
            .I(N__13673));
    LocalMux I__1561 (
            .O(N__13676),
            .I(\this_vga_signals.mult1_un75_sum_c3 ));
    LocalMux I__1560 (
            .O(N__13673),
            .I(\this_vga_signals.mult1_un75_sum_c3 ));
    InMux I__1559 (
            .O(N__13668),
            .I(N__13661));
    InMux I__1558 (
            .O(N__13667),
            .I(N__13658));
    InMux I__1557 (
            .O(N__13666),
            .I(N__13651));
    InMux I__1556 (
            .O(N__13665),
            .I(N__13651));
    InMux I__1555 (
            .O(N__13664),
            .I(N__13651));
    LocalMux I__1554 (
            .O(N__13661),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_2 ));
    LocalMux I__1553 (
            .O(N__13658),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_2 ));
    LocalMux I__1552 (
            .O(N__13651),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_2 ));
    CascadeMux I__1551 (
            .O(N__13644),
            .I(\this_vga_signals.mult1_un75_sum_c3_cascade_ ));
    InMux I__1550 (
            .O(N__13641),
            .I(N__13637));
    InMux I__1549 (
            .O(N__13640),
            .I(N__13634));
    LocalMux I__1548 (
            .O(N__13637),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_0 ));
    LocalMux I__1547 (
            .O(N__13634),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_0 ));
    InMux I__1546 (
            .O(N__13629),
            .I(N__13623));
    InMux I__1545 (
            .O(N__13628),
            .I(N__13620));
    InMux I__1544 (
            .O(N__13627),
            .I(N__13615));
    InMux I__1543 (
            .O(N__13626),
            .I(N__13615));
    LocalMux I__1542 (
            .O(N__13623),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1541 (
            .O(N__13620),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1540 (
            .O(N__13615),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    InMux I__1539 (
            .O(N__13608),
            .I(N__13603));
    InMux I__1538 (
            .O(N__13607),
            .I(N__13600));
    InMux I__1537 (
            .O(N__13606),
            .I(N__13597));
    LocalMux I__1536 (
            .O(N__13603),
            .I(\this_vga_signals.N_3_0 ));
    LocalMux I__1535 (
            .O(N__13600),
            .I(\this_vga_signals.N_3_0 ));
    LocalMux I__1534 (
            .O(N__13597),
            .I(\this_vga_signals.N_3_0 ));
    InMux I__1533 (
            .O(N__13590),
            .I(N__13580));
    InMux I__1532 (
            .O(N__13589),
            .I(N__13580));
    InMux I__1531 (
            .O(N__13588),
            .I(N__13580));
    InMux I__1530 (
            .O(N__13587),
            .I(N__13577));
    LocalMux I__1529 (
            .O(N__13580),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    LocalMux I__1528 (
            .O(N__13577),
            .I(\this_vga_signals.M_pcounter_q_i_3_1 ));
    CascadeMux I__1527 (
            .O(N__13572),
            .I(\this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_ ));
    InMux I__1526 (
            .O(N__13569),
            .I(N__13565));
    InMux I__1525 (
            .O(N__13568),
            .I(N__13562));
    LocalMux I__1524 (
            .O(N__13565),
            .I(\this_vga_signals.N_2_0 ));
    LocalMux I__1523 (
            .O(N__13562),
            .I(\this_vga_signals.N_2_0 ));
    InMux I__1522 (
            .O(N__13557),
            .I(N__13553));
    InMux I__1521 (
            .O(N__13556),
            .I(N__13550));
    LocalMux I__1520 (
            .O(N__13553),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    LocalMux I__1519 (
            .O(N__13550),
            .I(\this_vga_signals.M_pcounter_q_i_3_0 ));
    CascadeMux I__1518 (
            .O(N__13545),
            .I(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ));
    CascadeMux I__1517 (
            .O(N__13542),
            .I(\this_vga_signals.M_hcounter_d7_0_cascade_ ));
    InMux I__1516 (
            .O(N__13539),
            .I(N__13536));
    LocalMux I__1515 (
            .O(N__13536),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    CascadeMux I__1514 (
            .O(N__13533),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_x0_cascade_ ));
    CascadeMux I__1513 (
            .O(N__13530),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_ ));
    InMux I__1512 (
            .O(N__13527),
            .I(N__13524));
    LocalMux I__1511 (
            .O(N__13524),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0 ));
    CascadeMux I__1510 (
            .O(N__13521),
            .I(\this_vga_signals.g1_5_cascade_ ));
    InMux I__1509 (
            .O(N__13518),
            .I(N__13515));
    LocalMux I__1508 (
            .O(N__13515),
            .I(\this_vga_signals.g1_0_0 ));
    InMux I__1507 (
            .O(N__13512),
            .I(N__13509));
    LocalMux I__1506 (
            .O(N__13509),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_x1 ));
    InMux I__1505 (
            .O(N__13506),
            .I(N__13503));
    LocalMux I__1504 (
            .O(N__13503),
            .I(\this_vga_signals.g1_2 ));
    InMux I__1503 (
            .O(N__13500),
            .I(N__13489));
    InMux I__1502 (
            .O(N__13499),
            .I(N__13489));
    InMux I__1501 (
            .O(N__13498),
            .I(N__13486));
    InMux I__1500 (
            .O(N__13497),
            .I(N__13483));
    InMux I__1499 (
            .O(N__13496),
            .I(N__13478));
    InMux I__1498 (
            .O(N__13495),
            .I(N__13478));
    InMux I__1497 (
            .O(N__13494),
            .I(N__13475));
    LocalMux I__1496 (
            .O(N__13489),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    LocalMux I__1495 (
            .O(N__13486),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    LocalMux I__1494 (
            .O(N__13483),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    LocalMux I__1493 (
            .O(N__13478),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    LocalMux I__1492 (
            .O(N__13475),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns ));
    CascadeMux I__1491 (
            .O(N__13464),
            .I(\this_vga_signals.mult1_un68_sum_axb1_cascade_ ));
    InMux I__1490 (
            .O(N__13461),
            .I(N__13458));
    LocalMux I__1489 (
            .O(N__13458),
            .I(\this_vga_signals.mult1_un68_sum_c2_0 ));
    CascadeMux I__1488 (
            .O(N__13455),
            .I(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ));
    InMux I__1487 (
            .O(N__13452),
            .I(N__13449));
    LocalMux I__1486 (
            .O(N__13449),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0 ));
    InMux I__1485 (
            .O(N__13446),
            .I(N__13442));
    InMux I__1484 (
            .O(N__13445),
            .I(N__13439));
    LocalMux I__1483 (
            .O(N__13442),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0 ));
    LocalMux I__1482 (
            .O(N__13439),
            .I(\this_vga_signals.mult1_un68_sum_ac0_3_0_0 ));
    InMux I__1481 (
            .O(N__13434),
            .I(N__13430));
    InMux I__1480 (
            .O(N__13433),
            .I(N__13427));
    LocalMux I__1479 (
            .O(N__13430),
            .I(\this_vga_signals.if_i2_mux ));
    LocalMux I__1478 (
            .O(N__13427),
            .I(\this_vga_signals.if_i2_mux ));
    CascadeMux I__1477 (
            .O(N__13422),
            .I(\this_vga_signals.g0_1_1_x0_cascade_ ));
    CascadeMux I__1476 (
            .O(N__13419),
            .I(\this_vga_signals.g0_1_1_cascade_ ));
    InMux I__1475 (
            .O(N__13416),
            .I(N__13413));
    LocalMux I__1474 (
            .O(N__13413),
            .I(\this_vga_signals.N_4_0_0_0 ));
    CascadeMux I__1473 (
            .O(N__13410),
            .I(\this_vga_signals.g0_0_0_0_0_cascade_ ));
    InMux I__1472 (
            .O(N__13407),
            .I(N__13398));
    InMux I__1471 (
            .O(N__13406),
            .I(N__13398));
    InMux I__1470 (
            .O(N__13405),
            .I(N__13393));
    InMux I__1469 (
            .O(N__13404),
            .I(N__13393));
    InMux I__1468 (
            .O(N__13403),
            .I(N__13390));
    LocalMux I__1467 (
            .O(N__13398),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1466 (
            .O(N__13393),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1465 (
            .O(N__13390),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    InMux I__1464 (
            .O(N__13383),
            .I(N__13375));
    InMux I__1463 (
            .O(N__13382),
            .I(N__13375));
    InMux I__1462 (
            .O(N__13381),
            .I(N__13370));
    InMux I__1461 (
            .O(N__13380),
            .I(N__13370));
    LocalMux I__1460 (
            .O(N__13375),
            .I(N__13367));
    LocalMux I__1459 (
            .O(N__13370),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    Odrv4 I__1458 (
            .O(N__13367),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    CascadeMux I__1457 (
            .O(N__13362),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ));
    InMux I__1456 (
            .O(N__13359),
            .I(N__13356));
    LocalMux I__1455 (
            .O(N__13356),
            .I(N__13351));
    InMux I__1454 (
            .O(N__13355),
            .I(N__13346));
    InMux I__1453 (
            .O(N__13354),
            .I(N__13346));
    Span4Mux_v I__1452 (
            .O(N__13351),
            .I(N__13343));
    LocalMux I__1451 (
            .O(N__13346),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    Odrv4 I__1450 (
            .O(N__13343),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    CascadeMux I__1449 (
            .O(N__13338),
            .I(N__13335));
    InMux I__1448 (
            .O(N__13335),
            .I(N__13332));
    LocalMux I__1447 (
            .O(N__13332),
            .I(N__13329));
    Odrv4 I__1446 (
            .O(N__13329),
            .I(\this_vga_signals.g0_0_0_1 ));
    InMux I__1445 (
            .O(N__13326),
            .I(N__13323));
    LocalMux I__1444 (
            .O(N__13323),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i_0 ));
    CascadeMux I__1443 (
            .O(N__13320),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_cascade_ ));
    CascadeMux I__1442 (
            .O(N__13317),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_cascade_ ));
    InMux I__1441 (
            .O(N__13314),
            .I(N__13311));
    LocalMux I__1440 (
            .O(N__13311),
            .I(N__13308));
    Odrv12 I__1439 (
            .O(N__13308),
            .I(M_this_map_ram_write_data_0));
    InMux I__1438 (
            .O(N__13305),
            .I(N__13302));
    LocalMux I__1437 (
            .O(N__13302),
            .I(N__13299));
    Span4Mux_h I__1436 (
            .O(N__13299),
            .I(N__13296));
    Span4Mux_h I__1435 (
            .O(N__13296),
            .I(N__13293));
    Odrv4 I__1434 (
            .O(N__13293),
            .I(M_this_map_ram_write_data_7));
    InMux I__1433 (
            .O(N__13290),
            .I(N__13287));
    LocalMux I__1432 (
            .O(N__13287),
            .I(N__13284));
    Span4Mux_v I__1431 (
            .O(N__13284),
            .I(N__13281));
    Odrv4 I__1430 (
            .O(N__13281),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    InMux I__1429 (
            .O(N__13278),
            .I(N__13275));
    LocalMux I__1428 (
            .O(N__13275),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__1427 (
            .O(N__13272),
            .I(\this_vga_signals.N_1_4_1_cascade_ ));
    CascadeMux I__1426 (
            .O(N__13269),
            .I(\this_vga_signals.SUM_2_i_1_2_3_cascade_ ));
    InMux I__1425 (
            .O(N__13266),
            .I(N__13263));
    LocalMux I__1424 (
            .O(N__13263),
            .I(N__13255));
    InMux I__1423 (
            .O(N__13262),
            .I(N__13250));
    InMux I__1422 (
            .O(N__13261),
            .I(N__13250));
    InMux I__1421 (
            .O(N__13260),
            .I(N__13243));
    InMux I__1420 (
            .O(N__13259),
            .I(N__13243));
    InMux I__1419 (
            .O(N__13258),
            .I(N__13243));
    Odrv4 I__1418 (
            .O(N__13255),
            .I(N_880_0));
    LocalMux I__1417 (
            .O(N__13250),
            .I(N_880_0));
    LocalMux I__1416 (
            .O(N__13243),
            .I(N_880_0));
    CascadeMux I__1415 (
            .O(N__13236),
            .I(N__13233));
    InMux I__1414 (
            .O(N__13233),
            .I(N__13230));
    LocalMux I__1413 (
            .O(N__13230),
            .I(N__13227));
    Span4Mux_h I__1412 (
            .O(N__13227),
            .I(N__13224));
    Span4Mux_h I__1411 (
            .O(N__13224),
            .I(N__13221));
    Odrv4 I__1410 (
            .O(N__13221),
            .I(M_this_vga_signals_address_2));
    InMux I__1409 (
            .O(N__13218),
            .I(N__13215));
    LocalMux I__1408 (
            .O(N__13215),
            .I(\this_vga_signals.mult1_un82_sum_c2_0 ));
    CascadeMux I__1407 (
            .O(N__13212),
            .I(\this_vga_signals.mult1_un82_sum_c2_0_cascade_ ));
    InMux I__1406 (
            .O(N__13209),
            .I(N__13203));
    InMux I__1405 (
            .O(N__13208),
            .I(N__13203));
    LocalMux I__1404 (
            .O(N__13203),
            .I(\this_vga_signals.mult1_un82_sum_c3_0 ));
    CascadeMux I__1403 (
            .O(N__13200),
            .I(N__13197));
    InMux I__1402 (
            .O(N__13197),
            .I(N__13193));
    InMux I__1401 (
            .O(N__13196),
            .I(N__13190));
    LocalMux I__1400 (
            .O(N__13193),
            .I(\this_vga_signals.mult1_un75_sum_axbxc1 ));
    LocalMux I__1399 (
            .O(N__13190),
            .I(\this_vga_signals.mult1_un75_sum_axbxc1 ));
    CascadeMux I__1398 (
            .O(N__13185),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_2_0_cascade_ ));
    CascadeMux I__1397 (
            .O(N__13182),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_0_2_cascade_ ));
    InMux I__1396 (
            .O(N__13179),
            .I(N__13175));
    InMux I__1395 (
            .O(N__13178),
            .I(N__13172));
    LocalMux I__1394 (
            .O(N__13175),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1 ));
    LocalMux I__1393 (
            .O(N__13172),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1 ));
    InMux I__1392 (
            .O(N__13167),
            .I(N__13164));
    LocalMux I__1391 (
            .O(N__13164),
            .I(N__13161));
    Span12Mux_v I__1390 (
            .O(N__13161),
            .I(N__13158));
    Span12Mux_v I__1389 (
            .O(N__13158),
            .I(N__13155));
    Span12Mux_h I__1388 (
            .O(N__13155),
            .I(N__13152));
    Odrv12 I__1387 (
            .O(N__13152),
            .I(M_this_oam_ram_read_data_4));
    InMux I__1386 (
            .O(N__13149),
            .I(N__13146));
    LocalMux I__1385 (
            .O(N__13146),
            .I(N__13143));
    Span4Mux_v I__1384 (
            .O(N__13143),
            .I(N__13140));
    Span4Mux_v I__1383 (
            .O(N__13140),
            .I(N__13137));
    Span4Mux_h I__1382 (
            .O(N__13137),
            .I(N__13134));
    Odrv4 I__1381 (
            .O(N__13134),
            .I(M_this_map_ram_read_data_4));
    CascadeMux I__1380 (
            .O(N__13131),
            .I(N__13128));
    InMux I__1379 (
            .O(N__13128),
            .I(N__13122));
    CascadeMux I__1378 (
            .O(N__13127),
            .I(N__13119));
    CascadeMux I__1377 (
            .O(N__13126),
            .I(N__13114));
    CascadeMux I__1376 (
            .O(N__13125),
            .I(N__13108));
    LocalMux I__1375 (
            .O(N__13122),
            .I(N__13102));
    InMux I__1374 (
            .O(N__13119),
            .I(N__13099));
    CascadeMux I__1373 (
            .O(N__13118),
            .I(N__13096));
    CascadeMux I__1372 (
            .O(N__13117),
            .I(N__13093));
    InMux I__1371 (
            .O(N__13114),
            .I(N__13090));
    CascadeMux I__1370 (
            .O(N__13113),
            .I(N__13087));
    CascadeMux I__1369 (
            .O(N__13112),
            .I(N__13083));
    CascadeMux I__1368 (
            .O(N__13111),
            .I(N__13078));
    InMux I__1367 (
            .O(N__13108),
            .I(N__13075));
    CascadeMux I__1366 (
            .O(N__13107),
            .I(N__13072));
    CascadeMux I__1365 (
            .O(N__13106),
            .I(N__13069));
    CascadeMux I__1364 (
            .O(N__13105),
            .I(N__13066));
    Span4Mux_s3_v I__1363 (
            .O(N__13102),
            .I(N__13061));
    LocalMux I__1362 (
            .O(N__13099),
            .I(N__13061));
    InMux I__1361 (
            .O(N__13096),
            .I(N__13058));
    InMux I__1360 (
            .O(N__13093),
            .I(N__13055));
    LocalMux I__1359 (
            .O(N__13090),
            .I(N__13052));
    InMux I__1358 (
            .O(N__13087),
            .I(N__13049));
    CascadeMux I__1357 (
            .O(N__13086),
            .I(N__13046));
    InMux I__1356 (
            .O(N__13083),
            .I(N__13043));
    CascadeMux I__1355 (
            .O(N__13082),
            .I(N__13040));
    CascadeMux I__1354 (
            .O(N__13081),
            .I(N__13037));
    InMux I__1353 (
            .O(N__13078),
            .I(N__13033));
    LocalMux I__1352 (
            .O(N__13075),
            .I(N__13030));
    InMux I__1351 (
            .O(N__13072),
            .I(N__13027));
    InMux I__1350 (
            .O(N__13069),
            .I(N__13024));
    InMux I__1349 (
            .O(N__13066),
            .I(N__13021));
    Span4Mux_v I__1348 (
            .O(N__13061),
            .I(N__13014));
    LocalMux I__1347 (
            .O(N__13058),
            .I(N__13014));
    LocalMux I__1346 (
            .O(N__13055),
            .I(N__13014));
    Span4Mux_h I__1345 (
            .O(N__13052),
            .I(N__13009));
    LocalMux I__1344 (
            .O(N__13049),
            .I(N__13009));
    InMux I__1343 (
            .O(N__13046),
            .I(N__13006));
    LocalMux I__1342 (
            .O(N__13043),
            .I(N__13003));
    InMux I__1341 (
            .O(N__13040),
            .I(N__13000));
    InMux I__1340 (
            .O(N__13037),
            .I(N__12997));
    CascadeMux I__1339 (
            .O(N__13036),
            .I(N__12994));
    LocalMux I__1338 (
            .O(N__13033),
            .I(N__12991));
    Span4Mux_v I__1337 (
            .O(N__13030),
            .I(N__12988));
    LocalMux I__1336 (
            .O(N__13027),
            .I(N__12985));
    LocalMux I__1335 (
            .O(N__13024),
            .I(N__12982));
    LocalMux I__1334 (
            .O(N__13021),
            .I(N__12979));
    Span4Mux_v I__1333 (
            .O(N__13014),
            .I(N__12972));
    Span4Mux_v I__1332 (
            .O(N__13009),
            .I(N__12972));
    LocalMux I__1331 (
            .O(N__13006),
            .I(N__12972));
    Span4Mux_v I__1330 (
            .O(N__13003),
            .I(N__12967));
    LocalMux I__1329 (
            .O(N__13000),
            .I(N__12967));
    LocalMux I__1328 (
            .O(N__12997),
            .I(N__12964));
    InMux I__1327 (
            .O(N__12994),
            .I(N__12961));
    Span12Mux_h I__1326 (
            .O(N__12991),
            .I(N__12958));
    Sp12to4 I__1325 (
            .O(N__12988),
            .I(N__12953));
    Span12Mux_v I__1324 (
            .O(N__12985),
            .I(N__12953));
    Span12Mux_s6_v I__1323 (
            .O(N__12982),
            .I(N__12948));
    Span12Mux_v I__1322 (
            .O(N__12979),
            .I(N__12948));
    Span4Mux_h I__1321 (
            .O(N__12972),
            .I(N__12945));
    Span4Mux_v I__1320 (
            .O(N__12967),
            .I(N__12940));
    Span4Mux_h I__1319 (
            .O(N__12964),
            .I(N__12940));
    LocalMux I__1318 (
            .O(N__12961),
            .I(N__12937));
    Span12Mux_v I__1317 (
            .O(N__12958),
            .I(N__12934));
    Span12Mux_h I__1316 (
            .O(N__12953),
            .I(N__12929));
    Span12Mux_h I__1315 (
            .O(N__12948),
            .I(N__12929));
    Sp12to4 I__1314 (
            .O(N__12945),
            .I(N__12926));
    Span4Mux_h I__1313 (
            .O(N__12940),
            .I(N__12923));
    Span4Mux_h I__1312 (
            .O(N__12937),
            .I(N__12920));
    Odrv12 I__1311 (
            .O(N__12934),
            .I(M_this_ppu_sprites_addr_10));
    Odrv12 I__1310 (
            .O(N__12929),
            .I(M_this_ppu_sprites_addr_10));
    Odrv12 I__1309 (
            .O(N__12926),
            .I(M_this_ppu_sprites_addr_10));
    Odrv4 I__1308 (
            .O(N__12923),
            .I(M_this_ppu_sprites_addr_10));
    Odrv4 I__1307 (
            .O(N__12920),
            .I(M_this_ppu_sprites_addr_10));
    CascadeMux I__1306 (
            .O(N__12909),
            .I(\this_vga_signals.M_vcounter_d7lt3_cascade_ ));
    InMux I__1305 (
            .O(N__12906),
            .I(N__12903));
    LocalMux I__1304 (
            .O(N__12903),
            .I(\this_vga_ramdac.N_24_mux ));
    InMux I__1303 (
            .O(N__12900),
            .I(N__12897));
    LocalMux I__1302 (
            .O(N__12897),
            .I(N__12888));
    InMux I__1301 (
            .O(N__12896),
            .I(N__12885));
    InMux I__1300 (
            .O(N__12895),
            .I(N__12880));
    InMux I__1299 (
            .O(N__12894),
            .I(N__12880));
    InMux I__1298 (
            .O(N__12893),
            .I(N__12877));
    InMux I__1297 (
            .O(N__12892),
            .I(N__12872));
    InMux I__1296 (
            .O(N__12891),
            .I(N__12872));
    Odrv4 I__1295 (
            .O(N__12888),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    LocalMux I__1294 (
            .O(N__12885),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    LocalMux I__1293 (
            .O(N__12880),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    LocalMux I__1292 (
            .O(N__12877),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    LocalMux I__1291 (
            .O(N__12872),
            .I(M_pcounter_q_ret_2_RNIH7PG8));
    InMux I__1290 (
            .O(N__12861),
            .I(N__12857));
    CascadeMux I__1289 (
            .O(N__12860),
            .I(N__12854));
    LocalMux I__1288 (
            .O(N__12857),
            .I(N__12851));
    InMux I__1287 (
            .O(N__12854),
            .I(N__12848));
    Odrv4 I__1286 (
            .O(N__12851),
            .I(\this_vga_ramdac.N_3298_reto ));
    LocalMux I__1285 (
            .O(N__12848),
            .I(\this_vga_ramdac.N_3298_reto ));
    CascadeMux I__1284 (
            .O(N__12843),
            .I(\this_vga_signals.M_pcounter_q_3_1_cascade_ ));
    CascadeMux I__1283 (
            .O(N__12840),
            .I(N__12836));
    CascadeMux I__1282 (
            .O(N__12839),
            .I(N__12832));
    InMux I__1281 (
            .O(N__12836),
            .I(N__12825));
    InMux I__1280 (
            .O(N__12835),
            .I(N__12825));
    InMux I__1279 (
            .O(N__12832),
            .I(N__12825));
    LocalMux I__1278 (
            .O(N__12825),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    InMux I__1277 (
            .O(N__12822),
            .I(N__12817));
    InMux I__1276 (
            .O(N__12821),
            .I(N__12812));
    InMux I__1275 (
            .O(N__12820),
            .I(N__12812));
    LocalMux I__1274 (
            .O(N__12817),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__1273 (
            .O(N__12812),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    CascadeMux I__1272 (
            .O(N__12807),
            .I(N__12804));
    InMux I__1271 (
            .O(N__12804),
            .I(N__12801));
    LocalMux I__1270 (
            .O(N__12801),
            .I(N__12798));
    Span4Mux_h I__1269 (
            .O(N__12798),
            .I(N__12795));
    Span4Mux_h I__1268 (
            .O(N__12795),
            .I(N__12792));
    Odrv4 I__1267 (
            .O(N__12792),
            .I(M_this_vga_signals_address_1));
    CascadeMux I__1266 (
            .O(N__12789),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_1_cascade_ ));
    CascadeMux I__1265 (
            .O(N__12786),
            .I(N__12783));
    InMux I__1264 (
            .O(N__12783),
            .I(N__12780));
    LocalMux I__1263 (
            .O(N__12780),
            .I(N__12777));
    Span12Mux_h I__1262 (
            .O(N__12777),
            .I(N__12774));
    Odrv12 I__1261 (
            .O(N__12774),
            .I(M_this_vga_signals_address_0));
    CascadeMux I__1260 (
            .O(N__12771),
            .I(\this_vga_signals.g0_2_1_cascade_ ));
    InMux I__1259 (
            .O(N__12768),
            .I(N__12765));
    LocalMux I__1258 (
            .O(N__12765),
            .I(\this_vga_signals.N_5_0_0 ));
    InMux I__1257 (
            .O(N__12762),
            .I(N__12759));
    LocalMux I__1256 (
            .O(N__12759),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_x1 ));
    InMux I__1255 (
            .O(N__12756),
            .I(N__12753));
    LocalMux I__1254 (
            .O(N__12753),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_x0 ));
    CascadeMux I__1253 (
            .O(N__12750),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_ns_cascade_ ));
    InMux I__1252 (
            .O(N__12747),
            .I(N__12744));
    LocalMux I__1251 (
            .O(N__12744),
            .I(\this_vga_signals.g0_31_N_4L6 ));
    CascadeMux I__1250 (
            .O(N__12741),
            .I(\this_vga_signals.g0_31_N_2L1_cascade_ ));
    InMux I__1249 (
            .O(N__12738),
            .I(N__12735));
    LocalMux I__1248 (
            .O(N__12735),
            .I(\this_vga_signals.g0_31_N_5L8 ));
    CascadeMux I__1247 (
            .O(N__12732),
            .I(\this_vga_signals.M_pcounter_q_3_0_cascade_ ));
    CascadeMux I__1246 (
            .O(N__12729),
            .I(\this_vga_signals.N_2_0_cascade_ ));
    InMux I__1245 (
            .O(N__12726),
            .I(N__12723));
    LocalMux I__1244 (
            .O(N__12723),
            .I(\this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ));
    InMux I__1243 (
            .O(N__12720),
            .I(N__12715));
    InMux I__1242 (
            .O(N__12719),
            .I(N__12712));
    InMux I__1241 (
            .O(N__12718),
            .I(N__12709));
    LocalMux I__1240 (
            .O(N__12715),
            .I(N__12704));
    LocalMux I__1239 (
            .O(N__12712),
            .I(N__12704));
    LocalMux I__1238 (
            .O(N__12709),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv12 I__1237 (
            .O(N__12704),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__1236 (
            .O(N__12699),
            .I(\this_vga_signals.if_i1_mux_0_cascade_ ));
    CascadeMux I__1235 (
            .O(N__12696),
            .I(N__12693));
    InMux I__1234 (
            .O(N__12693),
            .I(N__12690));
    LocalMux I__1233 (
            .O(N__12690),
            .I(N__12687));
    Span4Mux_h I__1232 (
            .O(N__12687),
            .I(N__12684));
    Span4Mux_h I__1231 (
            .O(N__12684),
            .I(N__12681));
    Odrv4 I__1230 (
            .O(N__12681),
            .I(M_this_vga_signals_address_7));
    CascadeMux I__1229 (
            .O(N__12678),
            .I(\this_vga_signals.N_5_i_0_cascade_ ));
    InMux I__1228 (
            .O(N__12675),
            .I(N__12672));
    LocalMux I__1227 (
            .O(N__12672),
            .I(\this_vga_signals.mult1_un82_sum_c3 ));
    InMux I__1226 (
            .O(N__12669),
            .I(N__12666));
    LocalMux I__1225 (
            .O(N__12666),
            .I(\this_vga_signals.N_3_2_0_1 ));
    CascadeMux I__1224 (
            .O(N__12663),
            .I(\this_vga_signals.g0_i_x4_0_0_cascade_ ));
    InMux I__1223 (
            .O(N__12660),
            .I(N__12657));
    LocalMux I__1222 (
            .O(N__12657),
            .I(\this_vga_signals.N_3_3_0_0 ));
    CascadeMux I__1221 (
            .O(N__12654),
            .I(\this_vga_signals.g0_0_2_0_0_cascade_ ));
    InMux I__1220 (
            .O(N__12651),
            .I(N__12648));
    LocalMux I__1219 (
            .O(N__12648),
            .I(\this_vga_signals.g0_6_2 ));
    CascadeMux I__1218 (
            .O(N__12645),
            .I(\this_vga_signals.g1_1_0_0_0_cascade_ ));
    InMux I__1217 (
            .O(N__12642),
            .I(N__12639));
    LocalMux I__1216 (
            .O(N__12639),
            .I(\this_vga_signals.N_5_i_1_0_0 ));
    InMux I__1215 (
            .O(N__12636),
            .I(N__12633));
    LocalMux I__1214 (
            .O(N__12633),
            .I(N__12628));
    InMux I__1213 (
            .O(N__12632),
            .I(N__12623));
    InMux I__1212 (
            .O(N__12631),
            .I(N__12623));
    Odrv4 I__1211 (
            .O(N__12628),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__1210 (
            .O(N__12623),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    InMux I__1209 (
            .O(N__12618),
            .I(N__12615));
    LocalMux I__1208 (
            .O(N__12615),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    CascadeMux I__1207 (
            .O(N__12612),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ));
    CascadeMux I__1206 (
            .O(N__12609),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ));
    CascadeMux I__1205 (
            .O(N__12606),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    InMux I__1204 (
            .O(N__12603),
            .I(N__12600));
    LocalMux I__1203 (
            .O(N__12600),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_0 ));
    InMux I__1202 (
            .O(N__12597),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__1201 (
            .O(N__12594),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__1200 (
            .O(N__12591),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__1199 (
            .O(N__12588),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__1198 (
            .O(N__12585),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__1197 (
            .O(N__12582),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__1196 (
            .O(N__12579),
            .I(bfn_13_13_0_));
    InMux I__1195 (
            .O(N__12576),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    CascadeMux I__1194 (
            .O(N__12573),
            .I(N_880_0_cascade_));
    CascadeMux I__1193 (
            .O(N__12570),
            .I(N__12567));
    InMux I__1192 (
            .O(N__12567),
            .I(N__12564));
    LocalMux I__1191 (
            .O(N__12564),
            .I(N__12561));
    Span4Mux_v I__1190 (
            .O(N__12561),
            .I(N__12558));
    Odrv4 I__1189 (
            .O(N__12558),
            .I(M_this_vga_signals_address_5));
    CascadeMux I__1188 (
            .O(N__12555),
            .I(N__12552));
    InMux I__1187 (
            .O(N__12552),
            .I(N__12549));
    LocalMux I__1186 (
            .O(N__12549),
            .I(N__12546));
    Span4Mux_h I__1185 (
            .O(N__12546),
            .I(N__12543));
    Odrv4 I__1184 (
            .O(N__12543),
            .I(M_this_vga_signals_address_3));
    CascadeMux I__1183 (
            .O(N__12540),
            .I(N__12537));
    InMux I__1182 (
            .O(N__12537),
            .I(N__12534));
    LocalMux I__1181 (
            .O(N__12534),
            .I(N__12531));
    Span4Mux_h I__1180 (
            .O(N__12531),
            .I(N__12528));
    Odrv4 I__1179 (
            .O(N__12528),
            .I(M_this_vga_signals_address_4));
    InMux I__1178 (
            .O(N__12525),
            .I(N__12522));
    LocalMux I__1177 (
            .O(N__12522),
            .I(N__12519));
    Span12Mux_h I__1176 (
            .O(N__12519),
            .I(N__12516));
    Odrv12 I__1175 (
            .O(N__12516),
            .I(port_clk_c));
    InMux I__1174 (
            .O(N__12513),
            .I(N__12510));
    LocalMux I__1173 (
            .O(N__12510),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    InMux I__1172 (
            .O(N__12507),
            .I(N__12504));
    LocalMux I__1171 (
            .O(N__12504),
            .I(N__12501));
    Span4Mux_h I__1170 (
            .O(N__12501),
            .I(N__12498));
    Odrv4 I__1169 (
            .O(N__12498),
            .I(M_this_map_ram_write_data_1));
    InMux I__1168 (
            .O(N__12495),
            .I(N__12492));
    LocalMux I__1167 (
            .O(N__12492),
            .I(N__12489));
    Span4Mux_h I__1166 (
            .O(N__12489),
            .I(N__12486));
    Odrv4 I__1165 (
            .O(N__12486),
            .I(M_this_map_ram_write_data_5));
    InMux I__1164 (
            .O(N__12483),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    CascadeMux I__1163 (
            .O(N__12480),
            .I(\this_vga_ramdac.m19_cascade_ ));
    InMux I__1162 (
            .O(N__12477),
            .I(N__12474));
    LocalMux I__1161 (
            .O(N__12474),
            .I(N__12471));
    Span4Mux_h I__1160 (
            .O(N__12471),
            .I(N__12468));
    Sp12to4 I__1159 (
            .O(N__12468),
            .I(N__12464));
    InMux I__1158 (
            .O(N__12467),
            .I(N__12461));
    Odrv12 I__1157 (
            .O(N__12464),
            .I(\this_vga_ramdac.N_3302_reto ));
    LocalMux I__1156 (
            .O(N__12461),
            .I(\this_vga_ramdac.N_3302_reto ));
    InMux I__1155 (
            .O(N__12456),
            .I(N__12453));
    LocalMux I__1154 (
            .O(N__12453),
            .I(N__12449));
    InMux I__1153 (
            .O(N__12452),
            .I(N__12446));
    Odrv4 I__1152 (
            .O(N__12449),
            .I(\this_vga_ramdac.N_3303_reto ));
    LocalMux I__1151 (
            .O(N__12446),
            .I(\this_vga_ramdac.N_3303_reto ));
    CascadeMux I__1150 (
            .O(N__12441),
            .I(N__12437));
    CascadeMux I__1149 (
            .O(N__12440),
            .I(N__12434));
    InMux I__1148 (
            .O(N__12437),
            .I(N__12425));
    InMux I__1147 (
            .O(N__12434),
            .I(N__12425));
    InMux I__1146 (
            .O(N__12433),
            .I(N__12416));
    InMux I__1145 (
            .O(N__12432),
            .I(N__12416));
    InMux I__1144 (
            .O(N__12431),
            .I(N__12416));
    InMux I__1143 (
            .O(N__12430),
            .I(N__12416));
    LocalMux I__1142 (
            .O(N__12425),
            .I(N__12411));
    LocalMux I__1141 (
            .O(N__12416),
            .I(N__12411));
    Span4Mux_h I__1140 (
            .O(N__12411),
            .I(N__12408));
    Odrv4 I__1139 (
            .O(N__12408),
            .I(M_this_vram_read_data_0));
    CascadeMux I__1138 (
            .O(N__12405),
            .I(N__12400));
    InMux I__1137 (
            .O(N__12404),
            .I(N__12392));
    InMux I__1136 (
            .O(N__12403),
            .I(N__12392));
    InMux I__1135 (
            .O(N__12400),
            .I(N__12383));
    InMux I__1134 (
            .O(N__12399),
            .I(N__12383));
    InMux I__1133 (
            .O(N__12398),
            .I(N__12383));
    InMux I__1132 (
            .O(N__12397),
            .I(N__12383));
    LocalMux I__1131 (
            .O(N__12392),
            .I(N__12378));
    LocalMux I__1130 (
            .O(N__12383),
            .I(N__12378));
    Span4Mux_h I__1129 (
            .O(N__12378),
            .I(N__12375));
    Odrv4 I__1128 (
            .O(N__12375),
            .I(M_this_vram_read_data_3));
    CascadeMux I__1127 (
            .O(N__12372),
            .I(N__12365));
    CascadeMux I__1126 (
            .O(N__12371),
            .I(N__12362));
    InMux I__1125 (
            .O(N__12370),
            .I(N__12357));
    InMux I__1124 (
            .O(N__12369),
            .I(N__12357));
    InMux I__1123 (
            .O(N__12368),
            .I(N__12350));
    InMux I__1122 (
            .O(N__12365),
            .I(N__12350));
    InMux I__1121 (
            .O(N__12362),
            .I(N__12350));
    LocalMux I__1120 (
            .O(N__12357),
            .I(N__12345));
    LocalMux I__1119 (
            .O(N__12350),
            .I(N__12345));
    Span4Mux_h I__1118 (
            .O(N__12345),
            .I(N__12342));
    Odrv4 I__1117 (
            .O(N__12342),
            .I(M_this_vram_read_data_2));
    InMux I__1116 (
            .O(N__12339),
            .I(N__12329));
    InMux I__1115 (
            .O(N__12338),
            .I(N__12329));
    InMux I__1114 (
            .O(N__12337),
            .I(N__12320));
    InMux I__1113 (
            .O(N__12336),
            .I(N__12320));
    InMux I__1112 (
            .O(N__12335),
            .I(N__12320));
    InMux I__1111 (
            .O(N__12334),
            .I(N__12320));
    LocalMux I__1110 (
            .O(N__12329),
            .I(N__12315));
    LocalMux I__1109 (
            .O(N__12320),
            .I(N__12315));
    Span4Mux_h I__1108 (
            .O(N__12315),
            .I(N__12312));
    Odrv4 I__1107 (
            .O(N__12312),
            .I(M_this_vram_read_data_1));
    InMux I__1106 (
            .O(N__12309),
            .I(N__12306));
    LocalMux I__1105 (
            .O(N__12306),
            .I(\this_vga_ramdac.i2_mux_0 ));
    InMux I__1104 (
            .O(N__12303),
            .I(N__12297));
    InMux I__1103 (
            .O(N__12302),
            .I(N__12297));
    LocalMux I__1102 (
            .O(N__12297),
            .I(this_pixel_clk_M_counter_q_i_1));
    InMux I__1101 (
            .O(N__12294),
            .I(N__12289));
    InMux I__1100 (
            .O(N__12293),
            .I(N__12286));
    InMux I__1099 (
            .O(N__12292),
            .I(N__12283));
    LocalMux I__1098 (
            .O(N__12289),
            .I(this_pixel_clk_M_counter_q_0));
    LocalMux I__1097 (
            .O(N__12286),
            .I(this_pixel_clk_M_counter_q_0));
    LocalMux I__1096 (
            .O(N__12283),
            .I(this_pixel_clk_M_counter_q_0));
    InMux I__1095 (
            .O(N__12276),
            .I(N__12272));
    InMux I__1094 (
            .O(N__12275),
            .I(N__12269));
    LocalMux I__1093 (
            .O(N__12272),
            .I(N__12263));
    LocalMux I__1092 (
            .O(N__12269),
            .I(N__12263));
    InMux I__1091 (
            .O(N__12268),
            .I(N__12259));
    Span4Mux_v I__1090 (
            .O(N__12263),
            .I(N__12254));
    InMux I__1089 (
            .O(N__12262),
            .I(N__12251));
    LocalMux I__1088 (
            .O(N__12259),
            .I(N__12248));
    InMux I__1087 (
            .O(N__12258),
            .I(N__12245));
    CascadeMux I__1086 (
            .O(N__12257),
            .I(N__12241));
    Span4Mux_h I__1085 (
            .O(N__12254),
            .I(N__12236));
    LocalMux I__1084 (
            .O(N__12251),
            .I(N__12236));
    Span4Mux_h I__1083 (
            .O(N__12248),
            .I(N__12231));
    LocalMux I__1082 (
            .O(N__12245),
            .I(N__12231));
    InMux I__1081 (
            .O(N__12244),
            .I(N__12228));
    InMux I__1080 (
            .O(N__12241),
            .I(N__12225));
    Odrv4 I__1079 (
            .O(N__12236),
            .I(\this_vga_ramdac.N_880_i_reto ));
    Odrv4 I__1078 (
            .O(N__12231),
            .I(\this_vga_ramdac.N_880_i_reto ));
    LocalMux I__1077 (
            .O(N__12228),
            .I(\this_vga_ramdac.N_880_i_reto ));
    LocalMux I__1076 (
            .O(N__12225),
            .I(\this_vga_ramdac.N_880_i_reto ));
    InMux I__1075 (
            .O(N__12216),
            .I(N__12213));
    LocalMux I__1074 (
            .O(N__12213),
            .I(\this_vga_signals.if_m8_0_a3_1_1_1 ));
    CascadeMux I__1073 (
            .O(N__12210),
            .I(\this_vga_signals.if_N_5_cascade_ ));
    CascadeMux I__1072 (
            .O(N__12207),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ));
    InMux I__1071 (
            .O(N__12204),
            .I(N__12201));
    LocalMux I__1070 (
            .O(N__12201),
            .I(N__12198));
    Odrv4 I__1069 (
            .O(N__12198),
            .I(\this_vga_signals.mult1_un47_sum_c3_1_1_0 ));
    InMux I__1068 (
            .O(N__12195),
            .I(N__12192));
    LocalMux I__1067 (
            .O(N__12192),
            .I(N__12188));
    CascadeMux I__1066 (
            .O(N__12191),
            .I(N__12185));
    Span4Mux_v I__1065 (
            .O(N__12188),
            .I(N__12182));
    InMux I__1064 (
            .O(N__12185),
            .I(N__12179));
    Odrv4 I__1063 (
            .O(N__12182),
            .I(\this_vga_ramdac.N_3301_reto ));
    LocalMux I__1062 (
            .O(N__12179),
            .I(\this_vga_ramdac.N_3301_reto ));
    CascadeMux I__1061 (
            .O(N__12174),
            .I(\this_vga_signals.vvisibility_1_cascade_ ));
    InMux I__1060 (
            .O(N__12171),
            .I(N__12168));
    LocalMux I__1059 (
            .O(N__12168),
            .I(\this_vga_ramdac.m16 ));
    CascadeMux I__1058 (
            .O(N__12165),
            .I(N__12162));
    InMux I__1057 (
            .O(N__12162),
            .I(N__12159));
    LocalMux I__1056 (
            .O(N__12159),
            .I(\this_vga_signals.vaddress_5_0_6 ));
    InMux I__1055 (
            .O(N__12156),
            .I(N__12153));
    LocalMux I__1054 (
            .O(N__12153),
            .I(\this_vga_signals.N_5 ));
    InMux I__1053 (
            .O(N__12150),
            .I(N__12147));
    LocalMux I__1052 (
            .O(N__12147),
            .I(\this_vga_signals.if_m8_0_a3_1_1_0 ));
    CascadeMux I__1051 (
            .O(N__12144),
            .I(N__12141));
    InMux I__1050 (
            .O(N__12141),
            .I(N__12138));
    LocalMux I__1049 (
            .O(N__12138),
            .I(\this_vga_signals.g2_5 ));
    InMux I__1048 (
            .O(N__12135),
            .I(N__12132));
    LocalMux I__1047 (
            .O(N__12132),
            .I(\this_vga_signals.N_18_0 ));
    CascadeMux I__1046 (
            .O(N__12129),
            .I(\this_vga_signals.g0_7_0_cascade_ ));
    InMux I__1045 (
            .O(N__12126),
            .I(N__12123));
    LocalMux I__1044 (
            .O(N__12123),
            .I(N__12120));
    Odrv4 I__1043 (
            .O(N__12120),
            .I(\this_vga_signals.g1_0_0_0 ));
    CascadeMux I__1042 (
            .O(N__12117),
            .I(\this_vga_signals.N_4_0_0_cascade_ ));
    IoInMux I__1041 (
            .O(N__12114),
            .I(N__12111));
    LocalMux I__1040 (
            .O(N__12111),
            .I(N__12108));
    IoSpan4Mux I__1039 (
            .O(N__12108),
            .I(N__12105));
    Span4Mux_s3_v I__1038 (
            .O(N__12105),
            .I(N__12102));
    Span4Mux_h I__1037 (
            .O(N__12102),
            .I(N__12099));
    Sp12to4 I__1036 (
            .O(N__12099),
            .I(N__12096));
    Odrv12 I__1035 (
            .O(N__12096),
            .I(N_495));
    CascadeMux I__1034 (
            .O(N__12093),
            .I(\this_vga_signals.un2_vsynclt8_cascade_ ));
    IoInMux I__1033 (
            .O(N__12090),
            .I(N__12087));
    LocalMux I__1032 (
            .O(N__12087),
            .I(N__12084));
    Span4Mux_s2_v I__1031 (
            .O(N__12084),
            .I(N__12081));
    Span4Mux_h I__1030 (
            .O(N__12081),
            .I(N__12078));
    Span4Mux_v I__1029 (
            .O(N__12078),
            .I(N__12075));
    Sp12to4 I__1028 (
            .O(N__12075),
            .I(N__12072));
    Span12Mux_v I__1027 (
            .O(N__12072),
            .I(N__12069));
    Odrv12 I__1026 (
            .O(N__12069),
            .I(this_vga_signals_vsync_1_i));
    InMux I__1025 (
            .O(N__12066),
            .I(N__12063));
    LocalMux I__1024 (
            .O(N__12063),
            .I(\this_vga_signals.vsync_1_2 ));
    InMux I__1023 (
            .O(N__12060),
            .I(N__12057));
    LocalMux I__1022 (
            .O(N__12057),
            .I(\this_vga_signals.vsync_1_3 ));
    CascadeMux I__1021 (
            .O(N__12054),
            .I(\this_vga_signals.mult1_un47_sum_c3_1_1_0_cascade_ ));
    IoInMux I__1020 (
            .O(N__12051),
            .I(N__12048));
    LocalMux I__1019 (
            .O(N__12048),
            .I(N__12045));
    Span12Mux_s10_h I__1018 (
            .O(N__12045),
            .I(N__12042));
    Odrv12 I__1017 (
            .O(N__12042),
            .I(rgb_c_0));
    CascadeMux I__1016 (
            .O(N__12039),
            .I(\this_vga_ramdac.i2_mux_cascade_ ));
    InMux I__1015 (
            .O(N__12036),
            .I(N__12033));
    LocalMux I__1014 (
            .O(N__12033),
            .I(N__12029));
    InMux I__1013 (
            .O(N__12032),
            .I(N__12026));
    Odrv12 I__1012 (
            .O(N__12029),
            .I(\this_vga_ramdac.N_3300_reto ));
    LocalMux I__1011 (
            .O(N__12026),
            .I(\this_vga_ramdac.N_3300_reto ));
    CascadeMux I__1010 (
            .O(N__12021),
            .I(\this_vga_ramdac.m6_cascade_ ));
    InMux I__1009 (
            .O(N__12018),
            .I(N__12015));
    LocalMux I__1008 (
            .O(N__12015),
            .I(N__12012));
    Span4Mux_v I__1007 (
            .O(N__12012),
            .I(N__12008));
    InMux I__1006 (
            .O(N__12011),
            .I(N__12005));
    Odrv4 I__1005 (
            .O(N__12008),
            .I(\this_vga_ramdac.N_3299_reto ));
    LocalMux I__1004 (
            .O(N__12005),
            .I(\this_vga_ramdac.N_3299_reto ));
    IoInMux I__1003 (
            .O(N__12000),
            .I(N__11997));
    LocalMux I__1002 (
            .O(N__11997),
            .I(N__11994));
    Span4Mux_s2_h I__1001 (
            .O(N__11994),
            .I(N__11991));
    Span4Mux_h I__1000 (
            .O(N__11991),
            .I(N__11988));
    Span4Mux_h I__999 (
            .O(N__11988),
            .I(N__11985));
    Sp12to4 I__998 (
            .O(N__11985),
            .I(N__11982));
    Odrv12 I__997 (
            .O(N__11982),
            .I(rgb_c_5));
    CascadeMux I__996 (
            .O(N__11979),
            .I(N__11976));
    InMux I__995 (
            .O(N__11976),
            .I(N__11973));
    LocalMux I__994 (
            .O(N__11973),
            .I(N__11970));
    Odrv4 I__993 (
            .O(N__11970),
            .I(\this_vga_signals.N_729 ));
    InMux I__992 (
            .O(N__11967),
            .I(un1_M_this_map_address_q_cry_1));
    CascadeMux I__991 (
            .O(N__11964),
            .I(N__11961));
    CascadeBuf I__990 (
            .O(N__11961),
            .I(N__11958));
    CascadeMux I__989 (
            .O(N__11958),
            .I(N__11955));
    InMux I__988 (
            .O(N__11955),
            .I(N__11952));
    LocalMux I__987 (
            .O(N__11952),
            .I(N__11948));
    InMux I__986 (
            .O(N__11951),
            .I(N__11945));
    Span4Mux_h I__985 (
            .O(N__11948),
            .I(N__11942));
    LocalMux I__984 (
            .O(N__11945),
            .I(M_this_map_address_qZ0Z_3));
    Odrv4 I__983 (
            .O(N__11942),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__982 (
            .O(N__11937),
            .I(un1_M_this_map_address_q_cry_2));
    CascadeMux I__981 (
            .O(N__11934),
            .I(N__11931));
    CascadeBuf I__980 (
            .O(N__11931),
            .I(N__11928));
    CascadeMux I__979 (
            .O(N__11928),
            .I(N__11925));
    InMux I__978 (
            .O(N__11925),
            .I(N__11922));
    LocalMux I__977 (
            .O(N__11922),
            .I(N__11918));
    InMux I__976 (
            .O(N__11921),
            .I(N__11915));
    Span4Mux_h I__975 (
            .O(N__11918),
            .I(N__11912));
    LocalMux I__974 (
            .O(N__11915),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__973 (
            .O(N__11912),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__972 (
            .O(N__11907),
            .I(un1_M_this_map_address_q_cry_3));
    CascadeMux I__971 (
            .O(N__11904),
            .I(N__11901));
    CascadeBuf I__970 (
            .O(N__11901),
            .I(N__11898));
    CascadeMux I__969 (
            .O(N__11898),
            .I(N__11895));
    InMux I__968 (
            .O(N__11895),
            .I(N__11892));
    LocalMux I__967 (
            .O(N__11892),
            .I(N__11888));
    InMux I__966 (
            .O(N__11891),
            .I(N__11885));
    Span4Mux_h I__965 (
            .O(N__11888),
            .I(N__11882));
    LocalMux I__964 (
            .O(N__11885),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__963 (
            .O(N__11882),
            .I(M_this_map_address_qZ0Z_5));
    InMux I__962 (
            .O(N__11877),
            .I(un1_M_this_map_address_q_cry_4));
    CascadeMux I__961 (
            .O(N__11874),
            .I(N__11871));
    CascadeBuf I__960 (
            .O(N__11871),
            .I(N__11868));
    CascadeMux I__959 (
            .O(N__11868),
            .I(N__11865));
    InMux I__958 (
            .O(N__11865),
            .I(N__11862));
    LocalMux I__957 (
            .O(N__11862),
            .I(N__11858));
    InMux I__956 (
            .O(N__11861),
            .I(N__11855));
    Span4Mux_h I__955 (
            .O(N__11858),
            .I(N__11852));
    LocalMux I__954 (
            .O(N__11855),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__953 (
            .O(N__11852),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__952 (
            .O(N__11847),
            .I(un1_M_this_map_address_q_cry_5));
    CascadeMux I__951 (
            .O(N__11844),
            .I(N__11841));
    CascadeBuf I__950 (
            .O(N__11841),
            .I(N__11838));
    CascadeMux I__949 (
            .O(N__11838),
            .I(N__11835));
    InMux I__948 (
            .O(N__11835),
            .I(N__11832));
    LocalMux I__947 (
            .O(N__11832),
            .I(N__11828));
    InMux I__946 (
            .O(N__11831),
            .I(N__11825));
    Span4Mux_h I__945 (
            .O(N__11828),
            .I(N__11822));
    LocalMux I__944 (
            .O(N__11825),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__943 (
            .O(N__11822),
            .I(M_this_map_address_qZ0Z_7));
    InMux I__942 (
            .O(N__11817),
            .I(un1_M_this_map_address_q_cry_6));
    CascadeMux I__941 (
            .O(N__11814),
            .I(N__11811));
    CascadeBuf I__940 (
            .O(N__11811),
            .I(N__11808));
    CascadeMux I__939 (
            .O(N__11808),
            .I(N__11805));
    InMux I__938 (
            .O(N__11805),
            .I(N__11802));
    LocalMux I__937 (
            .O(N__11802),
            .I(N__11798));
    InMux I__936 (
            .O(N__11801),
            .I(N__11795));
    Span4Mux_h I__935 (
            .O(N__11798),
            .I(N__11792));
    LocalMux I__934 (
            .O(N__11795),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__933 (
            .O(N__11792),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__932 (
            .O(N__11787),
            .I(bfn_10_28_0_));
    InMux I__931 (
            .O(N__11784),
            .I(un1_M_this_map_address_q_cry_8));
    CascadeMux I__930 (
            .O(N__11781),
            .I(N__11778));
    CascadeBuf I__929 (
            .O(N__11778),
            .I(N__11775));
    CascadeMux I__928 (
            .O(N__11775),
            .I(N__11772));
    InMux I__927 (
            .O(N__11772),
            .I(N__11769));
    LocalMux I__926 (
            .O(N__11769),
            .I(N__11765));
    InMux I__925 (
            .O(N__11768),
            .I(N__11762));
    Span4Mux_h I__924 (
            .O(N__11765),
            .I(N__11759));
    LocalMux I__923 (
            .O(N__11762),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__922 (
            .O(N__11759),
            .I(M_this_map_address_qZ0Z_9));
    IoInMux I__921 (
            .O(N__11754),
            .I(N__11751));
    LocalMux I__920 (
            .O(N__11751),
            .I(N__11748));
    Span12Mux_s1_h I__919 (
            .O(N__11748),
            .I(N__11745));
    Odrv12 I__918 (
            .O(N__11745),
            .I(rgb_c_2));
    IoInMux I__917 (
            .O(N__11742),
            .I(N__11739));
    LocalMux I__916 (
            .O(N__11739),
            .I(N__11736));
    Odrv12 I__915 (
            .O(N__11736),
            .I(rgb_c_1));
    IoInMux I__914 (
            .O(N__11733),
            .I(N__11730));
    LocalMux I__913 (
            .O(N__11730),
            .I(N__11727));
    IoSpan4Mux I__912 (
            .O(N__11727),
            .I(N__11724));
    Span4Mux_s2_h I__911 (
            .O(N__11724),
            .I(N__11721));
    Span4Mux_h I__910 (
            .O(N__11721),
            .I(N__11718));
    Span4Mux_v I__909 (
            .O(N__11718),
            .I(N__11715));
    Span4Mux_v I__908 (
            .O(N__11715),
            .I(N__11712));
    Odrv4 I__907 (
            .O(N__11712),
            .I(rgb_c_4));
    InMux I__906 (
            .O(N__11709),
            .I(N__11706));
    LocalMux I__905 (
            .O(N__11706),
            .I(N__11703));
    Odrv4 I__904 (
            .O(N__11703),
            .I(M_this_map_ram_write_data_4));
    CascadeMux I__903 (
            .O(N__11700),
            .I(N__11697));
    InMux I__902 (
            .O(N__11697),
            .I(N__11694));
    LocalMux I__901 (
            .O(N__11694),
            .I(N__11691));
    Odrv4 I__900 (
            .O(N__11691),
            .I(N_393_0));
    IoInMux I__899 (
            .O(N__11688),
            .I(N__11685));
    LocalMux I__898 (
            .O(N__11685),
            .I(N__11682));
    IoSpan4Mux I__897 (
            .O(N__11682),
            .I(N__11679));
    Span4Mux_s1_h I__896 (
            .O(N__11679),
            .I(N__11676));
    Span4Mux_h I__895 (
            .O(N__11676),
            .I(N__11673));
    Span4Mux_h I__894 (
            .O(N__11673),
            .I(N__11670));
    Odrv4 I__893 (
            .O(N__11670),
            .I(rgb_c_3));
    CascadeMux I__892 (
            .O(N__11667),
            .I(N__11664));
    CascadeBuf I__891 (
            .O(N__11664),
            .I(N__11661));
    CascadeMux I__890 (
            .O(N__11661),
            .I(N__11658));
    InMux I__889 (
            .O(N__11658),
            .I(N__11654));
    InMux I__888 (
            .O(N__11657),
            .I(N__11651));
    LocalMux I__887 (
            .O(N__11654),
            .I(N__11648));
    LocalMux I__886 (
            .O(N__11651),
            .I(N__11643));
    Span4Mux_v I__885 (
            .O(N__11648),
            .I(N__11643));
    Odrv4 I__884 (
            .O(N__11643),
            .I(M_this_map_address_qZ0Z_0));
    CascadeMux I__883 (
            .O(N__11640),
            .I(N__11637));
    CascadeBuf I__882 (
            .O(N__11637),
            .I(N__11634));
    CascadeMux I__881 (
            .O(N__11634),
            .I(N__11631));
    InMux I__880 (
            .O(N__11631),
            .I(N__11628));
    LocalMux I__879 (
            .O(N__11628),
            .I(N__11624));
    InMux I__878 (
            .O(N__11627),
            .I(N__11621));
    Span4Mux_v I__877 (
            .O(N__11624),
            .I(N__11618));
    LocalMux I__876 (
            .O(N__11621),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__875 (
            .O(N__11618),
            .I(M_this_map_address_qZ0Z_1));
    InMux I__874 (
            .O(N__11613),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__873 (
            .O(N__11610),
            .I(N__11607));
    CascadeBuf I__872 (
            .O(N__11607),
            .I(N__11604));
    CascadeMux I__871 (
            .O(N__11604),
            .I(N__11601));
    InMux I__870 (
            .O(N__11601),
            .I(N__11598));
    LocalMux I__869 (
            .O(N__11598),
            .I(N__11594));
    InMux I__868 (
            .O(N__11597),
            .I(N__11591));
    Span4Mux_h I__867 (
            .O(N__11594),
            .I(N__11588));
    LocalMux I__866 (
            .O(N__11591),
            .I(M_this_map_address_qZ0Z_2));
    Odrv4 I__865 (
            .O(N__11588),
            .I(M_this_map_address_qZ0Z_2));
    IoInMux I__864 (
            .O(N__11583),
            .I(N__11580));
    LocalMux I__863 (
            .O(N__11580),
            .I(port_data_rw_i_i));
    IoInMux I__862 (
            .O(N__11577),
            .I(N__11574));
    LocalMux I__861 (
            .O(N__11574),
            .I(N__11571));
    Odrv12 I__860 (
            .O(N__11571),
            .I(port_nmib_0_i));
    IoInMux I__859 (
            .O(N__11568),
            .I(N__11565));
    LocalMux I__858 (
            .O(N__11565),
            .I(N__11562));
    Odrv12 I__857 (
            .O(N__11562),
            .I(this_vga_signals_vvisibility_i));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_20_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_6_0_));
    defparam IN_MUX_bfv_20_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_7_0_ (
            .carryinitin(\this_ppu.un1_M_vaddress_q_cry_7 ),
            .carryinitout(bfn_20_7_0_));
    defparam IN_MUX_bfv_19_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_5_0_));
    defparam IN_MUX_bfv_19_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_6_0_ (
            .carryinitin(\this_ppu.un1_M_haddress_q_cry_7 ),
            .carryinitout(bfn_19_6_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_21_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_22_0_));
    defparam IN_MUX_bfv_21_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_23_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_21_23_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_24_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_11_0_));
    defparam IN_MUX_bfv_21_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_6_0_));
    defparam IN_MUX_bfv_21_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_7_0_ (
            .carryinitin(\this_ppu.un1_M_vaddress_q_3_cry_7 ),
            .carryinitout(bfn_21_7_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_19_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_8_0_ (
            .carryinitin(\this_ppu.un1_M_haddress_q_2_cry_7 ),
            .carryinitout(bfn_19_8_0_));
    defparam IN_MUX_bfv_19_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_22_0_));
    defparam IN_MUX_bfv_19_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_23_0_ (
            .carryinitin(un1_M_this_sprites_address_q_cry_7),
            .carryinitout(bfn_19_23_0_));
    defparam IN_MUX_bfv_10_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_27_0_));
    defparam IN_MUX_bfv_10_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_28_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_10_28_0_));
    defparam IN_MUX_bfv_26_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_21_0_));
    defparam IN_MUX_bfv_26_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_22_0_ (
            .carryinitin(M_this_external_address_q_cry_7),
            .carryinitout(bfn_26_22_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__14700),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_1332_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_9  (
            .USERSIGNALTOGLOBALBUFFER(N__29698),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__25017),
            .GLOBALBUFFEROUTPUT(N_404_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.port_data_rw_i_i_LC_1_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.port_data_rw_i_i_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.port_data_rw_i_i_LC_1_21_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_vga_signals.port_data_rw_i_i_LC_1_21_1  (
            .in0(N__25547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24980),
            .lcout(port_data_rw_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNINGI76_7_LC_4_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINGI76_7_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINGI76_7_LC_4_11_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNINGI76_7_LC_4_11_7  (
            .in0(N__24979),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20603),
            .lcout(port_nmib_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_15_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_15_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_15_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_7_LC_5_29_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_7_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_7_LC_5_29_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_0_7_LC_5_29_3  (
            .in0(N__20604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_17_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__12036),
            .in2(_gnd_net_),
            .in3(N__12276),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_18_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_18_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(N__12018),
            .in2(_gnd_net_),
            .in3(N__12275),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_9_19_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_9_19_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_9_19_6  (
            .in0(N__12477),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12268),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_4_LC_9_28_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_4_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_4_LC_9_28_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_4_LC_9_28_4  (
            .in0(N__32417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25294),
            .lcout(M_this_map_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI88JG2_9_LC_10_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI88JG2_9_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI88JG2_9_LC_10_17_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI88JG2_9_LC_10_17_4  (
            .in0(N__20593),
            .in1(N__15831),
            .in2(N__11979),
            .in3(N__15678),
            .lcout(N_393_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_10_19_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_10_19_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_10_19_3  (
            .in0(N__12195),
            .in1(N__12258),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_0_LC_10_27_0.C_ON=1'b1;
    defparam M_this_map_address_q_0_LC_10_27_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_10_27_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_0_LC_10_27_0 (
            .in0(N__25346),
            .in1(N__11657),
            .in2(N__25291),
            .in3(N__25295),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_10_27_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_1_LC_10_27_1.C_ON=1'b1;
    defparam M_this_map_address_q_1_LC_10_27_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_10_27_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_1_LC_10_27_1 (
            .in0(N__25352),
            .in1(N__11627),
            .in2(_gnd_net_),
            .in3(N__11613),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_2_LC_10_27_2.C_ON=1'b1;
    defparam M_this_map_address_q_2_LC_10_27_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_10_27_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_2_LC_10_27_2 (
            .in0(N__25347),
            .in1(N__11597),
            .in2(_gnd_net_),
            .in3(N__11967),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_3_LC_10_27_3.C_ON=1'b1;
    defparam M_this_map_address_q_3_LC_10_27_3.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_10_27_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_3_LC_10_27_3 (
            .in0(N__25353),
            .in1(N__11951),
            .in2(_gnd_net_),
            .in3(N__11937),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_4_LC_10_27_4.C_ON=1'b1;
    defparam M_this_map_address_q_4_LC_10_27_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_10_27_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_4_LC_10_27_4 (
            .in0(N__25348),
            .in1(N__11921),
            .in2(_gnd_net_),
            .in3(N__11907),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_5_LC_10_27_5.C_ON=1'b1;
    defparam M_this_map_address_q_5_LC_10_27_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_10_27_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_5_LC_10_27_5 (
            .in0(N__25350),
            .in1(N__11891),
            .in2(_gnd_net_),
            .in3(N__11877),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_6_LC_10_27_6.C_ON=1'b1;
    defparam M_this_map_address_q_6_LC_10_27_6.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_10_27_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_6_LC_10_27_6 (
            .in0(N__25349),
            .in1(N__11861),
            .in2(_gnd_net_),
            .in3(N__11847),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_7_LC_10_27_7.C_ON=1'b1;
    defparam M_this_map_address_q_7_LC_10_27_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_10_27_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_7_LC_10_27_7 (
            .in0(N__25351),
            .in1(N__11831),
            .in2(_gnd_net_),
            .in3(N__11817),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(N__36963),
            .ce(),
            .sr(N__32207));
    defparam M_this_map_address_q_8_LC_10_28_0.C_ON=1'b1;
    defparam M_this_map_address_q_8_LC_10_28_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_10_28_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_8_LC_10_28_0 (
            .in0(N__25357),
            .in1(N__11801),
            .in2(_gnd_net_),
            .in3(N__11787),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_10_28_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(N__36966),
            .ce(),
            .sr(N__32205));
    defparam M_this_map_address_q_9_LC_10_28_1.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_10_28_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_10_28_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_map_address_q_9_LC_10_28_1 (
            .in0(N__11768),
            .in1(N__25358),
            .in2(_gnd_net_),
            .in3(N__11784),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36966),
            .ce(),
            .sr(N__32205));
    defparam \this_vga_signals.un5_vaddress_g0_39_LC_11_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_39_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_39_LC_11_14_2 .LUT_INIT=16'b1000010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_39_LC_11_14_2  (
            .in0(N__17331),
            .in1(N__17160),
            .in2(N__16505),
            .in3(N__17058),
            .lcout(\this_vga_signals.N_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_5_LC_11_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_5_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_5_LC_11_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_5_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__16783),
            .in2(_gnd_net_),
            .in3(N__16367),
            .lcout(\this_vga_signals.g2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_11_17_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_11_17_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_11_17_1  (
            .in0(N__12262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12861),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_11_17_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_11_17_2 .LUT_INIT=16'b0000011001110111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_11_17_2  (
            .in0(N__12403),
            .in1(N__12338),
            .in2(N__12440),
            .in3(N__12369),
            .lcout(),
            .ltout(\this_vga_ramdac.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_17_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_17_3 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_11_17_3  (
            .in0(N__12032),
            .in1(N__29685),
            .in2(N__12039),
            .in3(N__12895),
            .lcout(\this_vga_ramdac.N_3300_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36909),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6 .LUT_INIT=16'b0001000111111011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_11_17_6  (
            .in0(N__12404),
            .in1(N__12339),
            .in2(N__12441),
            .in3(N__12370),
            .lcout(),
            .ltout(\this_vga_ramdac.m6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_17_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_17_7 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_11_17_7  (
            .in0(N__12011),
            .in1(N__29684),
            .in2(N__12021),
            .in3(N__12894),
            .lcout(\this_vga_ramdac.N_3299_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36909),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_11_18_0 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_11_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12293),
            .lcout(this_pixel_clk_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36920),
            .ce(),
            .sr(N__36028));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_11_19_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_11_19_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_11_19_1  (
            .in0(N__12456),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12244),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_11_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_11_19_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__15599),
            .in2(_gnd_net_),
            .in3(N__15069),
            .lcout(\this_vga_signals.N_729 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_21_2 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_11_21_2  (
            .in0(N__15597),
            .in1(N__15825),
            .in2(_gnd_net_),
            .in3(N__15672),
            .lcout(N_495),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_13_0 .LUT_INIT=16'b0000000100001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_13_0  (
            .in0(N__14945),
            .in1(N__14873),
            .in2(N__16811),
            .in3(N__16909),
            .lcout(),
            .ltout(\this_vga_signals.un2_vsynclt8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_13_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_13_1  (
            .in0(N__12066),
            .in1(N__12060),
            .in2(N__12093),
            .in3(N__16447),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_13_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_13_2  (
            .in0(N__14946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17412),
            .lcout(\this_vga_signals.vsync_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_13_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_13_3  (
            .in0(N__16765),
            .in1(N__16350),
            .in2(N__14797),
            .in3(N__16224),
            .lcout(\this_vga_signals.vsync_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_12_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_12_13_4 .LUT_INIT=16'b0110110110110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_40_LC_12_13_4  (
            .in0(N__16223),
            .in1(N__17411),
            .in2(N__16476),
            .in3(N__14783),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_2_LC_12_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_2_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_2_LC_12_13_5 .LUT_INIT=16'b0110110010010011;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_2_LC_12_13_5  (
            .in0(N__16764),
            .in1(N__16446),
            .in2(N__16377),
            .in3(N__17140),
            .lcout(\this_vga_signals.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_12_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_12_13_6 .LUT_INIT=16'b1101010000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_38_LC_12_13_6  (
            .in0(N__17139),
            .in1(N__17302),
            .in2(N__12165),
            .in3(N__17045),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_1_1_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_12_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_12_13_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_36_LC_12_13_7  (
            .in0(N__17303),
            .in1(_gnd_net_),
            .in2(N__12054),
            .in3(N__16795),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_12_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_12_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_2_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__17313),
            .in2(_gnd_net_),
            .in3(N__15406),
            .lcout(\this_vga_signals.g0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_2_LC_12_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_2_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_2_LC_12_14_2 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_2_LC_12_14_2  (
            .in0(N__15408),
            .in1(N__16478),
            .in2(_gnd_net_),
            .in3(N__16365),
            .lcout(\this_vga_signals.vaddress_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_14_3 .LUT_INIT=16'b0110101111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_12_14_3  (
            .in0(N__17395),
            .in1(N__14367),
            .in2(N__16222),
            .in3(N__14753),
            .lcout(\this_vga_signals.if_m8_0_a3_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_1_LC_12_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_1_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_1_LC_12_14_4 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_1_LC_12_14_4  (
            .in0(N__15407),
            .in1(N__16477),
            .in2(_gnd_net_),
            .in3(N__16366),
            .lcout(\this_vga_signals.vaddress_5_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_0_LC_12_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_0_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_0_LC_12_14_5 .LUT_INIT=16'b0011000001110101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_0_LC_12_14_5  (
            .in0(N__12156),
            .in1(N__12150),
            .in2(N__12144),
            .in3(N__17314),
            .lcout(),
            .ltout(\this_vga_signals.g0_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_12_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_37_LC_12_14_6 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_37_LC_12_14_6  (
            .in0(N__16766),
            .in1(N__12135),
            .in2(N__12129),
            .in3(N__16109),
            .lcout(),
            .ltout(\this_vga_signals.N_4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_12_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_12_14_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_34_LC_12_14_7  (
            .in0(N__16110),
            .in1(N__12126),
            .in2(N__12117),
            .in3(N__14505),
            .lcout(\this_vga_signals.N_3_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_12_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_12_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_12_15_0  (
            .in0(N__16368),
            .in1(N__16217),
            .in2(N__16506),
            .in3(N__17406),
            .lcout(\this_vga_signals.M_vcounter_d7lto8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13359),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36893),
            .ce(N__14157),
            .sr(N__14109));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_12_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_12_15_3 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x0_LC_12_15_3  (
            .in0(N__17311),
            .in1(N__16148),
            .in2(N__16793),
            .in3(N__16093),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4  (
            .in0(N__12636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36893),
            .ce(N__14157),
            .sr(N__14109));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_15_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_15_5  (
            .in0(N__16364),
            .in1(N__12216),
            .in2(_gnd_net_),
            .in3(N__15405),
            .lcout(),
            .ltout(\this_vga_signals.if_N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_12_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_LC_12_15_6 .LUT_INIT=16'b0000110100001110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_LC_12_15_6  (
            .in0(N__15909),
            .in1(N__17310),
            .in2(N__12210),
            .in3(N__17118),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x1_LC_12_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x1_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x1_LC_12_15_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_x1_LC_12_15_7  (
            .in0(N__17312),
            .in1(N__16789),
            .in2(N__12207),
            .in3(N__16094),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_12_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_12_16_0 .LUT_INIT=16'b1110011100011000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_N_4L6_LC_12_16_0  (
            .in0(N__12204),
            .in1(N__17315),
            .in2(N__16819),
            .in3(N__16121),
            .lcout(\this_vga_signals.g0_31_N_4L6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_12_16_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_12_16_1 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_12_16_1  (
            .in0(N__12171),
            .in1(N__29711),
            .in2(N__12191),
            .in3(N__12896),
            .lcout(\this_vga_ramdac.N_3301_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36897),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBCAC_6_LC_12_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBCAC_6_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBCAC_6_LC_12_16_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBCAC_6_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__16501),
            .in2(_gnd_net_),
            .in3(N__15710),
            .lcout(),
            .ltout(\this_vga_signals.vvisibility_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_7_LC_12_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_7_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_7_LC_12_16_5 .LUT_INIT=16'b0000000011100111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5JIE1_7_LC_12_16_5  (
            .in0(N__16218),
            .in1(N__17407),
            .in2(N__12174),
            .in3(N__14798),
            .lcout(this_vga_signals_vvisibility),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_17_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_17_1 .LUT_INIT=16'b0100000110110111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_12_17_1  (
            .in0(N__12430),
            .in1(N__12398),
            .in2(N__12371),
            .in3(N__12334),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_12_17_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_12_17_2 .LUT_INIT=16'b0110001101001101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_12_17_2  (
            .in0(N__12337),
            .in1(N__12368),
            .in2(N__12405),
            .in3(N__12433),
            .lcout(),
            .ltout(\this_vga_ramdac.m19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_12_17_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_12_17_3 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_12_17_3  (
            .in0(N__12467),
            .in1(N__29680),
            .in2(N__12480),
            .in3(N__12891),
            .lcout(\this_vga_ramdac.N_3302_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36903),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_12_17_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_12_17_4 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_12_17_4  (
            .in0(N__12892),
            .in1(N__12452),
            .in2(N__29699),
            .in3(N__12309),
            .lcout(\this_vga_ramdac.N_3303_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36903),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_12_17_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_12_17_5 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_12_17_5  (
            .in0(N__12431),
            .in1(N__12397),
            .in2(_gnd_net_),
            .in3(N__12336),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_12_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_12_17_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_RNIH7PG8_LC_12_17_6  (
            .in0(N__12726),
            .in1(N__13606),
            .in2(_gnd_net_),
            .in3(N__13568),
            .lcout(M_pcounter_q_ret_2_RNIH7PG8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_12_17_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_12_17_7 .LUT_INIT=16'b0000101101100011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_12_17_7  (
            .in0(N__12432),
            .in1(N__12399),
            .in2(N__12372),
            .in3(N__12335),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_12_18_0 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_12_18_0 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_12_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_12_18_0  (
            .in0(N__36087),
            .in1(N__12303),
            .in2(_gnd_net_),
            .in3(N__12294),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36910),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.G_394_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.G_394_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.G_394_LC_12_18_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.G_394_LC_12_18_1  (
            .in0(N__12302),
            .in1(N__12292),
            .in2(_gnd_net_),
            .in3(N__36086),
            .lcout(\this_vga_signals.GZ0Z_394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_12_19_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_12_19_0 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_12_19_0  (
            .in0(N__29715),
            .in1(N__13260),
            .in2(N__12257),
            .in3(N__12900),
            .lcout(\this_vga_ramdac.N_880_i_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36921),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_12_19_1 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3SF72_9_LC_12_19_1  (
            .in0(N__15827),
            .in1(N__15673),
            .in2(N__20589),
            .in3(N__15598),
            .lcout(N_880_0),
            .ltout(N_880_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIITNT4_9_LC_12_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIITNT4_9_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIITNT4_9_LC_12_19_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIITNT4_9_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12573),
            .in3(N__13818),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNILLQLK_9_LC_12_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNILLQLK_9_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNILLQLK_9_LC_12_19_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNILLQLK_9_LC_12_19_5  (
            .in0(N__13258),
            .in1(N__13782),
            .in2(_gnd_net_),
            .in3(N__13668),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS7VH6_9_LC_12_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS7VH6_9_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS7VH6_9_LC_12_19_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIS7VH6_9_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__13259),
            .in2(_gnd_net_),
            .in3(N__14019),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_12_20_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12513),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36926),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_12_20_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_12_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12525),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36926),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_1_LC_12_27_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_1_LC_12_27_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_1_LC_12_27_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_1_LC_12_27_3  (
            .in0(N__33311),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25229),
            .lcout(M_this_map_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_5_LC_12_27_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_5_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_5_LC_12_27_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_5_LC_12_27_7  (
            .in0(N__36360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25230),
            .lcout(M_this_map_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_12_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_13_12_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_13_12_0  (
            .in0(N__17682),
            .in1(N__12718),
            .in2(N__13923),
            .in3(N__13921),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__36861),
            .ce(),
            .sr(N__14106));
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_12_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_12_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_13_12_1  (
            .in0(N__17684),
            .in1(N__14872),
            .in2(_gnd_net_),
            .in3(N__12483),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__36861),
            .ce(),
            .sr(N__14106));
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_12_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_12_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_13_12_2  (
            .in0(N__17683),
            .in1(N__14944),
            .in2(_gnd_net_),
            .in3(N__12597),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__36861),
            .ce(),
            .sr(N__14106));
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_12_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_12_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_13_12_3  (
            .in0(N__17685),
            .in1(N__16908),
            .in2(_gnd_net_),
            .in3(N__12594),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__36861),
            .ce(),
            .sr(N__14106));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_12_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__16718),
            .in2(_gnd_net_),
            .in3(N__12591),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_12_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__16375),
            .in2(_gnd_net_),
            .in3(N__12588),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_12_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__16495),
            .in2(_gnd_net_),
            .in3(N__12585),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_12_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__17421),
            .in2(_gnd_net_),
            .in3(N__12582),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_13_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__16233),
            .in2(_gnd_net_),
            .in3(N__12579),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_13_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_13_13_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__14790),
            .in2(_gnd_net_),
            .in3(N__12576),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36869),
            .ce(N__14154),
            .sr(N__14108));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_13_13_2  (
            .in0(N__12632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36869),
            .ce(N__14154),
            .sr(N__14108));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_13_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12631),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36869),
            .ce(N__14154),
            .sr(N__14108));
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_13_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_13_14_1 .LUT_INIT=16'b0100011010010001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_18_LC_13_14_1  (
            .in0(N__14415),
            .in1(N__17309),
            .in2(N__14406),
            .in3(N__17138),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_13_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_13_14_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_13_14_2  (
            .in0(N__13383),
            .in1(N__13290),
            .in2(N__14214),
            .in3(N__12618),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_13_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_13_14_3 .LUT_INIT=16'b0000101100011101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_13_14_3  (
            .in0(N__13407),
            .in1(N__14240),
            .in2(N__12612),
            .in3(N__14752),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_13_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_13_14_4 .LUT_INIT=16'b1101000010110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_13_14_4  (
            .in0(N__14366),
            .in1(N__12603),
            .in2(N__12609),
            .in3(N__15703),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_14_5 .LUT_INIT=16'b0001100011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_14_5  (
            .in0(N__15906),
            .in1(N__17308),
            .in2(N__12606),
            .in3(N__17026),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_13_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_13_14_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_a3_a7_LC_13_14_6  (
            .in0(N__13382),
            .in1(_gnd_net_),
            .in2(N__14213),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_13_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_13_14_7 .LUT_INIT=16'b0011111100101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_13_14_7  (
            .in0(N__13406),
            .in1(N__14239),
            .in2(N__14770),
            .in3(N__14365),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_13_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_13_15_0 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_13_15_0  (
            .in0(N__14876),
            .in1(N__14985),
            .in2(_gnd_net_),
            .in3(N__12642),
            .lcout(),
            .ltout(\this_vga_signals.if_i1_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIIADJ4E2_7_LC_13_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIIADJ4E2_7_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIIADJ4E2_7_LC_13_15_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIIADJ4E2_7_LC_13_15_1  (
            .in0(N__15531),
            .in1(N__13518),
            .in2(N__12699),
            .in3(N__12675),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_13_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_LC_13_15_2 .LUT_INIT=16'b1001010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_LC_13_15_2  (
            .in0(N__14316),
            .in1(N__12738),
            .in2(N__14973),
            .in3(N__13445),
            .lcout(),
            .ltout(\this_vga_signals.N_5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_13_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_13_15_3 .LUT_INIT=16'b1110001110000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_LC_13_15_3  (
            .in0(N__12720),
            .in1(N__14875),
            .in2(N__12678),
            .in3(N__12660),
            .lcout(\this_vga_signals.mult1_un82_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_2_LC_13_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_2_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_2_LC_13_15_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_2_LC_13_15_5  (
            .in0(N__13499),
            .in1(N__14500),
            .in2(N__16980),
            .in3(N__16114),
            .lcout(\this_vga_signals.g0_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_0_LC_13_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_0_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_0_LC_13_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_0_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__16791),
            .in2(_gnd_net_),
            .in3(N__13500),
            .lcout(),
            .ltout(\this_vga_signals.g0_i_x4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_13_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_13_15_7 .LUT_INIT=16'b0001111011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_13_15_7  (
            .in0(N__16952),
            .in1(N__12669),
            .in2(N__12663),
            .in3(N__12768),
            .lcout(\this_vga_signals.N_3_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_13_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_13_16_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_13_16_0  (
            .in0(N__16790),
            .in1(N__14499),
            .in2(N__16981),
            .in3(N__15348),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_13_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_13_16_1 .LUT_INIT=16'b1101111111110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_LC_13_16_1  (
            .in0(N__14981),
            .in1(N__14085),
            .in2(N__12654),
            .in3(N__12651),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_13_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_13_16_2 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_13_16_2  (
            .in0(N__16554),
            .in1(N__14307),
            .in2(N__12645),
            .in3(N__13446),
            .lcout(\this_vga_signals.N_5_i_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_2_LC_13_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_2_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_2_LC_13_16_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_2_LC_13_16_3  (
            .in0(N__16948),
            .in1(N__14073),
            .in2(_gnd_net_),
            .in3(N__16122),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_13_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_13_16_4 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_13_16_4  (
            .in0(N__14948),
            .in1(N__14497),
            .in2(N__12771),
            .in3(N__13498),
            .lcout(\this_vga_signals.N_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_13_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_13_16_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_ns_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(N__12762),
            .in2(N__14634),
            .in3(N__12756),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_ns ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_N_2L1_LC_13_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_2L1_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_2L1_LC_13_16_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_N_2L1_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12750),
            .in3(N__15999),
            .lcout(),
            .ltout(\this_vga_signals.g0_31_N_2L1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_13_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_13_16_7 .LUT_INIT=16'b0111111010111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_31_N_5L8_LC_13_16_7  (
            .in0(N__14498),
            .in1(N__12747),
            .in2(N__12741),
            .in3(N__16953),
            .lcout(\this_vga_signals.g0_31_N_5L8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_17_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_13_17_1  (
            .in0(N__13896),
            .in1(N__13587),
            .in2(_gnd_net_),
            .in3(N__13556),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_13_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_13_17_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_13_17_2  (
            .in0(N__17615),
            .in1(_gnd_net_),
            .in2(N__12732),
            .in3(N__12822),
            .lcout(\this_vga_signals.N_2_0 ),
            .ltout(\this_vga_signals.N_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_13_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_13_17_3 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12729),
            .in3(N__13608),
            .lcout(\this_vga_signals.M_this_vga_signals_pixel_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36898),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_17_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIRT8S_0_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__14874),
            .in2(_gnd_net_),
            .in3(N__12719),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_d7lt3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIK8V32_2_LC_13_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIK8V32_2_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIK8V32_2_LC_13_17_5 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIK8V32_2_LC_13_17_5  (
            .in0(N__14947),
            .in1(N__16947),
            .in2(N__12909),
            .in3(N__16794),
            .lcout(\this_vga_signals.M_vcounter_d7lt9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_17_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_17_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_13_17_7  (
            .in0(N__12906),
            .in1(N__29679),
            .in2(N__12860),
            .in3(N__12893),
            .lcout(\this_vga_ramdac.N_3298_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36898),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_18_0 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_13_18_0  (
            .in0(N__13588),
            .in1(N__12820),
            .in2(N__12839),
            .in3(N__13897),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_13_18_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__12835),
            .in2(N__12843),
            .in3(N__17614),
            .lcout(\this_vga_signals.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_13_18_2 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_1_LC_13_18_2  (
            .in0(N__13590),
            .in1(N__12821),
            .in2(N__12840),
            .in3(N__13899),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36904),
            .ce(N__17669),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_13_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_13_18_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_0_LC_13_18_3  (
            .in0(N__13898),
            .in1(N__13589),
            .in2(_gnd_net_),
            .in3(N__13557),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36904),
            .ce(N__17669),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS3ODH5_9_LC_13_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS3ODH5_9_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIS3ODH5_9_LC_13_19_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIS3ODH5_9_LC_13_19_0  (
            .in0(N__13262),
            .in1(N__13209),
            .in2(_gnd_net_),
            .in3(N__13725),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_13_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_13_19_1  (
            .in0(N__13629),
            .in1(N__13218),
            .in2(N__13200),
            .in3(N__13716),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un89_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI15V0FA_9_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI15V0FA_9_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI15V0FA_9_LC_13_19_2 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI15V0FA_9_LC_13_19_2  (
            .in0(N__13261),
            .in1(N__13208),
            .in2(N__12789),
            .in3(N__13724),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIDAFV71_9_LC_13_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIDAFV71_9_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIDAFV71_9_LC_13_19_5 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIDAFV71_9_LC_13_19_5  (
            .in0(N__13266),
            .in1(N__13680),
            .in2(_gnd_net_),
            .in3(N__13179),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_13_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_13_20_0 .LUT_INIT=16'b1000111000101011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c2_LC_13_20_0  (
            .in0(N__15332),
            .in1(N__13679),
            .in2(N__17760),
            .in3(N__13178),
            .lcout(\this_vga_signals.mult1_un82_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un82_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_13_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_13_20_1 .LUT_INIT=16'b1111001100110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__13196),
            .in2(N__13212),
            .in3(N__13628),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m1_0_LC_13_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m1_0_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m1_0_LC_13_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m1_0_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__15196),
            .in2(_gnd_net_),
            .in3(N__14007),
            .lcout(\this_vga_signals.if_m7_0_x4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc1_LC_13_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc1_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc1_LC_13_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc1_LC_13_20_4  (
            .in0(N__13771),
            .in1(N__15331),
            .in2(N__15272),
            .in3(N__13667),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_0_LC_13_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_0_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_0_LC_13_20_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_0_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__13842),
            .in2(_gnd_net_),
            .in3(N__14006),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_LC_13_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_LC_13_20_6 .LUT_INIT=16'b0111100000011110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_2_LC_13_20_6  (
            .in0(N__15195),
            .in1(N__13811),
            .in2(N__13185),
            .in3(N__15126),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0_2 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__13640),
            .in2(N__13182),
            .in3(N__13770),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI1VTU_4_LC_13_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI1VTU_4_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI1VTU_4_LC_13_21_5 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \this_ppu.M_state_q_RNI1VTU_4_LC_13_21_5  (
            .in0(N__13167),
            .in1(N__13149),
            .in2(N__33939),
            .in3(N__33792),
            .lcout(M_this_ppu_sprites_addr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_0_LC_13_28_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_0_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_0_LC_13_28_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_0_LC_13_28_5  (
            .in0(_gnd_net_),
            .in1(N__31263),
            .in2(_gnd_net_),
            .in3(N__25276),
            .lcout(M_this_map_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_7_LC_13_28_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_7_LC_13_28_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_7_LC_13_28_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_7_LC_13_28_6  (
            .in0(N__25277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34581),
            .lcout(M_this_map_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14254),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36856),
            .ce(N__14155),
            .sr(N__14104));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_12_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_12_1  (
            .in0(N__14255),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36856),
            .ce(N__14155),
            .sr(N__14104));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_12_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14273),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36856),
            .ce(N__14155),
            .sr(N__14104));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14168),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36856),
            .ce(N__14155),
            .sr(N__14104));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13354),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36862),
            .ce(N__14150),
            .sr(N__14107));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_14_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_14_13_1 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_14_13_1  (
            .in0(N__13381),
            .in1(_gnd_net_),
            .in2(N__14206),
            .in3(N__13278),
            .lcout(),
            .ltout(\this_vga_signals.N_1_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_RNIE4021_LC_14_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_RNIE4021_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_RNIE4021_LC_14_13_2 .LUT_INIT=16'b1011111110101111;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_RNIE4021_LC_14_13_2  (
            .in0(N__14353),
            .in1(N__14771),
            .in2(N__13272),
            .in3(N__13405),
            .lcout(\this_vga_signals.SUM_2_i_1_2_3 ),
            .ltout(\this_vga_signals.SUM_2_i_1_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_14_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_14_13_3 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_14_13_3  (
            .in0(N__15516),
            .in1(N__15489),
            .in2(N__13269),
            .in3(N__15426),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIG08B1_LC_14_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIG08B1_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIG08B1_LC_14_13_4 .LUT_INIT=16'b1001110111011101;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIG08B1_LC_14_13_4  (
            .in0(N__14742),
            .in1(N__13404),
            .in2(N__14364),
            .in3(N__14237),
            .lcout(\this_vga_signals.SUM_2_i_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_14_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_14_13_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIU9761_5_LC_14_13_5  (
            .in0(N__14196),
            .in1(N__14741),
            .in2(N__14241),
            .in3(N__13403),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_fast_esr_RNIU9761Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_14_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_14_13_6 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61_4_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__13380),
            .in2(N__13362),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fast_esr_RNI5QL61Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_13_7  (
            .in0(N__13355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36862),
            .ce(N__14150),
            .sr(N__14107));
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_14_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_14_14_0 .LUT_INIT=16'b0100000111101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_8_LC_14_14_0  (
            .in0(N__13434),
            .in1(N__14382),
            .in2(N__13338),
            .in3(N__16166),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_14_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__13326),
            .in2(N__13320),
            .in3(N__14373),
            .lcout(\this_vga_signals.N_4_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x1_LC_14_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x1_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x1_LC_14_14_2 .LUT_INIT=16'b0011110000110110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x1_LC_14_14_2  (
            .in0(N__16720),
            .in1(N__16092),
            .in2(N__17327),
            .in3(N__14532),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_654_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_14_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_14_14_3 .LUT_INIT=16'b0111110000110100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_LC_14_14_3  (
            .in0(N__17280),
            .in1(N__17027),
            .in2(N__15907),
            .in3(N__17114),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x0_LC_14_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x0_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x0_LC_14_14_4 .LUT_INIT=16'b0111010010001011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_x0_LC_14_14_4  (
            .in0(N__16719),
            .in1(N__17282),
            .in2(N__13317),
            .in3(N__16091),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_654_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_14_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_14_14_5 .LUT_INIT=16'b1100001110111110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x0_LC_14_14_5  (
            .in0(N__16931),
            .in1(N__15992),
            .in2(N__16596),
            .in3(N__14580),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_14_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_14_14_6 .LUT_INIT=16'b0110010000011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m2_1_LC_14_14_6  (
            .in0(N__17028),
            .in1(N__15899),
            .in2(N__17141),
            .in3(N__17281),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m4_0_LC_14_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m4_0_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m4_0_LC_14_14_7 .LUT_INIT=16'b0000110000000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m4_0_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__16721),
            .in2(N__13455),
            .in3(N__16910),
            .lcout(\this_vga_signals.if_i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_14_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_14_15_0 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_ns_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__14493),
            .in2(N__14571),
            .in3(N__13452),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_14_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_14_15_1 .LUT_INIT=16'b0011001110100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_14_15_1  (
            .in0(N__14624),
            .in1(N__16161),
            .in2(N__16376),
            .in3(N__13433),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_1_x0_LC_14_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_x0_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_x0_LC_14_15_2 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_1_x0_LC_14_15_2  (
            .in0(N__17325),
            .in1(N__14536),
            .in2(N__16982),
            .in3(N__16107),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_1_ns_LC_14_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_ns_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_ns_LC_14_15_3 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_1_ns_LC_14_15_3  (
            .in0(N__16108),
            .in1(N__16961),
            .in2(N__13422),
            .in3(N__13539),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_14_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_14_15_4 .LUT_INIT=16'b0111101110110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_LC_14_15_4  (
            .in0(N__13494),
            .in1(N__14972),
            .in2(N__13419),
            .in3(N__14492),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_14_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_0_LC_14_15_5 .LUT_INIT=16'b1011001111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_0_LC_14_15_5  (
            .in0(N__16932),
            .in1(N__13416),
            .in2(N__13410),
            .in3(N__14300),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_14_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_14_15_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_14_15_7  (
            .in0(N__14625),
            .in1(N__17324),
            .in2(_gnd_net_),
            .in3(N__16732),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x0_LC_14_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x0_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x0_LC_14_16_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x0_LC_14_16_0  (
            .in0(N__16969),
            .in1(N__13496),
            .in2(N__14986),
            .in3(N__15995),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_0_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_ns_LC_14_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_ns_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_ns_LC_14_16_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_ns_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__14496),
            .in2(N__13533),
            .in3(N__13512),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0 ),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIVJPKIE_3_LC_14_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIVJPKIE_3_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIVJPKIE_3_LC_14_16_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIVJPKIE_3_LC_14_16_2  (
            .in0(N__14511),
            .in1(N__13506),
            .in2(N__13530),
            .in3(N__13461),
            .lcout(),
            .ltout(\this_vga_signals.g1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI2J0JQ31_3_LC_14_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI2J0JQ31_3_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI2J0JQ31_3_LC_14_16_3 .LUT_INIT=16'b0001111011010010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI2J0JQ31_3_LC_14_16_3  (
            .in0(N__13527),
            .in1(N__14832),
            .in2(N__13521),
            .in3(N__14430),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x1_LC_14_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x1_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x1_LC_14_16_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un82_sum_axbxc3_0_x1_LC_14_16_4  (
            .in0(N__13497),
            .in1(N__16962),
            .in2(N__14987),
            .in3(N__15993),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI6FOR21_3_LC_14_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI6FOR21_3_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI6FOR21_3_LC_14_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI6FOR21_3_LC_14_16_5  (
            .in0(N__16788),
            .in1(N__14495),
            .in2(N__16983),
            .in3(N__16123),
            .lcout(\this_vga_signals.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_14_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_14_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_14_16_6  (
            .in0(N__14494),
            .in1(N__13495),
            .in2(N__16984),
            .in3(N__15994),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_14_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_14_16_7 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_c2_LC_14_16_7  (
            .in0(N__14980),
            .in1(N__16970),
            .in2(N__13464),
            .in3(N__14299),
            .lcout(\this_vga_signals.mult1_un68_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_14_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_14_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13607),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36894),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_e_0_RNISGJ64_1_LC_14_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_e_0_RNISGJ64_1_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_e_0_RNISGJ64_1_LC_14_17_2 .LUT_INIT=16'b0100000001010101;
    LogicCell40 \this_vga_signals.M_lcounter_q_e_0_RNISGJ64_1_LC_14_17_2  (
            .in0(N__13866),
            .in1(N__16528),
            .in2(N__14825),
            .in3(N__14792),
            .lcout(\this_vga_signals.M_lcounter_d_0_sqmuxa ),
            .ltout(\this_vga_signals.M_lcounter_d_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_14_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_14_17_3 .LUT_INIT=16'b0110001010101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_14_17_3  (
            .in0(N__13952),
            .in1(N__17681),
            .in2(N__13572),
            .in3(N__13908),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36894),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_14_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_14_17_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNIPGBM_0_LC_14_17_4  (
            .in0(N__13865),
            .in1(N__13951),
            .in2(_gnd_net_),
            .in3(N__14791),
            .lcout(\this_vga_signals.line_clk_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_0_LC_14_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_0_LC_14_17_5 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \this_ppu.M_state_q_0_LC_14_17_5  (
            .in0(N__18882),
            .in1(N__29678),
            .in2(N__19671),
            .in3(N__18861),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36894),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_14_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_14_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13569),
            .lcout(\this_vga_signals.M_pcounter_q_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36894),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_14_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_14_18_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_14_18_1  (
            .in0(N__14687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17628),
            .lcout(\this_vga_signals.N_966_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_14_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_14_18_3 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_14_18_3  (
            .in0(N__17560),
            .in1(N__15256),
            .in2(N__17759),
            .in3(N__14673),
            .lcout(),
            .ltout(\this_vga_signals.M_hcounter_d7lt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_14_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_14_18_4 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_14_18_4  (
            .in0(N__15656),
            .in1(N__13827),
            .in2(N__13545),
            .in3(N__15818),
            .lcout(\this_vga_signals.M_hcounter_d7_0 ),
            .ltout(\this_vga_signals.M_hcounter_d7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_14_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_14_18_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13542),
            .in3(N__17627),
            .lcout(\this_vga_signals.M_vcounter_q_501_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_0_LC_14_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_0_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_0_LC_14_19_0 .LUT_INIT=16'b0110001100111001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_0_LC_14_19_0  (
            .in0(N__15197),
            .in1(N__13791),
            .in2(N__15263),
            .in3(N__14015),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_1_1_LC_14_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_1_1_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_1_1_LC_14_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_1_1_LC_14_19_1  (
            .in0(N__13666),
            .in1(N__15253),
            .in2(_gnd_net_),
            .in3(N__13695),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_14_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_14_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_14_19_2  (
            .in0(N__13627),
            .in1(N__13710),
            .in2(N__13728),
            .in3(N__13769),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_14_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_14_19_3 .LUT_INIT=16'b0000100101101111;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_LC_14_19_3  (
            .in0(N__15325),
            .in1(N__13626),
            .in2(N__17758),
            .in3(N__13701),
            .lcout(\this_vga_signals.mult1_un89_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_14_19_4 .LUT_INIT=16'b0111000111010100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_14_19_4  (
            .in0(N__15318),
            .in1(N__13768),
            .in2(N__15265),
            .in3(N__13664),
            .lcout(\this_vga_signals.mult1_un75_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un75_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_14_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_14_19_5 .LUT_INIT=16'b0010000110110111;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_LC_14_19_5  (
            .in0(N__13694),
            .in1(N__17748),
            .in2(N__13704),
            .in3(N__17561),
            .lcout(\this_vga_signals.if_N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_14_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_14_19_6 .LUT_INIT=16'b0000111110110010;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_14_19_6  (
            .in0(N__15317),
            .in1(N__13833),
            .in2(N__15264),
            .in3(N__13693),
            .lcout(\this_vga_signals.mult1_un75_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un75_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_14_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_14_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_14_19_7  (
            .in0(N__13665),
            .in1(N__13778),
            .in2(N__13644),
            .in3(N__13641),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_14_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_14_20_0 .LUT_INIT=16'b1001110101010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_14_20_0  (
            .in0(N__15635),
            .in1(N__15566),
            .in2(N__15064),
            .in3(N__15794),
            .lcout(\this_vga_signals.SUM_3_i_1_0 ),
            .ltout(\this_vga_signals.SUM_3_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_14_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_14_20_1 .LUT_INIT=16'b1011011001101101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_0_1_LC_14_20_1  (
            .in0(N__15058),
            .in1(N__15114),
            .in2(N__13845),
            .in3(N__14033),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_0_1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_14_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_14_20_2 .LUT_INIT=16'b1011010000101101;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_14_20_2  (
            .in0(N__15180),
            .in1(N__13810),
            .in2(N__13836),
            .in3(N__15120),
            .lcout(\this_vga_signals.if_N_8_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_14_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_14_20_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__17670),
            .in2(_gnd_net_),
            .in3(N__17497),
            .lcout(\this_vga_signals.N_966_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_14_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_14_20_4 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_14_20_4  (
            .in0(N__15115),
            .in1(N__15567),
            .in2(N__15065),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_d7lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_14_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_14_20_5 .LUT_INIT=16'b0011101100100011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_14_20_5  (
            .in0(N__15059),
            .in1(N__14034),
            .in2(N__15125),
            .in3(N__14052),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_14_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_14_20_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__15178),
            .in2(N__13794),
            .in3(N__15119),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_14_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_14_20_7 .LUT_INIT=16'b0000110101001111;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_ac0_3_0_LC_14_20_7  (
            .in0(N__15235),
            .in1(N__15181),
            .in2(N__13785),
            .in3(N__14008),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_14_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_14_21_0 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIR18F4_9_LC_14_21_0  (
            .in0(N__15798),
            .in1(N__14058),
            .in2(N__15655),
            .in3(N__13983),
            .lcout(M_hcounter_q_esr_RNIR18F4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_14_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_14_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_14_21_2  (
            .in0(N__15255),
            .in1(N__15327),
            .in2(N__17565),
            .in3(N__17756),
            .lcout(),
            .ltout(\this_vga_signals.N_473_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_6_LC_14_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_6_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_6_LC_14_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIEVMV1_6_LC_14_21_3  (
            .in0(N__15056),
            .in1(N__15191),
            .in2(N__14061),
            .in3(N__15112),
            .lcout(\this_vga_signals.N_554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_14_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_14_21_4 .LUT_INIT=16'b1011110101000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_14_21_4  (
            .in0(N__15636),
            .in1(N__15568),
            .in2(N__15814),
            .in3(N__15054),
            .lcout(\this_vga_signals.N_735_0 ),
            .ltout(\this_vga_signals.N_735_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_2_LC_14_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_2_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_2_LC_14_21_5 .LUT_INIT=16'b0111011001100001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_2_LC_14_21_5  (
            .in0(N__15055),
            .in1(N__14051),
            .in2(N__14040),
            .in3(N__15110),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_14_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_14_21_6 .LUT_INIT=16'b1110010111010000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_14_21_6  (
            .in0(N__15111),
            .in1(N__15177),
            .in2(N__14037),
            .in3(N__14032),
            .lcout(\this_vga_signals.mult1_un61_sum_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_14_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_14_21_7 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_14_21_7  (
            .in0(N__15057),
            .in1(N__15581),
            .in2(N__13977),
            .in3(N__15113),
            .lcout(\this_vga_signals.hsync_1_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_14_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_14_22_0 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_14_22_0  (
            .in0(N__15198),
            .in1(N__17757),
            .in2(N__15336),
            .in3(N__15273),
            .lcout(\this_vga_signals.N_507_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_6_LC_14_29_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_6_LC_14_29_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_6_LC_14_29_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_6_LC_14_29_7  (
            .in0(N__34455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25293),
            .lcout(M_this_map_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_e_0_1_LC_15_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_e_0_1_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_e_0_1_LC_15_12_4 .LUT_INIT=16'b0110000010101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_e_0_1_LC_15_12_4  (
            .in0(N__13859),
            .in1(N__13959),
            .in2(N__13938),
            .in3(N__13922),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36851),
            .ce(N__17688),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_15_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_15_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14178),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36857),
            .ce(N__14156),
            .sr(N__14105));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_LC_15_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_LC_15_13_2 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_LC_15_13_2  (
            .in0(N__15385),
            .in1(N__16410),
            .in2(_gnd_net_),
            .in3(N__16302),
            .lcout(\this_vga_signals.vaddress_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_15_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_15_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14283),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36857),
            .ce(N__14156),
            .sr(N__14105));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_15_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_15_13_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_15_13_4  (
            .in0(N__15384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16301),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_15_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_15_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14262),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36857),
            .ce(N__14156),
            .sr(N__14105));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_15_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_15_13_6 .LUT_INIT=16'b1010101010010101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_0_LC_15_13_6  (
            .in0(N__14238),
            .in1(N__14205),
            .in2(N__15394),
            .in3(N__14354),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_15_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_15_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14177),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36857),
            .ce(N__14156),
            .sr(N__14105));
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_15_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_15_14_0 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_27_LC_15_14_0  (
            .in0(N__14544),
            .in1(_gnd_net_),
            .in2(N__16809),
            .in3(N__17244),
            .lcout(\this_vga_signals.g1_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_2_1_LC_15_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_2_1_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_2_1_LC_15_14_1 .LUT_INIT=16'b0101000001110110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_2_1_LC_15_14_1  (
            .in0(N__17243),
            .in1(N__14626),
            .in2(N__14538),
            .in3(N__16779),
            .lcout(\this_vga_signals.g0_2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_15_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_15_14_2 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_14_LC_15_14_2  (
            .in0(N__15428),
            .in1(N__15518),
            .in2(N__15464),
            .in3(N__15494),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_15_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_15_14_3 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_LC_15_14_3  (
            .in0(N__15517),
            .in1(N__15490),
            .in2(N__15460),
            .in3(N__15427),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i_2 ),
            .ltout(\this_vga_signals.mult1_un40_sum_axb1_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_15_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_15_14_4 .LUT_INIT=16'b1101001101000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_15_14_4  (
            .in0(N__17143),
            .in1(N__14396),
            .in2(N__14385),
            .in3(N__17241),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_2 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_15_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_15_14_5 .LUT_INIT=16'b1100100101101100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_LC_15_14_5  (
            .in0(N__17242),
            .in1(N__16971),
            .in2(N__14376),
            .in3(N__16778),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_15_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_15_14_6 .LUT_INIT=16'b1100000000111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__15386),
            .in2(N__16335),
            .in3(N__14355),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(\this_vga_signals.vaddress_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_15_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_15_14_7 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_15_14_7  (
            .in0(N__17240),
            .in1(N__17142),
            .in2(N__14322),
            .in3(N__17029),
            .lcout(\this_vga_signals.mult1_un47_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_15_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_15_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_15_15_0  (
            .in0(N__16035),
            .in1(N__16026),
            .in2(N__16592),
            .in3(N__15987),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_15_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_15_15_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_15_15_1  (
            .in0(N__14488),
            .in1(_gnd_net_),
            .in2(N__14319),
            .in3(N__15951),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_15_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_15_15_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__14487),
            .in2(N__16591),
            .in3(N__15985),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_ns_LC_15_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_ns_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_ns_LC_15_15_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_654_ns_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__14630),
            .in2(N__14598),
            .in3(N__14589),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_654_ns ),
            .ltout(\this_vga_signals.mult1_un68_sum_axb1_654_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m1_3_LC_15_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_3_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_3_LC_15_15_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_3_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__16957),
            .in2(N__14583),
            .in3(N__16784),
            .lcout(\this_vga_signals.if_m1_3 ),
            .ltout(\this_vga_signals.if_m1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_15_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_15_15_5 .LUT_INIT=16'b1110010111011010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_3_0_0_x1_LC_15_15_5  (
            .in0(N__15986),
            .in1(N__16985),
            .in2(N__14574),
            .in3(N__16582),
            .lcout(\this_vga_signals.mult1_un68_sum_ac0_3_0_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_15_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_15_15_6 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_20_LC_15_15_6  (
            .in0(N__17322),
            .in1(N__17165),
            .in2(N__14559),
            .in3(N__17049),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_LC_15_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_LC_15_15_7 .LUT_INIT=16'b1100100011111001;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_LC_15_15_7  (
            .in0(N__15870),
            .in1(N__17323),
            .in2(N__16810),
            .in3(N__14537),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_15_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_LC_15_16_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_LC_15_16_0  (
            .in0(N__15003),
            .in1(N__14501),
            .in2(N__15918),
            .in3(N__16125),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_15_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_15_16_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_LC_15_16_1  (
            .in0(N__14994),
            .in1(N__14421),
            .in2(N__14439),
            .in3(N__14436),
            .lcout(\this_vga_signals.N_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_15_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_15_16_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_28_LC_15_16_2  (
            .in0(N__15864),
            .in1(N__16499),
            .in2(N__16821),
            .in3(N__17166),
            .lcout(),
            .ltout(\this_vga_signals.N_11_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_15_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_15_16_3 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_11_LC_15_16_3  (
            .in0(N__17326),
            .in1(N__15933),
            .in2(N__14424),
            .in3(N__15846),
            .lcout(\this_vga_signals.N_4_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_15_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_15_16_4 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_15_16_4  (
            .in0(N__16029),
            .in1(N__16167),
            .in2(N__16820),
            .in3(N__16124),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_15_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_15_16_5 .LUT_INIT=16'b0000101010101111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_15_16_5  (
            .in0(N__16973),
            .in1(_gnd_net_),
            .in2(N__14997),
            .in3(N__16818),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_7_LC_15_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_7_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_7_LC_15_17_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \this_ppu.M_count_q_7_LC_15_17_0  (
            .in0(N__18881),
            .in1(N__17847),
            .in2(_gnd_net_),
            .in3(N__21523),
            .lcout(\this_ppu.M_count_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36884),
            .ce(),
            .sr(N__36015));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_15_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_15_17_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__15826),
            .in2(_gnd_net_),
            .in3(N__14793),
            .lcout(\this_vga_signals.g0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m5_s_LC_15_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m5_s_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m5_s_LC_15_17_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m5_s_LC_15_17_6  (
            .in0(N__14988),
            .in1(N__14883),
            .in2(_gnd_net_),
            .in3(N__14838),
            .lcout(\this_vga_signals.if_m5_s ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_18_1 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_15_18_1  (
            .in0(N__17487),
            .in1(N__16536),
            .in2(N__14826),
            .in3(N__14799),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNI670G_1_LC_15_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNI670G_1_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNI670G_1_LC_15_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNI670G_1_LC_15_18_4  (
            .in0(N__18758),
            .in1(N__17833),
            .in2(N__17811),
            .in3(N__17776),
            .lcout(\this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI4I6I_2_LC_15_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI4I6I_2_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI4I6I_2_LC_15_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI4I6I_2_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__15316),
            .in2(_gnd_net_),
            .in3(N__15179),
            .lcout(\this_vga_signals.M_hcounter_d7lto4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_15_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_15_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_15_19_2  (
            .in0(N__14667),
            .in1(N__14652),
            .in2(_gnd_net_),
            .in3(N__28109),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_15_20_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_15_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__17548),
            .in2(N__17749),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_15_20_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_15_20_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_15_20_1  (
            .in0(N__17674),
            .in1(N__15326),
            .in2(_gnd_net_),
            .in3(N__15276),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__36905),
            .ce(),
            .sr(N__17515));
    defparam \this_vga_signals.M_hcounter_q_3_LC_15_20_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_15_20_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_15_20_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_15_20_2  (
            .in0(N__17671),
            .in1(N__15254),
            .in2(_gnd_net_),
            .in3(N__15201),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__36905),
            .ce(),
            .sr(N__17515));
    defparam \this_vga_signals.M_hcounter_q_4_LC_15_20_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_15_20_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_15_20_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_15_20_3  (
            .in0(N__17675),
            .in1(N__15190),
            .in2(_gnd_net_),
            .in3(N__15129),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__36905),
            .ce(),
            .sr(N__17515));
    defparam \this_vga_signals.M_hcounter_q_5_LC_15_20_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_15_20_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_15_20_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_15_20_4  (
            .in0(N__17672),
            .in1(N__15124),
            .in2(_gnd_net_),
            .in3(N__15072),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__36905),
            .ce(),
            .sr(N__17515));
    defparam \this_vga_signals.M_hcounter_q_6_LC_15_20_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_15_20_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_15_20_5  (
            .in0(N__17676),
            .in1(N__15063),
            .in2(_gnd_net_),
            .in3(N__15012),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__36905),
            .ce(),
            .sr(N__17515));
    defparam \this_vga_signals.M_hcounter_q_7_LC_15_20_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_15_20_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_15_20_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_15_20_6  (
            .in0(N__17673),
            .in1(N__15580),
            .in2(_gnd_net_),
            .in3(N__15009),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__36905),
            .ce(),
            .sr(N__17515));
    defparam \this_vga_signals.M_hcounter_q_8_LC_15_20_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_15_20_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_15_20_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_15_20_7  (
            .in0(N__17677),
            .in1(N__15654),
            .in2(_gnd_net_),
            .in3(N__15006),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__36905),
            .ce(),
            .sr(N__17515));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_15_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_15_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__15810),
            .in2(_gnd_net_),
            .in3(N__15834),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36911),
            .ce(N__15759),
            .sr(N__17517));
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_15_25_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_15_25_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_wclke_3_LC_15_25_5  (
            .in0(N__34995),
            .in1(N__34914),
            .in2(N__34820),
            .in3(N__34678),
            .lcout(\this_sprites_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_2_LC_15_27_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_2_LC_15_27_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_2_LC_15_27_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_2_LC_15_27_7  (
            .in0(N__35137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25290),
            .lcout(M_this_map_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_16_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_16_13_1 .LUT_INIT=16'b0111011101111110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_16_13_1  (
            .in0(N__16236),
            .in1(N__17427),
            .in2(N__16472),
            .in3(N__15714),
            .lcout(),
            .ltout(\this_vga_signals.g2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3SF72_7_LC_16_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3SF72_7_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3SF72_7_LC_16_13_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3SF72_7_LC_16_13_2  (
            .in0(N__15690),
            .in1(N__15677),
            .in2(N__15603),
            .in3(N__15600),
            .lcout(\this_vga_signals.g0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_16_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_16_14_0 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_16_14_0  (
            .in0(N__15519),
            .in1(N__15498),
            .in2(N__15468),
            .in3(N__15435),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_0_LC_16_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_0_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_0_LC_16_14_2 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIFA121_0_LC_16_14_2  (
            .in0(N__16466),
            .in1(N__16360),
            .in2(_gnd_net_),
            .in3(N__15393),
            .lcout(\this_vga_signals.vaddress_0_0_6 ),
            .ltout(\this_vga_signals.vaddress_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_16_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_16_14_3 .LUT_INIT=16'b0010010010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_25_LC_16_14_3  (
            .in0(N__17259),
            .in1(N__17153),
            .in2(N__15351),
            .in3(N__17064),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_16_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_16_14_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_30_LC_16_14_4  (
            .in0(N__16467),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16750),
            .lcout(\this_vga_signals.g0_i_i_a5_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_16_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_16_14_5 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_16_14_5  (
            .in0(N__16027),
            .in1(N__16165),
            .in2(N__16792),
            .in3(N__16115),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_16_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_16_14_6 .LUT_INIT=16'b0000110011001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_1_0_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__16972),
            .in2(N__16038),
            .in3(N__16754),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_16_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_16_14_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_16_14_7  (
            .in0(N__16028),
            .in1(N__16589),
            .in2(N__16002),
            .in3(N__15988),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_16_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_16_15_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_29_LC_16_15_0  (
            .in0(N__17161),
            .in1(N__17304),
            .in2(N__15945),
            .in3(N__15859),
            .lcout(\this_vga_signals.g0_i_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_16_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_16_15_1 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_5_LC_16_15_1  (
            .in0(N__16756),
            .in1(N__16468),
            .in2(_gnd_net_),
            .in3(N__16362),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_16_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_16_15_2 .LUT_INIT=16'b0001100011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_LC_16_15_2  (
            .in0(N__17164),
            .in1(N__17307),
            .in2(N__15927),
            .in3(N__15924),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_16_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_16_15_3 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_16_15_3  (
            .in0(N__17305),
            .in1(N__17162),
            .in2(N__15908),
            .in3(N__17062),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_16_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_16_15_4 .LUT_INIT=16'b0111101110110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_16_15_4  (
            .in0(N__16361),
            .in1(N__16755),
            .in2(N__16494),
            .in3(N__15860),
            .lcout(\this_vga_signals.N_7_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_16_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_16_15_5 .LUT_INIT=16'b0001100010100101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_16_15_5  (
            .in0(N__17306),
            .in1(N__17163),
            .in2(N__17073),
            .in3(N__17063),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_16_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_16_15_6 .LUT_INIT=16'b1101001001001011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_LC_16_15_6  (
            .in0(N__16986),
            .in1(N__16757),
            .in2(N__16599),
            .in3(N__16590),
            .lcout(\this_vga_signals.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNINAB95_1_LC_16_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNINAB95_1_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNINAB95_1_LC_16_16_0 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \this_ppu.M_state_q_RNINAB95_1_LC_16_16_0  (
            .in0(N__19897),
            .in1(N__18950),
            .in2(N__19684),
            .in3(N__19711),
            .lcout(\this_ppu.un13_0 ),
            .ltout(\this_ppu.un13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_6_LC_16_16_1 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_6_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_6_LC_16_16_1 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_6_LC_16_16_1  (
            .in0(N__18831),
            .in1(N__17346),
            .in2(N__16542),
            .in3(N__18663),
            .lcout(\this_ppu.M_count_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36868),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_16_16_2 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_16_16_2 .LUT_INIT=16'b1010001010001010;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_16_16_2  (
            .in0(N__16251),
            .in1(N__16235),
            .in2(N__16260),
            .in3(N__17423),
            .lcout(\this_ppu.M_last_q ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36868),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIO1JM4_LC_16_16_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIO1JM4_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIO1JM4_LC_16_16_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIO1JM4_LC_16_16_3  (
            .in0(N__19709),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19896),
            .lcout(\this_ppu.M_line_clk_out_0 ),
            .ltout(\this_ppu.M_line_clk_out_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIC69A5_1_LC_16_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIC69A5_1_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIC69A5_1_LC_16_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIC69A5_1_LC_16_16_4  (
            .in0(N__19673),
            .in1(N__27714),
            .in2(N__16539),
            .in3(N__27802),
            .lcout(\this_ppu.un1_M_vaddress_q_2_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_5_LC_16_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_5_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_5_LC_16_16_5 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_5_LC_16_16_5  (
            .in0(N__16535),
            .in1(N__16500),
            .in2(_gnd_net_),
            .in3(N__16363),
            .lcout(\this_vga_signals.un4_lvisibility_1 ),
            .ltout(\this_vga_signals.un4_lvisibility_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIV6084_7_LC_16_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIV6084_7_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIV6084_7_LC_16_16_6 .LUT_INIT=16'b1010001010001010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIV6084_7_LC_16_16_6  (
            .in0(N__16250),
            .in1(N__16234),
            .in2(N__16170),
            .in3(N__17422),
            .lcout(M_this_vga_signals_line_clk_0),
            .ltout(M_this_vga_signals_line_clk_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIN5VV4_LC_16_16_7 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIN5VV4_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIN5VV4_LC_16_16_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIN5VV4_LC_16_16_7  (
            .in0(N__19710),
            .in1(_gnd_net_),
            .in2(N__17364),
            .in3(N__19672),
            .lcout(\this_ppu.M_count_d_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_17_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__18580),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_17_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__28749),
            .in2(N__17781),
            .in3(N__17361),
            .lcout(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_17_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__17834),
            .in2(N__28807),
            .in3(N__17358),
            .lcout(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_17_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__28753),
            .in2(N__18759),
            .in3(N__17355),
            .lcout(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_17_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__17809),
            .in2(N__28808),
            .in3(N__17352),
            .lcout(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_17_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__28757),
            .in2(N__18606),
            .in3(N__17349),
            .lcout(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_17_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__18662),
            .in2(N__28809),
            .in3(N__17337),
            .lcout(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_17_7 .LUT_INIT=16'b1111000000011110;
    LogicCell40 \this_ppu.M_count_q_RNO_0_7_LC_16_17_7  (
            .in0(N__18951),
            .in1(N__21519),
            .in2(N__18644),
            .in3(N__17334),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_2_LC_16_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_2_LC_16_18_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_2_LC_16_18_0 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_2_LC_16_18_0  (
            .in0(N__18829),
            .in1(N__17841),
            .in2(N__18794),
            .in3(N__17835),
            .lcout(\this_ppu.M_count_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36883),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_4_LC_16_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_4_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_4_LC_16_18_4 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_4_LC_16_18_4  (
            .in0(N__18830),
            .in1(N__17817),
            .in2(N__18795),
            .in3(N__17810),
            .lcout(\this_ppu.M_count_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36883),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_1_LC_16_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_1_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_1_LC_16_18_7 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_1_LC_16_18_7  (
            .in0(N__17780),
            .in1(N__18787),
            .in2(N__17790),
            .in3(N__18828),
            .lcout(\this_ppu.M_count_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36883),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_16_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_16_19_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_16_19_0  (
            .in0(N__17556),
            .in1(N__17686),
            .in2(_gnd_net_),
            .in3(N__17732),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36892),
            .ce(),
            .sr(N__17516));
    defparam \this_vga_signals.M_hcounter_q_0_LC_16_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_16_19_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_16_19_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_16_19_1  (
            .in0(N__17687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17555),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36892),
            .ce(),
            .sr(N__17516));
    defparam \this_delay_clk.M_pipe_q_3_LC_16_20_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_16_20_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_16_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17457),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36896),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_16_20_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_16_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17466),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36896),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_21_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_21_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_21_0  (
            .in0(N__34994),
            .in1(N__34912),
            .in2(N__34819),
            .in3(N__34699),
            .lcout(\this_sprites_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_RNO_0_LC_16_21_1.C_ON=1'b0;
    defparam M_this_substate_q_RNO_0_LC_16_21_1.SEQ_MODE=4'b0000;
    defparam M_this_substate_q_RNO_0_LC_16_21_1.LUT_INIT=16'b1000100111111111;
    LogicCell40 M_this_substate_q_RNO_0_LC_16_21_1 (
            .in0(N__25711),
            .in1(N__25665),
            .in2(N__25833),
            .in3(N__31638),
            .lcout(M_this_substate_q_s_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_i_LC_16_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_i_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_i_LC_16_21_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_i_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__24900),
            .in2(_gnd_net_),
            .in3(N__36095),
            .lcout(N_49),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_464_tz_LC_16_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_464_tz_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_464_tz_LC_16_22_5 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_464_tz_LC_16_22_5  (
            .in0(N__26430),
            .in1(N__31147),
            .in2(N__23536),
            .in3(N__26519),
            .lcout(N_1294_tz_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_7_LC_16_23_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_7_LC_16_23_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_7_LC_16_23_0.LUT_INIT=16'b1010000011110011;
    LogicCell40 M_this_sprites_address_q_RNO_0_7_LC_16_23_0 (
            .in0(N__27050),
            .in1(N__26125),
            .in2(N__23782),
            .in3(N__26205),
            .lcout(M_this_sprites_address_qc_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_7_LC_16_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_7_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_7_LC_16_23_1 .LUT_INIT=16'b0000011100000101;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_7_LC_16_23_1  (
            .in0(N__23748),
            .in1(N__27052),
            .in2(N__31337),
            .in3(N__31149),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_7_LC_16_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_7_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_7_LC_16_23_2 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_7_LC_16_23_2  (
            .in0(N__25503),
            .in1(N__23705),
            .in2(N__17877),
            .in3(N__26438),
            .lcout(),
            .ltout(N_597_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_7_LC_16_23_3.C_ON=1'b0;
    defparam M_this_sprites_address_q_7_LC_16_23_3.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_7_LC_16_23_3.LUT_INIT=16'b0000111000000000;
    LogicCell40 M_this_sprites_address_q_7_LC_16_23_3 (
            .in0(N__23706),
            .in1(N__17865),
            .in2(N__17874),
            .in3(N__17871),
            .lcout(M_this_sprites_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36919),
            .ce(),
            .sr(N__32203));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_468_tz_LC_16_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_468_tz_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_468_tz_LC_16_23_4 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_468_tz_LC_16_23_4  (
            .in0(N__31148),
            .in1(N__26553),
            .in2(N__23783),
            .in3(N__26436),
            .lcout(N_1298_tz_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_8_LC_16_23_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_8_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_8_LC_16_23_5 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_8_LC_16_23_5  (
            .in0(N__26437),
            .in1(N__25504),
            .in2(N__20397),
            .in3(N__23468),
            .lcout(),
            .ltout(N_602_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_8_LC_16_23_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_8_LC_16_23_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_8_LC_16_23_6.LUT_INIT=16'b0000111000000000;
    LogicCell40 M_this_sprites_address_q_8_LC_16_23_6 (
            .in0(N__23469),
            .in1(N__17859),
            .in2(N__17850),
            .in3(N__18561),
            .lcout(M_this_sprites_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36919),
            .ce(),
            .sr(N__32203));
    defparam M_this_sprites_address_q_RNO_0_8_LC_16_23_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_8_LC_16_23_7.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_8_LC_16_23_7.LUT_INIT=16'b1100110101000101;
    LogicCell40 M_this_sprites_address_q_RNO_0_8_LC_16_23_7 (
            .in0(N__26204),
            .in1(N__23510),
            .in2(N__26130),
            .in3(N__27051),
            .lcout(M_this_sprites_address_qc_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_LC_16_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_LC_16_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_LC_16_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__27054),
            .in2(_gnd_net_),
            .in3(N__31146),
            .lcout(\this_vga_signals.N_415_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_3_LC_16_27_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_3_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_3_LC_16_27_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_ram_write_data_0_a2_0_a4_3_LC_16_27_1  (
            .in0(N__35830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25266),
            .lcout(M_this_map_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_17_9_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_17_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19469),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36847),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI0VTU_0_4_LC_17_11_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI0VTU_0_4_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI0VTU_0_4_LC_17_11_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \this_ppu.M_state_q_RNI0VTU_0_4_LC_17_11_0  (
            .in0(N__18543),
            .in1(N__33773),
            .in2(N__18531),
            .in3(N__33863),
            .lcout(M_this_ppu_sprites_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIEH4G1_2_LC_17_11_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIEH4G1_2_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIEH4G1_2_LC_17_11_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIEH4G1_2_LC_17_11_7  (
            .in0(N__33772),
            .in1(N__27605),
            .in2(N__33888),
            .in3(N__19596),
            .lcout(M_this_ppu_sprites_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_17_12_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_17_12_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_17_12_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__19485),
            .in2(_gnd_net_),
            .in3(N__18123),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36852),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_17_12_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_17_12_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_17_12_4 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_17_12_4  (
            .in0(N__19484),
            .in1(N__18132),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36852),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIBD3G1_1_LC_17_13_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIBD3G1_1_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIBD3G1_1_LC_17_13_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIBD3G1_1_LC_17_13_1  (
            .in0(N__27713),
            .in1(N__33771),
            .in2(N__33846),
            .in3(N__19611),
            .lcout(M_this_ppu_sprites_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_17_14_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_17_14_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__19486),
            .in2(_gnd_net_),
            .in3(N__18675),
            .lcout(\this_reset_cond.M_stage_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36863),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_1_LC_17_14_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_17_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNO_0_1_LC_17_14_3  (
            .in0(N__20686),
            .in1(N__18944),
            .in2(N__33845),
            .in3(N__36097),
            .lcout(),
            .ltout(\this_ppu.M_state_q_srsts_i_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_1_LC_17_14_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_17_14_4 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \this_ppu.M_state_q_1_LC_17_14_4  (
            .in0(N__20646),
            .in1(N__19740),
            .in2(N__18666),
            .in3(N__18857),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36863),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIEF0G_7_LC_17_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIEF0G_7_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIEF0G_7_LC_17_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNIEF0G_7_LC_17_15_6  (
            .in0(N__18661),
            .in1(N__18605),
            .in2(N__18645),
            .in3(N__18582),
            .lcout(\this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5 ),
            .ltout(\this_ppu.M_count_d_0_sqmuxa_1_0_a3_7_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_2_LC_17_15_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_2_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_2_LC_17_15_7 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \this_ppu.M_state_q_2_LC_17_15_7  (
            .in0(N__18945),
            .in1(N__18906),
            .in2(N__18618),
            .in3(N__36103),
            .lcout(\this_ppu.M_state_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36870),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_1_LC_17_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_1_LC_17_16_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_1_LC_17_16_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_vaddress_q_1_LC_17_16_2  (
            .in0(N__27788),
            .in1(N__19683),
            .in2(N__27715),
            .in3(N__18856),
            .lcout(\this_ppu.M_vaddress_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36876),
            .ce(),
            .sr(N__21484));
    defparam \this_ppu.M_vaddress_q_0_LC_17_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_0_LC_17_16_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_0_LC_17_16_5 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \this_ppu.M_vaddress_q_0_LC_17_16_5  (
            .in0(N__19715),
            .in1(N__27787),
            .in2(N__19688),
            .in3(N__19905),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36876),
            .ce(),
            .sr(N__21484));
    defparam \this_ppu.M_count_q_5_LC_17_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_5_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_5_LC_17_17_0 .LUT_INIT=16'b1000100010000010;
    LogicCell40 \this_ppu.M_count_q_5_LC_17_17_0  (
            .in0(N__18827),
            .in1(N__18604),
            .in2(N__18615),
            .in3(N__18786),
            .lcout(\this_ppu.M_count_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36885),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_0_LC_17_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_0_LC_17_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_0_LC_17_17_1 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \this_ppu.M_count_q_0_LC_17_17_1  (
            .in0(N__18581),
            .in1(N__18777),
            .in2(_gnd_net_),
            .in3(N__18826),
            .lcout(\this_ppu.M_count_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36885),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_9_LC_17_17_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_9_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_9_LC_17_17_2 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \this_reset_cond.M_stage_q_9_LC_17_17_2  (
            .in0(N__18957),
            .in1(_gnd_net_),
            .in2(N__19509),
            .in3(_gnd_net_),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36885),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_8_LC_17_17_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_8_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_8_LC_17_17_3 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \this_reset_cond.M_stage_q_8_LC_17_17_3  (
            .in0(N__18681),
            .in1(N__19501),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36885),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIKRC91_1_LC_17_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIKRC91_1_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIKRC91_1_LC_17_17_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_state_q_RNIKRC91_1_LC_17_17_5  (
            .in0(N__18946),
            .in1(N__18915),
            .in2(_gnd_net_),
            .in3(N__18905),
            .lcout(\this_ppu.M_count_d_0_sqmuxa_1 ),
            .ltout(\this_ppu.M_count_d_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIN6OG6_0_LC_17_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIN6OG6_0_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIN6OG6_0_LC_17_17_6 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \this_ppu.M_state_q_RNIN6OG6_0_LC_17_17_6  (
            .in0(N__19670),
            .in1(N__29662),
            .in2(N__18864),
            .in3(N__18849),
            .lcout(\this_ppu.N_1417_0 ),
            .ltout(\this_ppu.N_1417_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_3_LC_17_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_3_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_3_LC_17_17_7 .LUT_INIT=16'b1100000010010000;
    LogicCell40 \this_ppu.M_count_q_3_LC_17_17_7  (
            .in0(N__18804),
            .in1(N__18751),
            .in2(N__18798),
            .in3(N__18778),
            .lcout(\this_ppu.M_count_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36885),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_6_LC_17_18_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_6_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_6_LC_17_18_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_6_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__19507),
            .in2(_gnd_net_),
            .in3(N__19434),
            .lcout(\this_reset_cond.M_stage_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36895),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_17_18_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_17_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_17_18_2  (
            .in0(N__28086),
            .in1(N__18729),
            .in2(_gnd_net_),
            .in3(N__18714),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_4_LC_17_18_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_4_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_4_LC_17_18_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_4_LC_17_18_3  (
            .in0(N__19505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18696),
            .lcout(\this_reset_cond.M_stage_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36895),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_7_LC_17_18_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_7_LC_17_18_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_7_LC_17_18_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_7_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__19508),
            .in2(_gnd_net_),
            .in3(N__18687),
            .lcout(\this_reset_cond.M_stage_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36895),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_5_LC_17_18_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_5_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_5_LC_17_18_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_5_LC_17_18_5  (
            .in0(N__19506),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19440),
            .lcout(\this_reset_cond.M_stage_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36895),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_17_19_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_17_19_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_17_19_0  (
            .in0(N__28068),
            .in1(N__19428),
            .in2(_gnd_net_),
            .in3(N__19410),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_11_LC_17_19_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_11_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_11_LC_17_19_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \this_sprites_ram.mem_radreg_11_LC_17_19_1  (
            .in0(N__33785),
            .in1(N__19395),
            .in2(N__19374),
            .in3(N__33906),
            .lcout(\this_sprites_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36899),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_13_LC_17_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_13_LC_17_19_3 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_13_LC_17_19_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \this_sprites_ram.mem_radreg_13_LC_17_19_3  (
            .in0(N__33786),
            .in1(N__19353),
            .in2(N__19335),
            .in3(N__33907),
            .lcout(\this_sprites_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36899),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_17_19_4  (
            .in0(N__28069),
            .in1(N__19311),
            .in2(_gnd_net_),
            .in3(N__19296),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_5 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_17_19_5  (
            .in0(N__21662),
            .in1(N__21757),
            .in2(N__19284),
            .in3(N__19281),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI0VTU_4_LC_17_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI0VTU_4_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI0VTU_4_LC_17_19_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \this_ppu.M_state_q_RNI0VTU_4_LC_17_19_6  (
            .in0(N__19275),
            .in1(N__19251),
            .in2(N__33927),
            .in3(N__33784),
            .lcout(M_this_ppu_sprites_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_17_19_7  (
            .in0(N__18990),
            .in1(N__18975),
            .in2(_gnd_net_),
            .in3(N__28070),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_LC_17_20_4.C_ON=1'b0;
    defparam M_this_substate_q_LC_17_20_4.SEQ_MODE=4'b1000;
    defparam M_this_substate_q_LC_17_20_4.LUT_INIT=16'b1111111110100010;
    LogicCell40 M_this_substate_q_LC_17_20_4 (
            .in0(N__31555),
            .in1(N__23377),
            .in2(N__19539),
            .in3(N__25533),
            .lcout(M_this_substate_qZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36906),
            .ce(),
            .sr(N__36018));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_480_LC_17_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_480_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_480_LC_17_21_0 .LUT_INIT=16'b0101010100000001;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_480_LC_17_21_0  (
            .in0(N__22128),
            .in1(N__24359),
            .in2(N__22203),
            .in3(N__26555),
            .lcout(),
            .ltout(M_this_sprites_address_q_0_0_i_480_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_4_LC_17_21_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_4_LC_17_21_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_4_LC_17_21_1.LUT_INIT=16'b0000110000000100;
    LogicCell40 M_this_sprites_address_q_4_LC_17_21_1 (
            .in0(N__19515),
            .in1(N__19527),
            .in2(N__19530),
            .in3(N__19521),
            .lcout(M_this_sprites_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36912),
            .ce(),
            .sr(N__32210));
    defparam M_this_sprites_address_q_RNO_0_4_LC_17_21_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_4_LC_17_21_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_4_LC_17_21_2.LUT_INIT=16'b1111000100110001;
    LogicCell40 M_this_sprites_address_q_RNO_0_4_LC_17_21_2 (
            .in0(N__24275),
            .in1(N__26216),
            .in2(N__22202),
            .in3(N__26413),
            .lcout(M_this_sprites_address_qc_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_4_LC_17_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_4_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_4_LC_17_21_3 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_4_LC_17_21_3  (
            .in0(N__25468),
            .in1(N__22127),
            .in2(_gnd_net_),
            .in3(N__27049),
            .lcout(N_511_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_4_LC_17_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_4_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_4_LC_17_21_4 .LUT_INIT=16'b0000010100001101;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_4_LC_17_21_4  (
            .in0(N__22170),
            .in1(N__31103),
            .in2(N__32441),
            .in3(N__26412),
            .lcout(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_5_LC_17_21_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_5_LC_17_21_6.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_5_LC_17_21_6.LUT_INIT=16'b0010001000000010;
    LogicCell40 M_this_sprites_address_q_5_LC_17_21_6 (
            .in0(N__20277),
            .in1(N__20349),
            .in2(N__19584),
            .in3(N__20283),
            .lcout(M_this_sprites_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36912),
            .ce(),
            .sr(N__32210));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_484_LC_17_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_484_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_484_LC_17_22_0 .LUT_INIT=16'b0000111100000001;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_484_LC_17_22_0  (
            .in0(N__22421),
            .in1(N__24358),
            .in2(N__22392),
            .in3(N__26537),
            .lcout(M_this_sprites_address_q_0_0_i_484),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_492_LC_17_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_492_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_492_LC_17_22_1 .LUT_INIT=16'b0000000010101011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_492_LC_17_22_1  (
            .in0(N__26536),
            .in1(N__22926),
            .in2(N__24367),
            .in3(N__22887),
            .lcout(M_this_sprites_address_q_0_0_i_492),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_3_LC_17_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_3_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_3_LC_17_22_2 .LUT_INIT=16'b0000010100001101;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_3_LC_17_22_2  (
            .in0(N__22422),
            .in1(N__31115),
            .in2(N__35831),
            .in3(N__26435),
            .lcout(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_5_LC_17_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_5_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_5_LC_17_22_3 .LUT_INIT=16'b0000011100000011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_5_LC_17_22_3  (
            .in0(N__26434),
            .in1(N__21919),
            .in2(N__36356),
            .in3(N__31117),
            .lcout(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_i_0_0_a4_4_LC_17_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_0_0_a4_4_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_0_0_a4_4_LC_17_22_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_0_0_a4_4_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(N__31178),
            .in2(_gnd_net_),
            .in3(N__31116),
            .lcout(),
            .ltout(\this_vga_signals.N_659_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_17_22_5.C_ON=1'b0;
    defparam M_this_state_q_4_LC_17_22_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_17_22_5.LUT_INIT=16'b1111100011110000;
    LogicCell40 M_this_state_q_4_LC_17_22_5 (
            .in0(N__25829),
            .in1(N__25744),
            .in2(N__19575),
            .in3(N__27073),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36922),
            .ce(),
            .sr(N__36023));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_2_LC_17_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_2_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_2_LC_17_23_0 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_2_LC_17_23_0  (
            .in0(N__25505),
            .in1(N__22625),
            .in2(N__19563),
            .in3(N__27053),
            .lcout(),
            .ltout(N_572_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_2_LC_17_23_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_2_LC_17_23_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_2_LC_17_23_1.LUT_INIT=16'b0000111000000000;
    LogicCell40 M_this_sprites_address_q_2_LC_17_23_1 (
            .in0(N__22626),
            .in1(N__19626),
            .in2(N__19572),
            .in3(N__19569),
            .lcout(M_this_sprites_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36927),
            .ce(),
            .sr(N__32206));
    defparam M_this_sprites_address_q_RNO_0_2_LC_17_23_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_2_LC_17_23_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_2_LC_17_23_2.LUT_INIT=16'b1000100011001111;
    LogicCell40 M_this_sprites_address_q_RNO_0_2_LC_17_23_2 (
            .in0(N__26432),
            .in1(N__22691),
            .in2(N__24280),
            .in3(N__26206),
            .lcout(M_this_sprites_address_qc_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_2_LC_17_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_2_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_2_LC_17_23_3 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_2_LC_17_23_3  (
            .in0(N__31144),
            .in1(N__22703),
            .in2(N__35238),
            .in3(N__26431),
            .lcout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_3_LC_17_23_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_3_LC_17_23_6.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_3_LC_17_23_6.LUT_INIT=16'b1000100011001111;
    LogicCell40 M_this_sprites_address_q_RNO_0_3_LC_17_23_6 (
            .in0(N__26433),
            .in1(N__22420),
            .in2(N__24281),
            .in3(N__26207),
            .lcout(),
            .ltout(M_this_sprites_address_qc_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_3_LC_17_23_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_3_LC_17_23_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_3_LC_17_23_7.LUT_INIT=16'b0011000000010000;
    LogicCell40 M_this_sprites_address_q_3_LC_17_23_7 (
            .in0(N__19554),
            .in1(N__19548),
            .in2(N__19542),
            .in3(N__20403),
            .lcout(M_this_sprites_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36927),
            .ce(),
            .sr(N__32206));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_6_LC_17_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_6_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_6_LC_17_24_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_6_LC_17_24_0  (
            .in0(N__25663),
            .in1(N__25746),
            .in2(_gnd_net_),
            .in3(N__25803),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2_1_LC_17_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2_1_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2_1_LC_17_24_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a2_1_LC_17_24_4  (
            .in0(N__25662),
            .in1(N__31646),
            .in2(_gnd_net_),
            .in3(N__23382),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_488_tz_LC_17_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_488_tz_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_488_tz_LC_17_24_5 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_488_tz_LC_17_24_5  (
            .in0(N__24345),
            .in1(N__22690),
            .in2(_gnd_net_),
            .in3(N__26548),
            .lcout(N_1318_tz_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_10_LC_17_25_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_10_LC_17_25_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_10_LC_17_25_0.LUT_INIT=16'b1111000100110001;
    LogicCell40 M_this_sprites_address_q_RNO_0_10_LC_17_25_0 (
            .in0(N__26105),
            .in1(N__26217),
            .in2(N__24493),
            .in3(N__27045),
            .lcout(M_this_sprites_address_qc_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_11_LC_17_25_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_11_LC_17_25_6.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_11_LC_17_25_6.LUT_INIT=16'b1111000100110001;
    LogicCell40 M_this_sprites_address_q_RNO_0_11_LC_17_25_6 (
            .in0(N__26106),
            .in1(N__26218),
            .in2(N__34676),
            .in3(N__27046),
            .lcout(M_this_sprites_address_qc_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_18_11_0 .C_ON=1'b1;
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_0_c_inv_LC_18_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un2_vscroll_cry_0_c_inv_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__19617),
            .in2(N__27823),
            .in3(N__27868),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\this_ppu.un2_vscroll_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_18_11_1 .C_ON=1'b1;
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_18_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__19590),
            .in2(N__27720),
            .in3(N__19602),
            .lcout(\this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0 ),
            .ltout(),
            .carryin(\this_ppu.un2_vscroll_cry_0 ),
            .carryout(\this_ppu.un2_vscroll_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_18_11_2 .C_ON=1'b0;
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_18_11_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_18_11_2  (
            .in0(N__27539),
            .in1(N__27604),
            .in2(_gnd_net_),
            .in3(N__19599),
            .lcout(\this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_18_11_5 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_18_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27659),
            .lcout(M_this_oam_ram_read_data_i_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_0_LC_18_13_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_0_LC_18_13_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_0_LC_18_13_2 .LUT_INIT=16'b1100011011000011;
    LogicCell40 \this_ppu.M_haddress_q_0_LC_18_13_2  (
            .in0(N__33725),
            .in1(N__34267),
            .in2(N__20642),
            .in3(N__19842),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36864),
            .ce(),
            .sr(N__21068));
    defparam \this_ppu.M_state_q_RNIQKAOF_3_LC_18_14_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIQKAOF_3_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIQKAOF_3_LC_18_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_RNIQKAOF_3_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__20669),
            .in2(_gnd_net_),
            .in3(N__19841),
            .lcout(\this_ppu.N_124 ),
            .ltout(\this_ppu.N_124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_4_LC_18_14_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_4_LC_18_14_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_4_LC_18_14_1 .LUT_INIT=16'b0011000000110010;
    LogicCell40 \this_ppu.M_state_q_4_LC_18_14_1  (
            .in0(N__20687),
            .in1(N__29697),
            .in2(N__19734),
            .in3(N__24852),
            .lcout(\this_ppu.M_state_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36871),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_2_LC_18_15_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_2_LC_18_15_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_2_LC_18_15_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_vaddress_q_2_LC_18_15_5  (
            .in0(N__27789),
            .in1(N__27703),
            .in2(N__27602),
            .in3(N__21528),
            .lcout(\this_ppu.M_vaddress_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36877),
            .ce(),
            .sr(N__21494));
    defparam \this_ppu.M_vaddress_q_6_LC_18_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_6_LC_18_15_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_6_LC_18_15_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_vaddress_q_6_LC_18_15_6  (
            .in0(N__27249),
            .in1(N__27319),
            .in2(_gnd_net_),
            .in3(N__19727),
            .lcout(M_this_ppu_map_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36877),
            .ce(),
            .sr(N__21494));
    defparam \this_ppu.M_vaddress_q_RNI3FOP5_4_LC_18_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI3FOP5_4_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI3FOP5_4_LC_18_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNI3FOP5_4_LC_18_16_0  (
            .in0(N__27461),
            .in1(N__27399),
            .in2(N__27606),
            .in3(N__20620),
            .lcout(\this_ppu.un1_M_vaddress_q_2_c5 ),
            .ltout(\this_ppu.un1_M_vaddress_q_2_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_5_LC_18_16_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_5_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_5_LC_18_16_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_ppu.M_vaddress_q_5_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19731),
            .in3(N__27317),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36886),
            .ce(),
            .sr(N__21474));
    defparam \this_ppu.M_vaddress_q_7_LC_18_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_7_LC_18_16_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_7_LC_18_16_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_vaddress_q_7_LC_18_16_3  (
            .in0(N__27250),
            .in1(N__27318),
            .in2(N__27958),
            .in3(N__19728),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36886),
            .ce(),
            .sr(N__21474));
    defparam \this_ppu.M_vaddress_q_3_LC_18_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_3_LC_18_16_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_3_LC_18_16_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_ppu.M_vaddress_q_3_LC_18_16_5  (
            .in0(N__20621),
            .in1(N__27601),
            .in2(_gnd_net_),
            .in3(N__27462),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36886),
            .ce(),
            .sr(N__21474));
    defparam \this_ppu.line_clk.M_last_q_RNI3BB75_LC_18_16_6 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI3BB75_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI3BB75_LC_18_16_6 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI3BB75_LC_18_16_6  (
            .in0(N__19716),
            .in1(N__36098),
            .in2(N__19689),
            .in3(N__19904),
            .lcout(\this_ppu.M_last_q_RNI3BB75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_17_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_18_17_1  (
            .in0(N__28094),
            .in1(N__19881),
            .in2(_gnd_net_),
            .in3(N__19860),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vram_en_i_a2_0_LC_18_17_3 .C_ON=1'b0;
    defparam \this_ppu.vram_en_i_a2_0_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vram_en_i_a2_0_LC_18_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.vram_en_i_a2_0_LC_18_17_3  (
            .in0(N__19796),
            .in1(N__21716),
            .in2(N__20006),
            .in3(N__19751),
            .lcout(\this_ppu.vram_en_i_a2Z0Z_0 ),
            .ltout(\this_ppu.vram_en_i_a2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIUTM1G_3_LC_18_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIUTM1G_3_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIUTM1G_3_LC_18_17_4 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \this_ppu.M_state_q_RNIUTM1G_3_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__33760),
            .in2(N__19824),
            .in3(N__20670),
            .lcout(M_this_ppu_vram_en_0),
            .ltout(M_this_ppu_vram_en_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNINDU1G_1_LC_18_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNINDU1G_1_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNINDU1G_1_LC_18_17_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNINDU1G_1_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__33031),
            .in2(N__19821),
            .in3(N__34283),
            .lcout(\this_ppu.un1_M_haddress_q_3_c2 ),
            .ltout(\this_ppu.un1_M_haddress_q_3_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI4T92G_4_LC_18_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI4T92G_4_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI4T92G_4_LC_18_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNI4T92G_4_LC_18_17_6  (
            .in0(N__21416),
            .in1(N__21334),
            .in2(N__19818),
            .in3(N__32743),
            .lcout(\this_ppu.un1_M_haddress_q_3_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_18_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_18_0 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_18_18_0  (
            .in0(N__19815),
            .in1(N__20235),
            .in2(N__21766),
            .in3(N__19809),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_18_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_18_4 .LUT_INIT=16'b0000101101011011;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_18_18_4  (
            .in0(N__21753),
            .in1(N__19785),
            .in2(N__21666),
            .in3(N__19779),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_18_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_18_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_18_18_5  (
            .in0(N__21765),
            .in1(N__19773),
            .in2(N__19761),
            .in3(N__28020),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_18_19_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_18_19_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_18_19_0  (
            .in0(N__28088),
            .in1(N__20268),
            .in2(_gnd_net_),
            .in3(N__20250),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIITVO4_0_7_LC_18_19_1.C_ON=1'b0;
    defparam M_this_state_q_RNIITVO4_0_7_LC_18_19_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIITVO4_0_7_LC_18_19_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 M_this_state_q_RNIITVO4_0_7_LC_18_19_1 (
            .in0(N__24951),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dma_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_19_2  (
            .in0(N__28087),
            .in1(N__20052),
            .in2(_gnd_net_),
            .in3(N__20037),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_18_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_18_19_3 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_18_19_3  (
            .in0(N__21661),
            .in1(N__21763),
            .in2(N__20019),
            .in3(N__21831),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_18_19_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_18_19_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_18_19_4  (
            .in0(N__21764),
            .in1(N__19911),
            .in2(N__20016),
            .in3(N__19950),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_18_19_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_18_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_18_19_6  (
            .in0(N__28089),
            .in1(N__19983),
            .in2(_gnd_net_),
            .in3(N__19965),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_18_19_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_18_19_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_18_19_7  (
            .in0(N__19944),
            .in1(N__19929),
            .in2(_gnd_net_),
            .in3(N__28090),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_9_LC_18_20_0.C_ON=1'b0;
    defparam M_this_state_q_9_LC_18_20_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_18_20_0.LUT_INIT=16'b0000000011100000;
    LogicCell40 M_this_state_q_9_LC_18_20_0 (
            .in0(N__25047),
            .in1(N__25118),
            .in2(N__27180),
            .in3(N__25162),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36913),
            .ce(),
            .sr(N__36016));
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_0_LC_18_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_0_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_0_LC_18_20_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_19_i_0_o2_0_LC_18_20_1  (
            .in0(N__25119),
            .in1(N__25155),
            .in2(_gnd_net_),
            .in3(N__25046),
            .lcout(\this_vga_signals.N_419_0 ),
            .ltout(\this_vga_signals.N_419_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_LC_18_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_LC_18_20_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_19_i_0_o2_LC_18_20_2  (
            .in0(N__25599),
            .in1(N__25568),
            .in2(N__20313),
            .in3(N__35253),
            .lcout(N_440_0),
            .ltout(N_440_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o4_0_LC_18_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o4_0_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o4_0_LC_18_20_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_19_i_0_o4_0_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20310),
            .in3(N__31639),
            .lcout(\this_vga_signals.N_467_0 ),
            .ltout(\this_vga_signals.N_467_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_18_20_4.C_ON=1'b0;
    defparam M_this_state_q_5_LC_18_20_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_18_20_4.LUT_INIT=16'b1010000011101100;
    LogicCell40 M_this_state_q_5_LC_18_20_4 (
            .in0(N__20385),
            .in1(N__28192),
            .in2(N__20307),
            .in3(N__31126),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36913),
            .ce(),
            .sr(N__36016));
    defparam M_this_state_q_6_LC_18_20_5.C_ON=1'b0;
    defparam M_this_state_q_6_LC_18_20_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_18_20_5.LUT_INIT=16'b1101010111000000;
    LogicCell40 M_this_state_q_6_LC_18_20_5 (
            .in0(N__31125),
            .in1(N__20304),
            .in2(N__20298),
            .in3(N__29316),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36913),
            .ce(),
            .sr(N__36016));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_7_LC_18_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_7_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_7_LC_18_20_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_7_LC_18_20_6  (
            .in0(N__29315),
            .in1(N__30404),
            .in2(_gnd_net_),
            .in3(N__26241),
            .lcout(\this_vga_signals.N_732 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o4_LC_18_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o4_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o4_LC_18_21_0 .LUT_INIT=16'b0011001111101110;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_19_i_0_o4_LC_18_21_0  (
            .in0(N__25815),
            .in1(N__25664),
            .in2(_gnd_net_),
            .in3(N__25745),
            .lcout(\this_vga_signals.N_459_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_5_LC_18_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_5_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_5_LC_18_21_1 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_5_LC_18_21_1  (
            .in0(N__25483),
            .in1(N__21884),
            .in2(_gnd_net_),
            .in3(N__27048),
            .lcout(N_510_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_5_LC_18_21_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_5_LC_18_21_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_5_LC_18_21_2.LUT_INIT=16'b1111000100110001;
    LogicCell40 M_this_sprites_address_q_RNO_0_5_LC_18_21_2 (
            .in0(N__24268),
            .in1(N__26214),
            .in2(N__21936),
            .in3(N__26403),
            .lcout(M_this_sprites_address_qc_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0Z0Z_0_LC_18_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0Z0Z_0_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0Z0Z_0_LC_18_21_3 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0Z0Z_0_LC_18_21_3  (
            .in0(N__25482),
            .in1(N__23123),
            .in2(N__20334),
            .in3(N__27047),
            .lcout(),
            .ltout(N_562_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_0_LC_18_21_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_0_LC_18_21_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_0_LC_18_21_4.LUT_INIT=16'b0000101100000011;
    LogicCell40 M_this_sprites_address_q_RNO_0_0_LC_18_21_4 (
            .in0(N__23184),
            .in1(N__26215),
            .in2(N__20352),
            .in3(N__26404),
            .lcout(M_this_sprites_address_qc_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_476_LC_18_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_476_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_476_LC_18_21_5 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_476_LC_18_21_5  (
            .in0(N__21935),
            .in1(N__21885),
            .in2(N__24368),
            .in3(N__26554),
            .lcout(M_this_sprites_address_q_0_0_i_476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_496_LC_18_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_496_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_496_LC_18_22_0 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_496_LC_18_22_0  (
            .in0(N__23183),
            .in1(N__23127),
            .in2(N__24369),
            .in3(N__26538),
            .lcout(),
            .ltout(M_this_sprites_address_q_0_0_i_496_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_0_LC_18_22_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_0_LC_18_22_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_0_LC_18_22_1.LUT_INIT=16'b0000101100000000;
    LogicCell40 M_this_sprites_address_q_0_LC_18_22_1 (
            .in0(N__23185),
            .in1(N__24279),
            .in2(N__20343),
            .in3(N__20340),
            .lcout(M_this_sprites_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36928),
            .ce(),
            .sr(N__32211));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_0_LC_18_22_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_0_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_0_LC_18_22_4 .LUT_INIT=16'b0000010100001101;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_0_LC_18_22_4  (
            .in0(N__23182),
            .in1(N__31111),
            .in2(N__31355),
            .in3(N__26417),
            .lcout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_0_LC_18_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_0_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_0_LC_18_22_5 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_0_LC_18_22_5  (
            .in0(N__26416),
            .in1(N__25472),
            .in2(N__31143),
            .in3(N__27043),
            .lcout(N_773),
            .ltout(N_773_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_1_LC_18_22_6.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_1_LC_18_22_6.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_1_LC_18_22_6.LUT_INIT=16'b1010101100100011;
    LogicCell40 M_this_sprites_address_q_RNO_0_1_LC_18_22_6 (
            .in0(N__22925),
            .in1(N__26219),
            .in2(N__20325),
            .in3(N__26418),
            .lcout(),
            .ltout(M_this_sprites_address_qc_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_1_LC_18_22_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_1_LC_18_22_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_1_LC_18_22_7.LUT_INIT=16'b0011000000010000;
    LogicCell40 M_this_sprites_address_q_1_LC_18_22_7 (
            .in0(N__20370),
            .in1(N__20322),
            .in2(N__20316),
            .in3(N__20409),
            .lcout(M_this_sprites_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36928),
            .ce(),
            .sr(N__32211));
    defparam M_this_sprites_address_q_13_LC_18_23_0.C_ON=1'b0;
    defparam M_this_sprites_address_q_13_LC_18_23_0.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_13_LC_18_23_0.LUT_INIT=16'b0000000010101000;
    LogicCell40 M_this_sprites_address_q_13_LC_18_23_0 (
            .in0(N__26253),
            .in1(N__23400),
            .in2(N__26268),
            .in3(N__24378),
            .lcout(M_this_sprites_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36931),
            .ce(),
            .sr(N__32208));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_13_LC_18_23_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_13_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_13_LC_18_23_2 .LUT_INIT=16'b0000011100000101;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_13_LC_18_23_2  (
            .in0(N__34771),
            .in1(N__27006),
            .in2(N__34439),
            .in3(N__31120),
            .lcout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_1_LC_18_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_1_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_1_LC_18_23_3 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_1_LC_18_23_3  (
            .in0(N__25498),
            .in1(N__22883),
            .in2(_gnd_net_),
            .in3(N__27017),
            .lcout(N_896_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_3_LC_18_23_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_3_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_3_LC_18_23_4 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_3_LC_18_23_4  (
            .in0(N__25484),
            .in1(N__22385),
            .in2(_gnd_net_),
            .in3(N__27007),
            .lcout(N_512_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_8_LC_18_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_8_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_8_LC_18_23_7 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_8_LC_18_23_7  (
            .in0(N__31121),
            .in1(N__23518),
            .in2(N__33372),
            .in3(N__27016),
            .lcout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_5_LC_18_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_5_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_5_LC_18_24_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_5_LC_18_24_1  (
            .in0(N__25743),
            .in1(N__25649),
            .in2(_gnd_net_),
            .in3(N__25828),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_11_LC_18_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_11_LC_18_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_11_LC_18_24_4 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_11_LC_18_24_4  (
            .in0(N__31122),
            .in1(N__34651),
            .in2(N__32426),
            .in3(N__27044),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_11_LC_18_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_11_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_11_LC_18_24_5 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_11_LC_18_24_5  (
            .in0(N__26420),
            .in1(N__25501),
            .in2(N__20373),
            .in3(N__23444),
            .lcout(N_617),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_1_LC_18_24_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_1_LC_18_24_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_1_LC_18_24_7 .LUT_INIT=16'b0000011100000011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_1_LC_18_24_7  (
            .in0(N__26419),
            .in1(N__22947),
            .in2(N__33360),
            .in3(N__31123),
            .lcout(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_456_tz_LC_18_25_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_456_tz_LC_18_25_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_456_tz_LC_18_25_0 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_456_tz_LC_18_25_0  (
            .in0(N__26415),
            .in1(N__24459),
            .in2(N__31145),
            .in3(N__26556),
            .lcout(),
            .ltout(N_1286_tz_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_10_LC_18_25_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_10_LC_18_25_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_10_LC_18_25_1.LUT_INIT=16'b0010001000100000;
    LogicCell40 M_this_sprites_address_q_10_LC_18_25_1 (
            .in0(N__20361),
            .in1(N__24396),
            .in2(N__20355),
            .in3(N__24414),
            .lcout(M_this_sprites_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36941),
            .ce(),
            .sr(N__32204));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_7_LC_18_25_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_7_LC_18_25_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_7_LC_18_25_5 .LUT_INIT=16'b0011000010100000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_7_LC_18_25_5  (
            .in0(N__27038),
            .in1(N__31127),
            .in2(N__25499),
            .in3(N__26414),
            .lcout(N_762),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_11_LC_18_25_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_11_LC_18_25_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_11_LC_18_25_7.LUT_INIT=16'b0100010001000000;
    LogicCell40 M_this_sprites_address_q_11_LC_18_25_7 (
            .in0(N__20421),
            .in1(N__20415),
            .in2(N__24003),
            .in3(N__23448),
            .lcout(M_this_sprites_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36941),
            .ce(),
            .sr(N__32204));
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_5_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_5_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_5_0  (
            .in0(_gnd_net_),
            .in1(N__32798),
            .in2(N__20535),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_5_0_),
            .carryout(\this_ppu.un1_M_haddress_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_5_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_5_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_5_1  (
            .in0(_gnd_net_),
            .in1(N__20514),
            .in2(N__32000),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_0 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_5_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_5_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_5_2  (
            .in0(_gnd_net_),
            .in1(N__20496),
            .in2(N__33130),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_1 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_5_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_5_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_5_3  (
            .in0(_gnd_net_),
            .in1(N__31811),
            .in2(N__20481),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_2 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_5_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_5_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_5_4  (
            .in0(_gnd_net_),
            .in1(N__31839),
            .in2(N__20460),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_3 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_5_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_5_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_5_5  (
            .in0(_gnd_net_),
            .in1(N__31743),
            .in2(N__20442),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_4 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_5_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_5_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_5_6  (
            .in0(_gnd_net_),
            .in1(N__31770),
            .in2(N__20739),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_5 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_5_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_5_7  (
            .in0(_gnd_net_),
            .in1(N__31875),
            .in2(N__20718),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_cry_6 ),
            .carryout(\this_ppu.un1_M_haddress_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_cry_7_THRU_LUT4_0_LC_19_6_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_haddress_q_cry_7_THRU_LUT4_0_LC_19_6_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_cry_7_THRU_LUT4_0_LC_19_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_cry_7_THRU_LUT4_0_LC_19_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20538),
            .lcout(\this_ppu.un1_M_haddress_q_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_19_7_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_19_7_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_19_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_19_7_0  (
            .in0(_gnd_net_),
            .in1(N__32799),
            .in2(N__20531),
            .in3(N__34297),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_0 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_19_7_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_19_7_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_19_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_19_7_1  (
            .in0(_gnd_net_),
            .in1(N__32001),
            .in2(N__20513),
            .in3(N__33060),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_0 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_19_7_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_19_7_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_19_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(N__20492),
            .in2(N__33135),
            .in3(N__32720),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_1 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_19_7_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_19_7_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_19_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(N__24825),
            .in2(N__20477),
            .in3(N__21361),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_0 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_2 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_19_7_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_19_7_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_19_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(N__20453),
            .in2(N__24390),
            .in3(N__21424),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_3 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_19_7_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_19_7_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_19_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_19_7_5  (
            .in0(_gnd_net_),
            .in1(N__31902),
            .in2(N__20438),
            .in3(N__21235),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_4 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_19_7_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_19_7_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_19_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_19_7_6  (
            .in0(_gnd_net_),
            .in1(N__31722),
            .in2(N__20735),
            .in3(N__21160),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_3 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_5 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_19_7_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_19_7_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_19_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_19_7_7  (
            .in0(N__21290),
            .in1(N__31854),
            .in2(N__20714),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_4 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_haddress_q_2_cry_6 ),
            .carryout(\this_ppu.un1_M_haddress_q_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_THRU_LUT4_0_LC_19_8_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_THRU_LUT4_0_LC_19_8_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_THRU_LUT4_0_LC_19_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_7_THRU_LUT4_0_LC_19_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20697),
            .lcout(\this_ppu.un1_M_haddress_q_2_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_5_LC_19_9_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_5_LC_19_9_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_5_LC_19_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_5_LC_19_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36355),
            .lcout(M_this_data_tmp_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36849),
            .ce(N__30229),
            .sr(N__36027));
    defparam \this_ppu.M_state_q_3_LC_19_12_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_3_LC_19_12_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_3_LC_19_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_state_q_3_LC_19_12_5  (
            .in0(N__20694),
            .in1(N__36105),
            .in2(_gnd_net_),
            .in3(N__24848),
            .lcout(\this_ppu.M_state_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36865),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI6GOI_3_LC_19_13_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI6GOI_3_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI6GOI_3_LC_19_13_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_state_q_RNI6GOI_3_LC_19_13_1  (
            .in0(_gnd_net_),
            .in1(N__33713),
            .in2(_gnd_net_),
            .in3(N__20665),
            .lcout(\this_ppu.N_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_5_LC_19_13_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_5_LC_19_13_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_5_LC_19_13_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_5_LC_19_13_6  (
            .in0(_gnd_net_),
            .in1(N__33844),
            .in2(_gnd_net_),
            .in3(N__36104),
            .lcout(\this_ppu.M_state_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36872),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_4_LC_19_14_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_4_LC_19_14_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_4_LC_19_14_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_vaddress_q_4_LC_19_14_6  (
            .in0(N__27472),
            .in1(N__27585),
            .in2(N__27400),
            .in3(N__20625),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36878),
            .ce(),
            .sr(N__21495));
    defparam \this_ppu.M_haddress_q_2_LC_19_15_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_2_LC_19_15_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_2_LC_19_15_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_haddress_q_2_LC_19_15_3  (
            .in0(N__33039),
            .in1(N__34290),
            .in2(N__32737),
            .in3(N__21092),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36887),
            .ce(),
            .sr(N__21067));
    defparam \this_ppu.line_clk.M_last_q_RNIQRTEB_LC_19_16_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIQRTEB_LC_19_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIQRTEB_LC_19_16_3 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIQRTEB_LC_19_16_3  (
            .in0(N__20585),
            .in1(N__29700),
            .in2(N__24939),
            .in3(N__21524),
            .lcout(\this_ppu.M_last_q_RNIQRTEB ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_4_LC_19_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_4_LC_19_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_4_LC_19_17_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \this_ppu.M_haddress_q_4_LC_19_17_0  (
            .in0(N__21384),
            .in1(N__21336),
            .in2(N__32738),
            .in3(N__21417),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36900),
            .ce(),
            .sr(N__21069));
    defparam \this_ppu.M_haddress_q_3_LC_19_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_3_LC_19_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_3_LC_19_17_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_3_LC_19_17_1  (
            .in0(N__21335),
            .in1(N__32721),
            .in2(_gnd_net_),
            .in3(N__21383),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36900),
            .ce(),
            .sr(N__21069));
    defparam \this_ppu.M_haddress_q_7_LC_19_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_7_LC_19_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_7_LC_19_17_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_haddress_q_7_LC_19_17_2  (
            .in0(N__21258),
            .in1(N__21280),
            .in2(N__21219),
            .in3(N__21135),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36900),
            .ce(),
            .sr(N__21069));
    defparam \this_ppu.M_haddress_q_5_LC_19_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_5_LC_19_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_5_LC_19_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_haddress_q_5_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__21202),
            .in2(_gnd_net_),
            .in3(N__21256),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36900),
            .ce(),
            .sr(N__21069));
    defparam \this_ppu.M_haddress_q_6_LC_19_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_6_LC_19_17_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_6_LC_19_17_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_ppu.M_haddress_q_6_LC_19_17_4  (
            .in0(N__21257),
            .in1(_gnd_net_),
            .in2(N__21218),
            .in3(N__21134),
            .lcout(M_this_ppu_map_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36900),
            .ce(),
            .sr(N__21069));
    defparam \this_ppu.M_haddress_q_1_LC_19_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_1_LC_19_17_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_1_LC_19_17_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_1_LC_19_17_7  (
            .in0(N__33032),
            .in1(N__34303),
            .in2(_gnd_net_),
            .in3(N__21085),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36900),
            .ce(),
            .sr(N__21069));
    defparam M_this_state_q_fast_9_LC_19_18_4.C_ON=1'b0;
    defparam M_this_state_q_fast_9_LC_19_18_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_fast_9_LC_19_18_4.LUT_INIT=16'b0010001000100000;
    LogicCell40 M_this_state_q_fast_9_LC_19_18_4 (
            .in0(N__27179),
            .in1(N__25164),
            .in2(N__25117),
            .in3(N__25056),
            .lcout(M_this_state_q_fastZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36907),
            .ce(),
            .sr(N__36008));
    defparam \this_ppu.M_state_q_RNI0VTU_1_4_LC_19_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI0VTU_1_4_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI0VTU_1_4_LC_19_19_0 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_ppu.M_state_q_RNI0VTU_1_4_LC_19_19_0  (
            .in0(N__33776),
            .in1(N__21036),
            .in2(N__33934),
            .in3(N__21015),
            .lcout(M_this_ppu_sprites_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_19_19_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_19_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_19_19_1  (
            .in0(N__28096),
            .in1(N__21807),
            .in2(_gnd_net_),
            .in3(N__21789),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_19_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_19_19_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_19_19_2  (
            .in0(N__21660),
            .in1(N__21767),
            .in2(N__21771),
            .in3(N__21609),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_19_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_19_19_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_19_19_3  (
            .in0(N__21768),
            .in1(N__21534),
            .in2(N__21723),
            .in3(N__21567),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_12_LC_19_19_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_12_LC_19_19_4 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_12_LC_19_19_4 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \this_sprites_ram.mem_radreg_12_LC_19_19_4  (
            .in0(N__33777),
            .in1(N__21699),
            .in2(N__33935),
            .in3(N__21684),
            .lcout(\this_sprites_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36914),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_19_19_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_19_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_19_19_5  (
            .in0(N__28095),
            .in1(N__21633),
            .in2(_gnd_net_),
            .in3(N__21618),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_19_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_19_19_6  (
            .in0(N__21603),
            .in1(N__21585),
            .in2(_gnd_net_),
            .in3(N__28097),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_19_19_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_19_19_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_19_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_19_19_7  (
            .in0(N__28098),
            .in1(N__21561),
            .in2(_gnd_net_),
            .in3(N__21552),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_9_LC_19_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_9_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_9_LC_19_20_1 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_9_LC_19_20_1  (
            .in0(N__30945),
            .in1(N__25951),
            .in2(N__35224),
            .in3(N__27042),
            .lcout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_tr30_0_0_a2_0_a2_LC_19_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_tr30_0_0_a2_0_a2_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_tr30_0_0_a2_0_a2_LC_19_20_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_vga_signals.M_this_state_q_tr30_0_0_a2_0_a2_LC_19_20_3  (
            .in0(N__30944),
            .in1(_gnd_net_),
            .in2(N__29376),
            .in3(_gnd_net_),
            .lcout(M_this_map_ram_write_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_19_20_4 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_19_20_4 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_19_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_19_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21870),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36923),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_20_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_20_5  (
            .in0(N__28108),
            .in1(N__21861),
            .in2(_gnd_net_),
            .in3(N__21846),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_m2_LC_19_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_m2_LC_19_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_m2_LC_19_20_6 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_6_0_0_m2_LC_19_20_6  (
            .in0(N__26240),
            .in1(N__26518),
            .in2(N__30416),
            .in3(N__30943),
            .lcout(\this_vga_signals.N_505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_19_20_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_19_20_7 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_19_20_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_19_20_7  (
            .in0(N__25108),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25054),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36923),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2_0_LC_19_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2_0_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2_0_LC_19_21_0 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_i_a4_2_0_LC_19_21_0  (
            .in0(N__31624),
            .in1(N__29299),
            .in2(N__25173),
            .in3(N__27125),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_i_a4_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_0_i_a2_9_LC_19_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_0_i_a2_9_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_0_i_a2_9_LC_19_21_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_0_i_a2_9_LC_19_21_1  (
            .in0(N__29297),
            .in1(N__35229),
            .in2(N__26787),
            .in3(N__30946),
            .lcout(\this_vga_signals.N_746 ),
            .ltout(\this_vga_signals.N_746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_i_LC_19_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_i_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_i_LC_19_21_2 .LUT_INIT=16'b0101000001110011;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_6_0_0_i_LC_19_21_2  (
            .in0(N__36325),
            .in1(N__29298),
            .in2(N__21825),
            .in3(N__21822),
            .lcout(un1_M_this_state_q_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4_0_LC_19_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4_0_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4_0_LC_19_21_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_i_a4_4_0_LC_19_21_3  (
            .in0(N__31213),
            .in1(N__28191),
            .in2(N__21816),
            .in3(N__26509),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_i_a4_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_3_LC_19_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_3_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_3_LC_19_21_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_3_LC_19_21_4  (
            .in0(N__30948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27126),
            .lcout(\this_vga_signals.N_648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_1_0_LC_19_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_1_0_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_1_0_LC_19_21_5 .LUT_INIT=16'b0000000011010101;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_i_1_0_LC_19_21_5  (
            .in0(N__31625),
            .in1(N__23388),
            .in2(N__23381),
            .in3(N__30947),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_i_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNIRO0N6_0_LC_19_22_0.C_ON=1'b1;
    defparam M_this_sprites_address_q_RNIRO0N6_0_LC_19_22_0.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNIRO0N6_0_LC_19_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_sprites_address_q_RNIRO0N6_0_LC_19_22_0 (
            .in0(_gnd_net_),
            .in1(N__23181),
            .in2(N__23142),
            .in3(N__23141),
            .lcout(M_this_sprites_address_q_RNIRO0N6Z0Z_0),
            .ltout(),
            .carryin(bfn_19_22_0_),
            .carryout(un1_M_this_sprites_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_0_c_RNIUIDH_LC_19_22_1 (
            .in0(_gnd_net_),
            .in1(N__22924),
            .in2(_gnd_net_),
            .in3(N__22872),
            .lcout(un1_M_this_sprites_address_q_cry_0_c_RNIUIDHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_0),
            .carryout(un1_M_this_sprites_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_sprites_address_q_cry_1_c_RNI0MEH_LC_19_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22775),
            .in3(N__22611),
            .lcout(un1_M_this_sprites_address_q_cry_1_c_RNI0MEHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_1),
            .carryout(un1_M_this_sprites_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_2_c_RNI2PFH_LC_19_22_3 (
            .in0(_gnd_net_),
            .in1(N__22448),
            .in2(_gnd_net_),
            .in3(N__22371),
            .lcout(un1_M_this_sprites_address_q_cry_2_c_RNI2PFHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_2),
            .carryout(un1_M_this_sprites_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_3_c_RNI4SGH_LC_19_22_4 (
            .in0(_gnd_net_),
            .in1(N__22204),
            .in2(_gnd_net_),
            .in3(N__22113),
            .lcout(un1_M_this_sprites_address_q_cry_3_c_RNI4SGHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_3),
            .carryout(un1_M_this_sprites_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_4_c_RNI6VHH_LC_19_22_5 (
            .in0(_gnd_net_),
            .in1(N__21947),
            .in2(_gnd_net_),
            .in3(N__21876),
            .lcout(un1_M_this_sprites_address_q_cry_4_c_RNI6VHHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_4),
            .carryout(un1_M_this_sprites_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_5_c_RNI82JH_LC_19_22_6 (
            .in0(_gnd_net_),
            .in1(N__24071),
            .in2(_gnd_net_),
            .in3(N__21873),
            .lcout(un1_M_this_sprites_address_q_cry_5_c_RNI82JHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_5),
            .carryout(un1_M_this_sprites_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_6_c_RNIA5KH_LC_19_22_7 (
            .in0(_gnd_net_),
            .in1(N__23811),
            .in2(_gnd_net_),
            .in3(N__23691),
            .lcout(un1_M_this_sprites_address_q_cry_6_c_RNIA5KHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_6),
            .carryout(un1_M_this_sprites_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_7_c_RNIC8LH_LC_19_23_0 (
            .in0(_gnd_net_),
            .in1(N__23517),
            .in2(_gnd_net_),
            .in3(N__23457),
            .lcout(un1_M_this_sprites_address_q_cry_7_c_RNIC8LHZ0),
            .ltout(),
            .carryin(bfn_19_23_0_),
            .carryout(un1_M_this_sprites_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_8_c_RNIEBMH_LC_19_23_1 (
            .in0(_gnd_net_),
            .in1(N__25875),
            .in2(_gnd_net_),
            .in3(N__23454),
            .lcout(un1_M_this_sprites_address_q_cry_8_c_RNIEBMHZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_8),
            .carryout(un1_M_this_sprites_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_9_c_RNIN4NQ_LC_19_23_2 (
            .in0(_gnd_net_),
            .in1(N__24492),
            .in2(_gnd_net_),
            .in3(N__23451),
            .lcout(un1_M_this_sprites_address_q_cry_9_c_RNIN4NQZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_9),
            .carryout(un1_M_this_sprites_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_10_c_RNI09GE_LC_19_23_3 (
            .in0(_gnd_net_),
            .in1(N__34675),
            .in2(_gnd_net_),
            .in3(N__23433),
            .lcout(un1_M_this_sprites_address_q_cry_10_c_RNI09GEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_10),
            .carryout(un1_M_this_sprites_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4.C_ON=1'b1;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_sprites_address_q_cry_11_c_RNI2CHE_LC_19_23_4 (
            .in0(_gnd_net_),
            .in1(N__34953),
            .in2(_gnd_net_),
            .in3(N__23430),
            .lcout(un1_M_this_sprites_address_q_cry_11_c_RNI2CHEZ0),
            .ltout(),
            .carryin(un1_M_this_sprites_address_q_cry_11),
            .carryout(un1_M_this_sprites_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5.C_ON=1'b0;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_M_this_sprites_address_q_cry_12_c_RNI4FIE_LC_19_23_5 (
            .in0(_gnd_net_),
            .in1(N__34748),
            .in2(_gnd_net_),
            .in3(N__23427),
            .lcout(un1_M_this_sprites_address_q_cry_12_c_RNI4FIEZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_9_LC_19_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_9_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_9_LC_19_23_6 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_9_LC_19_23_6  (
            .in0(N__26424),
            .in1(N__25486),
            .in2(N__23424),
            .in3(N__23990),
            .lcout(N_607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_13_LC_19_23_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_13_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_13_LC_19_23_7 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_13_LC_19_23_7  (
            .in0(N__25485),
            .in1(N__26425),
            .in2(N__23409),
            .in3(N__23399),
            .lcout(N_627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_6_LC_19_24_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_6_LC_19_24_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_6_LC_19_24_0 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_o2_0_6_LC_19_24_0  (
            .in0(N__26989),
            .in1(N__25502),
            .in2(_gnd_net_),
            .in3(N__24305),
            .lcout(),
            .ltout(N_509_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_6_LC_19_24_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_6_LC_19_24_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_6_LC_19_24_1.LUT_INIT=16'b0000000011000100;
    LogicCell40 M_this_sprites_address_q_6_LC_19_24_1 (
            .in0(N__24288),
            .in1(N__24009),
            .in2(N__24372),
            .in3(N__24294),
            .lcout(M_this_sprites_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36942),
            .ce(),
            .sr(N__32209));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_472_LC_19_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_472_LC_19_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_472_LC_19_24_2 .LUT_INIT=16'b0000000010101011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_472_LC_19_24_2  (
            .in0(N__26550),
            .in1(N__24366),
            .in2(N__24109),
            .in3(N__24306),
            .lcout(M_this_sprites_address_q_0_0_i_472),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_6_LC_19_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_6_LC_19_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_6_LC_19_24_3 .LUT_INIT=16'b0001001100000011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_6_LC_19_24_3  (
            .in0(N__26422),
            .in1(N__34445),
            .in2(N__24153),
            .in3(N__31105),
            .lcout(this_vga_signals_M_this_sprites_address_q_0_0_i_a4_0_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_6_LC_19_24_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_6_LC_19_24_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_6_LC_19_24_4.LUT_INIT=16'b1111010100010001;
    LogicCell40 M_this_sprites_address_q_RNO_0_6_LC_19_24_4 (
            .in0(N__26184),
            .in1(N__24282),
            .in2(N__26439),
            .in3(N__24108),
            .lcout(M_this_sprites_address_qc_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_452_tz_LC_19_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_452_tz_LC_19_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_452_tz_LC_19_24_5 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_452_tz_LC_19_24_5  (
            .in0(N__26421),
            .in1(N__31104),
            .in2(N__34677),
            .in3(N__26549),
            .lcout(N_1282_tz_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_460_tz_LC_19_24_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_460_tz_LC_19_24_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_460_tz_LC_19_24_6 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_460_tz_LC_19_24_6  (
            .in0(N__26551),
            .in1(N__31124),
            .in2(N__25953),
            .in3(N__26423),
            .lcout(),
            .ltout(N_1290_tz_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_9_LC_19_24_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_9_LC_19_24_7.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_9_LC_19_24_7.LUT_INIT=16'b0000000011001000;
    LogicCell40 M_this_sprites_address_q_9_LC_19_24_7 (
            .in0(N__23991),
            .in1(N__25839),
            .in2(N__23979),
            .in3(N__23976),
            .lcout(M_this_sprites_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36942),
            .ce(),
            .sr(N__32209));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_10_LC_19_25_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_10_LC_19_25_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_10_LC_19_25_6 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_10_LC_19_25_6  (
            .in0(N__31102),
            .in1(N__24455),
            .in2(N__35863),
            .in3(N__27005),
            .lcout(),
            .ltout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_10_LC_19_25_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_10_LC_19_25_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_10_LC_19_25_7 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_10_LC_19_25_7  (
            .in0(N__25500),
            .in1(N__24413),
            .in2(N__24399),
            .in3(N__26429),
            .lcout(N_612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_map_address_q_0_i_a4_9_LC_19_27_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_map_address_q_0_i_a4_9_LC_19_27_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_map_address_q_0_i_a4_9_LC_19_27_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_map_address_q_0_i_a4_9_LC_19_27_5  (
            .in0(N__36344),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31706),
            .lcout(N_560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_20_5_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_20_5_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc1_LC_20_5_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc1_LC_20_5_1  (
            .in0(_gnd_net_),
            .in1(N__31838),
            .in2(_gnd_net_),
            .in3(N__31810),
            .lcout(\this_ppu.un1_M_haddress_q_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_6_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_6_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_6_0  (
            .in0(_gnd_net_),
            .in1(N__27870),
            .in2(N__27738),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_6_0_),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_6_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_6_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_6_1  (
            .in0(_gnd_net_),
            .in1(N__27660),
            .in2(N__27624),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_0 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_6_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_6_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_6_2  (
            .in0(_gnd_net_),
            .in1(N__27498),
            .in2(N__27543),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_1 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_6_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_6_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_6_3  (
            .in0(_gnd_net_),
            .in1(N__32070),
            .in2(N__27435),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_2 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_6_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_6_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_6_4  (
            .in0(_gnd_net_),
            .in1(N__32103),
            .in2(N__27362),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_3 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_6_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_6_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_6_5  (
            .in0(_gnd_net_),
            .in1(N__27290),
            .in2(N__32142),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_4 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_6_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_6_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_6_6  (
            .in0(_gnd_net_),
            .in1(N__29241),
            .in2(N__27222),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_5 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_6_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_6_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_6_7  (
            .in0(_gnd_net_),
            .in1(N__29214),
            .in2(N__27927),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_cry_6 ),
            .carryout(\this_ppu.un1_M_vaddress_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIF7IO_LC_20_7_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIF7IO_LC_20_7_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIF7IO_LC_20_7_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIF7IO_LC_20_7_0  (
            .in0(N__27903),
            .in1(N__24870),
            .in2(N__24864),
            .in3(N__24855),
            .lcout(\this_ppu.vscroll8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_20_7_6 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_20_7_6 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_20_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_20_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31815),
            .lcout(M_this_oam_ram_read_data_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_2_LC_20_9_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_2_LC_20_9_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_2_LC_20_9_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_2_LC_20_9_6 (
            .in0(N__35136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36853),
            .ce(N__30228),
            .sr(N__36024));
    defparam M_this_oam_address_q_0_LC_20_13_6.C_ON=1'b0;
    defparam M_this_oam_address_q_0_LC_20_13_6.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_0_LC_20_13_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 M_this_oam_address_q_0_LC_20_13_6 (
            .in0(N__30844),
            .in1(N__30648),
            .in2(_gnd_net_),
            .in3(N__33239),
            .lcout(M_this_oam_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36879),
            .ce(),
            .sr(N__32214));
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_20_14_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNINGCA_0_LC_20_14_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.M_vaddress_q_RNINGCA_0_LC_20_14_1  (
            .in0(_gnd_net_),
            .in1(N__27815),
            .in2(_gnd_net_),
            .in3(N__27869),
            .lcout(\this_ppu.un2_vscroll_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIO1A21_0_LC_20_15_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIO1A21_0_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIO1A21_0_LC_20_15_3 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \this_ppu.M_vaddress_q_RNIO1A21_0_LC_20_15_3  (
            .in0(N__24819),
            .in1(N__33748),
            .in2(N__33897),
            .in3(N__27816),
            .lcout(M_this_ppu_sprites_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI0A0E_6_LC_20_15_4.C_ON=1'b0;
    defparam M_this_state_q_RNI0A0E_6_LC_20_15_4.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI0A0E_6_LC_20_15_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 M_this_state_q_RNI0A0E_6_LC_20_15_4 (
            .in0(_gnd_net_),
            .in1(N__29334),
            .in2(_gnd_net_),
            .in3(N__27037),
            .lcout(M_this_state_q_RNI0A0EZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI244K2_6_LC_20_17_1.C_ON=1'b0;
    defparam M_this_state_q_RNI244K2_6_LC_20_17_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI244K2_6_LC_20_17_1.LUT_INIT=16'b0001010100111111;
    LogicCell40 M_this_state_q_RNI244K2_6_LC_20_17_1 (
            .in0(N__28143),
            .in1(N__24996),
            .in2(N__24879),
            .in3(N__29552),
            .lcout(),
            .ltout(M_this_state_q_RNI244K2Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIITVO4_7_LC_20_17_2.C_ON=1'b0;
    defparam M_this_state_q_RNIITVO4_7_LC_20_17_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIITVO4_7_LC_20_17_2.LUT_INIT=16'b0000110010001100;
    LogicCell40 M_this_state_q_RNIITVO4_7_LC_20_17_2 (
            .in0(N__25518),
            .in1(N__24885),
            .in2(N__24987),
            .in3(N__30376),
            .lcout(dma_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a4_5_LC_20_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a4_5_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a4_5_LC_20_17_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a4_5_LC_20_17_4  (
            .in0(N__35233),
            .in1(N__36334),
            .in2(_gnd_net_),
            .in3(N__29762),
            .lcout(N_661),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_82_i_0_o2_LC_20_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.N_82_i_0_o2_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_82_i_0_o2_LC_20_18_3 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.N_82_i_0_o2_LC_20_18_3  (
            .in0(N__27169),
            .in1(N__25163),
            .in2(N__25127),
            .in3(N__25055),
            .lcout(\this_vga_signals.N_428_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_a2_LC_20_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_a2_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_a2_LC_20_18_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_a2_LC_20_18_5  (
            .in0(N__29363),
            .in1(N__24909),
            .in2(_gnd_net_),
            .in3(N__30586),
            .lcout(N_861),
            .ltout(N_861_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIG5R81_10_LC_20_18_6.C_ON=1'b0;
    defparam M_this_state_q_RNIG5R81_10_LC_20_18_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIG5R81_10_LC_20_18_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 M_this_state_q_RNIG5R81_10_LC_20_18_6 (
            .in0(N__29418),
            .in1(N__28009),
            .in2(N__24888),
            .in3(N__27168),
            .lcout(dma_c4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un20_i_a2_4_a3_0_a4_2_1_LC_20_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un20_i_a2_4_a3_0_a4_2_1_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un20_i_a2_4_a3_0_a4_2_1_LC_20_18_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un20_i_a2_4_a3_0_a4_2_1_LC_20_18_7  (
            .in0(N__28008),
            .in1(N__30375),
            .in2(N__29374),
            .in3(N__27123),
            .lcout(this_vga_signals_un20_i_a2_4_a3_0_a4_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_13_LC_20_19_2.C_ON=1'b0;
    defparam M_this_state_q_13_LC_20_19_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_13_LC_20_19_2.LUT_INIT=16'b1111001000100010;
    LogicCell40 M_this_state_q_13_LC_20_19_2 (
            .in0(N__30597),
            .in1(N__31002),
            .in2(N__27197),
            .in3(N__29417),
            .lcout(M_this_state_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36924),
            .ce(),
            .sr(N__36009));
    defparam \this_vga_signals.M_this_state_q_ns_i_0_0_o2_13_LC_20_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_i_0_0_o2_13_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_i_0_0_o2_13_LC_20_19_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_i_0_0_o2_13_LC_20_19_3  (
            .in0(_gnd_net_),
            .in1(N__31539),
            .in2(_gnd_net_),
            .in3(N__30285),
            .lcout(N_460_0),
            .ltout(N_460_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_11_LC_20_19_4.C_ON=1'b0;
    defparam M_this_state_q_11_LC_20_19_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_20_19_4.LUT_INIT=16'b0011001000100010;
    LogicCell40 M_this_state_q_11_LC_20_19_4 (
            .in0(N__29373),
            .in1(N__31001),
            .in2(N__25365),
            .in3(N__28010),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36924),
            .ce(),
            .sr(N__36009));
    defparam M_this_state_q_10_LC_20_19_5.C_ON=1'b0;
    defparam M_this_state_q_10_LC_20_19_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_20_19_5.LUT_INIT=16'b1111111111111000;
    LogicCell40 M_this_state_q_10_LC_20_19_5 (
            .in0(N__28011),
            .in1(N__30488),
            .in2(N__25362),
            .in3(N__25205),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36924),
            .ce(),
            .sr(N__36009));
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_a2_0_LC_20_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_a2_0_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_a2_0_LC_20_20_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_qlde_i_0_a2_0_LC_20_20_0  (
            .in0(N__26775),
            .in1(N__29318),
            .in2(_gnd_net_),
            .in3(N__30966),
            .lcout(\this_vga_signals.N_745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_o2_1_LC_20_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_o2_1_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_o2_1_LC_20_20_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_o2_1_LC_20_20_1  (
            .in0(N__25126),
            .in1(N__25153),
            .in2(_gnd_net_),
            .in3(N__25044),
            .lcout(N_888_0),
            .ltout(N_888_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a2_5_LC_20_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a2_5_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a2_5_LC_20_20_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_oam_address_q_0_i_o3_0_a2_5_LC_20_20_2  (
            .in0(N__26776),
            .in1(N__35218),
            .in2(N__25176),
            .in3(N__29319),
            .lcout(M_this_oam_address_q_0_i_o3_0_a2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_0_0_LC_20_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_0_0_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_0_0_LC_20_20_4 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_i_a2_0_0_LC_20_20_4  (
            .in0(N__36313),
            .in1(_gnd_net_),
            .in2(N__26783),
            .in3(N__35219),
            .lcout(\this_vga_signals.N_779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_0_o4_LC_20_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_0_o4_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_0_o4_LC_20_20_5 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_0_o4_LC_20_20_5  (
            .in0(N__30593),
            .in1(N__25154),
            .in2(N__25128),
            .in3(N__25045),
            .lcout(N_413_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2_LC_20_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2_LC_20_20_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2_LC_20_20_6  (
            .in0(_gnd_net_),
            .in1(N__28193),
            .in2(_gnd_net_),
            .in3(N__29317),
            .lcout(un1_M_this_substate_q4_2_i_0_265_i_a2_0_a3_0_a2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_20_20_7.C_ON=1'b0;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_20_20_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_20_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_20_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36092),
            .lcout(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5L8_LC_20_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5L8_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5L8_LC_20_21_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5L8_LC_20_21_1  (
            .in0(N__25658),
            .in1(N__25595),
            .in2(N__25726),
            .in3(N__25817),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_5LZ0Z8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_LC_20_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_LC_20_21_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_1_LC_20_21_2  (
            .in0(N__35337),
            .in1(N__25569),
            .in2(N__25536),
            .in3(N__35346),
            .lcout(M_this_substate_d_0_sqmuxa),
            .ltout(M_this_substate_d_0_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_20_21_3.C_ON=1'b0;
    defparam M_this_state_q_1_LC_20_21_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_20_21_3.LUT_INIT=16'b1111000011111010;
    LogicCell40 M_this_state_q_1_LC_20_21_3 (
            .in0(N__26316),
            .in1(_gnd_net_),
            .in2(N__25521),
            .in3(N__31003),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36932),
            .ce(),
            .sr(N__36012));
    defparam M_this_state_q_RNITB0L_3_LC_20_21_6.C_ON=1'b0;
    defparam M_this_state_q_RNITB0L_3_LC_20_21_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNITB0L_3_LC_20_21_6.LUT_INIT=16'b0000000000010001;
    LogicCell40 M_this_state_q_RNITB0L_3_LC_20_21_6 (
            .in0(N__28202),
            .in1(N__27124),
            .in2(_gnd_net_),
            .in3(N__26315),
            .lcout(dma_c4_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_2_LC_20_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_2_LC_20_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_2_LC_20_21_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0_2_LC_20_21_7  (
            .in0(N__25707),
            .in1(N__25816),
            .in2(_gnd_net_),
            .in3(N__31566),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_12_LC_20_22_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_12_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_12_LC_20_22_0 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_12_LC_20_22_0  (
            .in0(N__26314),
            .in1(N__25506),
            .in2(N__25374),
            .in3(N__25391),
            .lcout(),
            .ltout(N_622_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_12_LC_20_22_1.C_ON=1'b0;
    defparam M_this_sprites_address_q_12_LC_20_22_1.SEQ_MODE=4'b1000;
    defparam M_this_sprites_address_q_12_LC_20_22_1.LUT_INIT=16'b0000111000000000;
    LogicCell40 M_this_sprites_address_q_12_LC_20_22_1 (
            .in0(N__25392),
            .in1(N__25380),
            .in2(N__25383),
            .in3(N__26562),
            .lcout(M_this_sprites_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36936),
            .ce(),
            .sr(N__32212));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_448_tz_LC_20_22_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_448_tz_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_448_tz_LC_20_22_2 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_448_tz_LC_20_22_2  (
            .in0(N__26313),
            .in1(N__31101),
            .in2(N__26552),
            .in3(N__34955),
            .lcout(N_1278_tz_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_12_LC_20_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_12_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_12_LC_20_22_3 .LUT_INIT=16'b0001000100110001;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0_12_LC_20_22_3  (
            .in0(N__34954),
            .in1(N__36314),
            .in2(N__31142),
            .in3(N__26941),
            .lcout(\this_vga_signals.M_this_sprites_address_q_0_0_i_a4_0_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_12_LC_20_22_4.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_12_LC_20_22_4.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_12_LC_20_22_4.LUT_INIT=16'b1010111100000011;
    LogicCell40 M_this_sprites_address_q_RNO_0_12_LC_20_22_4 (
            .in0(N__26942),
            .in1(N__26123),
            .in2(N__26220),
            .in3(N__34956),
            .lcout(M_this_sprites_address_qc_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_o2_2_0_LC_20_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_o2_2_0_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_o2_2_0_LC_20_22_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_i_o2_2_0_LC_20_22_5  (
            .in0(_gnd_net_),
            .in1(N__26939),
            .in2(_gnd_net_),
            .in3(N__26311),
            .lcout(\this_vga_signals.N_427_0 ),
            .ltout(\this_vga_signals.N_427_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_444_tz_LC_20_22_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_444_tz_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_444_tz_LC_20_22_6 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_444_tz_LC_20_22_6  (
            .in0(N__26312),
            .in1(N__34831),
            .in2(N__26271),
            .in3(N__31097),
            .lcout(N_1274_tz_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_13_LC_20_22_7.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_13_LC_20_22_7.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_13_LC_20_22_7.LUT_INIT=16'b1101110100000101;
    LogicCell40 M_this_sprites_address_q_RNO_0_13_LC_20_22_7 (
            .in0(N__26173),
            .in1(N__26940),
            .in2(N__26129),
            .in3(N__34818),
            .lcout(M_this_sprites_address_qc_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_o2_LC_20_23_0 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_o2_LC_20_23_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_o2_LC_20_23_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_6_0_0_o2_LC_20_23_0  (
            .in0(_gnd_net_),
            .in1(N__27154),
            .in2(_gnd_net_),
            .in3(N__27110),
            .lcout(\this_vga_signals.N_889_0 ),
            .ltout(\this_vga_signals.N_889_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_LC_20_23_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_LC_20_23_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_LC_20_23_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vga_signals.M_this_sprites_address_q_0_0_i_a2_0_LC_20_23_1  (
            .in0(N__36323),
            .in1(N__31702),
            .in2(N__26223),
            .in3(N__30431),
            .lcout(N_750),
            .ltout(N_750_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_sprites_address_q_RNO_0_9_LC_20_23_2.C_ON=1'b0;
    defparam M_this_sprites_address_q_RNO_0_9_LC_20_23_2.SEQ_MODE=4'b0000;
    defparam M_this_sprites_address_q_RNO_0_9_LC_20_23_2.LUT_INIT=16'b1100110100001101;
    LogicCell40 M_this_sprites_address_q_RNO_0_9_LC_20_23_2 (
            .in0(N__26124),
            .in1(N__25952),
            .in2(N__25842),
            .in3(N__26985),
            .lcout(M_this_sprites_address_qc_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_20_23_4.C_ON=1'b0;
    defparam M_this_state_q_3_LC_20_23_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_20_23_4.LUT_INIT=16'b1101110011001100;
    LogicCell40 M_this_state_q_3_LC_20_23_4 (
            .in0(N__25818),
            .in1(N__25755),
            .in2(N__25742),
            .in3(N__27080),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36943),
            .ce(),
            .sr(N__36019));
    defparam M_this_state_q_8_LC_20_23_5.C_ON=1'b0;
    defparam M_this_state_q_8_LC_20_23_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_20_23_5.LUT_INIT=16'b0101010101000000;
    LogicCell40 M_this_state_q_8_LC_20_23_5 (
            .in0(N__31084),
            .in1(N__30377),
            .in2(N__27204),
            .in3(N__27161),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36943),
            .ce(),
            .sr(N__36019));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_o2_0_LC_20_23_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_o2_0_LC_20_23_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_o2_0_LC_20_23_6 .LUT_INIT=16'b1010101100001111;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_i_i_o2_0_LC_20_23_6  (
            .in0(N__27160),
            .in1(N__27111),
            .in2(N__30442),
            .in3(N__31082),
            .lcout(\this_vga_signals.N_431_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_20_23_7.C_ON=1'b0;
    defparam M_this_state_q_2_LC_20_23_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_20_23_7.LUT_INIT=16'b1101110001010000;
    LogicCell40 M_this_state_q_2_LC_20_23_7 (
            .in0(N__31083),
            .in1(N__27090),
            .in2(N__27036),
            .in3(N__27081),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36943),
            .ce(),
            .sr(N__36019));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_3_LC_20_24_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_3_LC_20_24_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_3_LC_20_24_1 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_3_LC_20_24_1  (
            .in0(N__28523),
            .in1(N__35826),
            .in2(N__34577),
            .in3(N__28547),
            .lcout(N_250),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3_0_LC_20_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3_0_LC_20_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3_0_LC_20_24_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3_0_LC_20_24_2  (
            .in0(N__32383),
            .in1(N__34573),
            .in2(N__35846),
            .in3(N__31324),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_0_LC_20_24_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_0_LC_20_24_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_0_LC_20_24_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_i_a2_1_0_LC_20_24_3  (
            .in0(_gnd_net_),
            .in1(N__34444),
            .in2(N__26790),
            .in3(N__33355),
            .lcout(\this_vga_signals.N_743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_1_LC_20_24_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_1_LC_20_24_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_1_LC_20_24_4 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_1_LC_20_24_4  (
            .in0(N__33354),
            .in1(N__28545),
            .in2(N__36348),
            .in3(N__28521),
            .lcout(N_228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_2_LC_20_24_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_2_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_2_LC_20_24_5 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_2_LC_20_24_5  (
            .in0(N__28522),
            .in1(N__34443),
            .in2(N__35207),
            .in3(N__28546),
            .lcout(N_248),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_6_LC_21_5_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_6_LC_21_5_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_6_LC_21_5_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_6_LC_21_5_0 (
            .in0(N__34441),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36848),
            .ce(N__30230),
            .sr(N__36029));
    defparam M_this_data_tmp_q_esr_1_LC_21_5_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_1_LC_21_5_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_1_LC_21_5_5.LUT_INIT=16'b1100110011001100;
    LogicCell40 M_this_data_tmp_q_esr_1_LC_21_5_5 (
            .in0(_gnd_net_),
            .in1(N__33411),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36848),
            .ce(N__30230),
            .sr(N__36029));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_21_6_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_21_6_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_21_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_21_6_0  (
            .in0(_gnd_net_),
            .in1(N__27864),
            .in2(N__27737),
            .in3(N__27825),
            .lcout(\this_ppu.M_this_ppu_vram_addr_i_7 ),
            .ltout(),
            .carryin(bfn_21_6_0_),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_21_6_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_21_6_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_21_6_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_21_6_1  (
            .in0(N__27716),
            .in1(N__27655),
            .in2(N__27623),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_vaddress_q_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_0 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_21_6_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_21_6_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_21_6_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_21_6_2  (
            .in0(N__27603),
            .in1(N__27497),
            .in2(N__27538),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_vaddress_q_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_1 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_21_6_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_21_6_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_21_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_21_6_3  (
            .in0(_gnd_net_),
            .in1(N__27882),
            .in2(N__27434),
            .in3(N__27476),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_5 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_2 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_21_6_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_21_6_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_21_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_21_6_4  (
            .in0(_gnd_net_),
            .in1(N__29142),
            .in2(N__27363),
            .in3(N__27404),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_6 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_3 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_21_6_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_21_6_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_21_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_21_6_5  (
            .in0(_gnd_net_),
            .in1(N__32031),
            .in2(N__27291),
            .in3(N__27335),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_7 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_4 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_21_6_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_21_6_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_21_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_21_6_6  (
            .in0(_gnd_net_),
            .in1(N__29265),
            .in2(N__27221),
            .in3(N__27272),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_8 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_5 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_21_6_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_21_6_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_21_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_21_6_7  (
            .in0(_gnd_net_),
            .in1(N__29178),
            .in2(N__27923),
            .in3(N__27968),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_9 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_vaddress_q_3_cry_6 ),
            .carryout(\this_ppu.un1_M_vaddress_q_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_21_7_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_21_7_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_21_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_21_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27906),
            .lcout(\this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_16_LC_21_7_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_16_LC_21_7_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_16_LC_21_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a4_16_LC_21_7_2  (
            .in0(_gnd_net_),
            .in1(N__27876),
            .in2(_gnd_net_),
            .in3(N__35707),
            .lcout(M_this_oam_ram_write_data_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_7_4 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_7_4 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32066),
            .lcout(M_this_oam_ram_read_data_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_16_LC_21_8_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_16_LC_21_8_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_16_LC_21_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_16_LC_21_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31350),
            .lcout(M_this_data_tmp_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36854),
            .ce(N__34019),
            .sr(N__36025));
    defparam M_this_data_tmp_q_esr_17_LC_21_8_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_17_LC_21_8_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_17_LC_21_8_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_17_LC_21_8_1 (
            .in0(N__33407),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36854),
            .ce(N__34019),
            .sr(N__36025));
    defparam M_this_data_tmp_q_esr_23_LC_21_8_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_23_LC_21_8_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_23_LC_21_8_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_23_LC_21_8_3 (
            .in0(N__34542),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36854),
            .ce(N__34019),
            .sr(N__36025));
    defparam M_this_data_tmp_q_esr_3_LC_21_10_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_3_LC_21_10_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_3_LC_21_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_3_LC_21_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35868),
            .lcout(M_this_data_tmp_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36866),
            .ce(N__30215),
            .sr(N__36020));
    defparam M_this_data_tmp_q_esr_7_LC_21_10_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_7_LC_21_10_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_7_LC_21_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_7_LC_21_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34514),
            .lcout(M_this_data_tmp_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36866),
            .ce(N__30215),
            .sr(N__36020));
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_21_11_0.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_21_11_0.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_21_11_0.LUT_INIT=16'b1111111100010000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_1_LC_21_11_0 (
            .in0(N__30558),
            .in1(N__30658),
            .in2(N__30853),
            .in3(N__36102),
            .lcout(N_1412_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un20_i_a2_0_a3_0_a4_2_2_LC_21_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un20_i_a2_0_a3_0_a4_2_2_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un20_i_a2_0_a3_0_a4_2_2_LC_21_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un20_i_a2_0_a3_0_a4_2_2_LC_21_17_7  (
            .in0(N__31205),
            .in1(N__29402),
            .in2(N__30605),
            .in3(N__30378),
            .lcout(this_vga_signals_un20_i_a2_0_a3_0_a4_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_a2_LC_21_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_a2_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_6_0_0_a2_LC_21_18_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_6_0_0_a2_LC_21_18_2  (
            .in0(N__35220),
            .in1(N__36333),
            .in2(_gnd_net_),
            .in3(N__29763),
            .lcout(\this_vga_signals.N_747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_en_iv_i_0_0_LC_21_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_iv_i_0_0_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_en_iv_i_0_0_LC_21_18_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_en_iv_i_0_0_LC_21_18_4  (
            .in0(_gnd_net_),
            .in1(N__28510),
            .in2(_gnd_net_),
            .in3(N__30438),
            .lcout(N_25_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_18_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_18_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_18_7  (
            .in0(N__28137),
            .in1(N__28122),
            .in2(_gnd_net_),
            .in3(N__28110),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_LC_21_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_LC_21_19_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_o2_LC_21_19_4  (
            .in0(N__29416),
            .in1(N__28007),
            .in2(_gnd_net_),
            .in3(N__30361),
            .lcout(\this_vga_signals.N_433_0 ),
            .ltout(\this_vga_signals.N_433_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_0_LC_21_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_0_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_0_LC_21_19_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_o2_0_LC_21_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27987),
            .in3(N__30279),
            .lcout(\this_vga_signals.N_442_0 ),
            .ltout(\this_vga_signals.N_442_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_a4_0_LC_21_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_a4_0_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_a4_0_LC_21_19_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_a4_0_LC_21_19_6  (
            .in0(N__29329),
            .in1(N__28203),
            .in2(N__27984),
            .in3(N__31000),
            .lcout(),
            .ltout(\this_vga_signals.N_719_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_1_LC_21_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_1_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_1_LC_21_19_7 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_1_LC_21_19_7  (
            .in0(N__29548),
            .in1(N__30323),
            .in2(N__27981),
            .in3(N__30480),
            .lcout(\this_vga_signals.M_this_data_count_qlde_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_21_20_0.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_21_20_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_21_20_0.LUT_INIT=16'b1000100011110000;
    LogicCell40 M_this_data_count_q_2_LC_21_20_0 (
            .in0(N__28215),
            .in1(N__31670),
            .in2(N__28233),
            .in3(N__31486),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36933),
            .ce(N__31392),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_a3_0_a4_0_2_LC_21_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_a3_0_a4_0_2_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_a3_0_a4_0_2_LC_21_20_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_a3_0_a4_0_2_LC_21_20_1  (
            .in0(N__28195),
            .in1(_gnd_net_),
            .in2(N__36332),
            .in3(N__36090),
            .lcout(this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2),
            .ltout(this_vga_signals_M_this_data_count_q_3_0_a3_0_a4_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_i_i_10_LC_21_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_i_i_10_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_i_i_10_LC_21_20_2 .LUT_INIT=16'b0001001111011111;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_i_i_10_LC_21_20_2  (
            .in0(N__29751),
            .in1(N__35211),
            .in2(N__28209),
            .in3(N__28260),
            .lcout(),
            .ltout(N_307_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_21_20_3.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_21_20_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_21_20_3.LUT_INIT=16'b0100111000011011;
    LogicCell40 M_this_data_count_q_10_LC_21_20_3 (
            .in0(N__31487),
            .in1(N__28302),
            .in2(N__28206),
            .in3(N__29518),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36933),
            .ce(N__31392),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_i_i_a2_10_LC_21_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_i_i_a2_10_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_i_i_a2_10_LC_21_20_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_i_i_a2_10_LC_21_20_4  (
            .in0(N__36089),
            .in1(N__28194),
            .in2(_gnd_net_),
            .in3(N__31076),
            .lcout(N_755),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_a4_0_1_13_LC_21_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_a4_0_1_13_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_a4_0_1_13_LC_21_20_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_0_a4_0_1_13_LC_21_20_5  (
            .in0(N__36303),
            .in1(N__29750),
            .in2(N__35228),
            .in3(N__36088),
            .lcout(\this_vga_signals.N_665_1 ),
            .ltout(\this_vga_signals.N_665_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_13_LC_21_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_13_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_q_3_0_0_13_LC_21_20_6 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \this_vga_signals.M_this_data_count_q_3_0_0_13_LC_21_20_6  (
            .in0(_gnd_net_),
            .in1(N__36302),
            .in2(N__28149),
            .in3(N__28259),
            .lcout(),
            .ltout(M_this_data_count_q_3_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_21_20_7.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_21_20_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_21_20_7.LUT_INIT=16'b0100111000011011;
    LogicCell40 M_this_data_count_q_13_LC_21_20_7 (
            .in0(N__31488),
            .in1(N__29136),
            .in2(N__28146),
            .in3(N__29819),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36933),
            .ce(N__31392),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_21_21_0.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_21_21_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_21_21_0.LUT_INIT=16'b1110001000100010;
    LogicCell40 M_this_data_count_q_11_LC_21_21_0 (
            .in0(N__28290),
            .in1(N__31479),
            .in2(N__35847),
            .in3(N__28263),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36937),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_21_21_2.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_21_21_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_21_21_2.LUT_INIT=16'b1110001000100010;
    LogicCell40 M_this_data_count_q_12_LC_21_21_2 (
            .in0(N__28278),
            .in1(N__31480),
            .in2(N__32413),
            .in3(N__28264),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36937),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_14_LC_21_21_3.C_ON=1'b0;
    defparam M_this_data_count_q_14_LC_21_21_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_14_LC_21_21_3.LUT_INIT=16'b1010000011001100;
    LogicCell40 M_this_data_count_q_14_LC_21_21_3 (
            .in0(N__28261),
            .in1(N__28578),
            .in2(N__34442),
            .in3(N__31483),
            .lcout(M_this_data_count_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36937),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_15_LC_21_21_4.C_ON=1'b0;
    defparam M_this_data_count_q_15_LC_21_21_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_15_LC_21_21_4.LUT_INIT=16'b1110001000100010;
    LogicCell40 M_this_data_count_q_15_LC_21_21_4 (
            .in0(N__28563),
            .in1(N__31481),
            .in2(N__34569),
            .in3(N__28265),
            .lcout(M_this_data_count_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36937),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_21_21_5.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_21_21_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_21_21_5.LUT_INIT=16'b1010000011001100;
    LogicCell40 M_this_data_count_q_8_LC_21_21_5 (
            .in0(N__28262),
            .in1(N__28329),
            .in2(N__31362),
            .in3(N__31484),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36937),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_21_21_6.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_21_21_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_21_21_6.LUT_INIT=16'b1110001000100010;
    LogicCell40 M_this_data_count_q_9_LC_21_21_6 (
            .in0(N__28317),
            .in1(N__31482),
            .in2(N__33391),
            .in3(N__28266),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36937),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_21_21_7.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_21_21_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_21_21_7.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_0_LC_21_21_7 (
            .in0(_gnd_net_),
            .in1(N__31485),
            .in2(_gnd_net_),
            .in3(N__29586),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36937),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_c_0_LC_21_22_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_21_22_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_21_22_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_21_22_0 (
            .in0(_gnd_net_),
            .in1(N__29585),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_22_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_21_22_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_21_22_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_21_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_0_THRU_LUT4_0_LC_21_22_1 (
            .in0(_gnd_net_),
            .in1(N__28980),
            .in2(N__30030),
            .in3(N__28236),
            .lcout(M_this_data_count_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_2_LC_21_22_2.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_2_LC_21_22_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_2_LC_21_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_2_LC_21_22_2 (
            .in0(_gnd_net_),
            .in1(N__29601),
            .in2(N__29046),
            .in3(N__28221),
            .lcout(M_this_data_count_q_s_2),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_21_22_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_21_22_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_21_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_2_THRU_LUT4_0_LC_21_22_3 (
            .in0(_gnd_net_),
            .in1(N__28981),
            .in2(N__30000),
            .in3(N__28218),
            .lcout(M_this_data_count_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_21_22_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_21_22_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_21_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_3_THRU_LUT4_0_LC_21_22_4 (
            .in0(_gnd_net_),
            .in1(N__29969),
            .in2(N__29047),
            .in3(N__28341),
            .lcout(M_this_data_count_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_21_22_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_21_22_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_21_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_4_THRU_LUT4_0_LC_21_22_5 (
            .in0(_gnd_net_),
            .in1(N__28985),
            .in2(N__29946),
            .in3(N__28338),
            .lcout(M_this_data_count_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_21_22_6.C_ON=1'b1;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_21_22_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_21_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_5_THRU_LUT4_0_LC_21_22_6 (
            .in0(_gnd_net_),
            .in1(N__29917),
            .in2(N__29048),
            .in3(N__28335),
            .lcout(M_this_data_count_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_21_22_7.C_ON=1'b1;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_21_22_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_21_22_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_6_THRU_LUT4_0_LC_21_22_7 (
            .in0(_gnd_net_),
            .in1(N__28989),
            .in2(N__31431),
            .in3(N__28332),
            .lcout(M_this_data_count_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_8_LC_21_23_0.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_8_LC_21_23_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_8_LC_21_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_8_LC_21_23_0 (
            .in0(_gnd_net_),
            .in1(N__29003),
            .in2(N__29460),
            .in3(N__28320),
            .lcout(M_this_data_count_q_s_8),
            .ltout(),
            .carryin(bfn_21_23_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_9_LC_21_23_1.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_9_LC_21_23_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_9_LC_21_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_9_LC_21_23_1 (
            .in0(_gnd_net_),
            .in1(N__29496),
            .in2(N__29063),
            .in3(N__28305),
            .lcout(M_this_data_count_q_s_9),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_21_23_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_21_23_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_9_THRU_LUT4_0_LC_21_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_9_THRU_LUT4_0_LC_21_23_2 (
            .in0(_gnd_net_),
            .in1(N__29010),
            .in2(N__29526),
            .in3(N__28293),
            .lcout(M_this_data_count_q_cry_9_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_11_LC_21_23_3.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_11_LC_21_23_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_11_LC_21_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_11_LC_21_23_3 (
            .in0(_gnd_net_),
            .in1(N__29480),
            .in2(N__29062),
            .in3(N__28281),
            .lcout(M_this_data_count_q_s_11),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_12_LC_21_23_4.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_12_LC_21_23_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_12_LC_21_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_12_LC_21_23_4 (
            .in0(_gnd_net_),
            .in1(N__29001),
            .in2(N__29781),
            .in3(N__28269),
            .lcout(M_this_data_count_q_s_12),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_21_23_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_21_23_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_12_THRU_LUT4_0_LC_21_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_12_THRU_LUT4_0_LC_21_23_5 (
            .in0(_gnd_net_),
            .in1(N__29820),
            .in2(N__29064),
            .in3(N__29127),
            .lcout(M_this_data_count_q_cry_12_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_12),
            .carryout(M_this_data_count_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_14_LC_21_23_6.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_14_LC_21_23_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_14_LC_21_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_14_LC_21_23_6 (
            .in0(_gnd_net_),
            .in1(N__29002),
            .in2(N__29838),
            .in3(N__28569),
            .lcout(M_this_data_count_q_s_14),
            .ltout(),
            .carryin(M_this_data_count_q_cry_13),
            .carryout(M_this_data_count_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_15_LC_21_23_7.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_15_LC_21_23_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_15_LC_21_23_7.LUT_INIT=16'b1100110000110011;
    LogicCell40 M_this_data_count_q_RNO_0_15_LC_21_23_7 (
            .in0(_gnd_net_),
            .in1(N__29799),
            .in2(_gnd_net_),
            .in3(N__28566),
            .lcout(M_this_data_count_q_s_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_0_LC_21_25_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_0_LC_21_25_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_0_LC_21_25_2 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_i_i_i_0_LC_21_25_2  (
            .in0(N__31356),
            .in1(N__28551),
            .in2(N__32405),
            .in3(N__28527),
            .lcout(N_226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_6_LC_22_5_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_6_LC_22_5_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_6_LC_22_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_6_LC_22_5_0  (
            .in0(_gnd_net_),
            .in1(N__28401),
            .in2(_gnd_net_),
            .in3(N__35690),
            .lcout(M_this_oam_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_2_LC_22_5_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_2_LC_22_5_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_2_LC_22_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_2_LC_22_5_4  (
            .in0(_gnd_net_),
            .in1(N__28383),
            .in2(_gnd_net_),
            .in3(N__35689),
            .lcout(M_this_oam_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_1_LC_22_5_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_1_LC_22_5_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_1_LC_22_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_1_LC_22_5_6  (
            .in0(_gnd_net_),
            .in1(N__28359),
            .in2(_gnd_net_),
            .in3(N__35688),
            .lcout(M_this_oam_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_4_LC_22_6_2.C_ON=1'b0;
    defparam M_this_oam_address_q_4_LC_22_6_2.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_4_LC_22_6_2.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_4_LC_22_6_2 (
            .in0(N__30066),
            .in1(N__33257),
            .in2(_gnd_net_),
            .in3(N__30770),
            .lcout(M_this_oam_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36850),
            .ce(),
            .sr(N__32217));
    defparam M_this_oam_address_q_5_LC_22_6_3.C_ON=1'b0;
    defparam M_this_oam_address_q_5_LC_22_6_3.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_5_LC_22_6_3.LUT_INIT=16'b0000011000001100;
    LogicCell40 M_this_oam_address_q_5_LC_22_6_3 (
            .in0(N__30771),
            .in1(N__30106),
            .in2(N__33261),
            .in3(N__30067),
            .lcout(M_this_oam_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36850),
            .ce(),
            .sr(N__32217));
    defparam \this_ppu.un1_oam_data_ac0_1_LC_22_7_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_ac0_1_LC_22_7_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_ac0_1_LC_22_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.un1_oam_data_ac0_1_LC_22_7_1  (
            .in0(_gnd_net_),
            .in1(N__32098),
            .in2(_gnd_net_),
            .in3(N__32064),
            .lcout(\this_ppu.un1_oam_data_c2 ),
            .ltout(\this_ppu.un1_oam_data_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc3_LC_22_7_2 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc3_LC_22_7_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc3_LC_22_7_2 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \this_ppu.un1_oam_data_axbxc3_LC_22_7_2  (
            .in0(N__29239),
            .in1(_gnd_net_),
            .in2(N__29268),
            .in3(N__32137),
            .lcout(\this_ppu.un1_M_vaddress_q_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_23_LC_22_7_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_23_LC_22_7_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_23_LC_22_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_23_LC_22_7_3  (
            .in0(_gnd_net_),
            .in1(N__29259),
            .in2(_gnd_net_),
            .in3(N__35627),
            .lcout(M_this_oam_ram_write_data_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc4_LC_22_7_4 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc4_LC_22_7_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc4_LC_22_7_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.un1_oam_data_axbxc4_LC_22_7_4  (
            .in0(N__29240),
            .in1(N__32138),
            .in2(N__29213),
            .in3(N__29184),
            .lcout(\this_ppu.un1_M_vaddress_q_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_25_LC_22_7_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_25_LC_22_7_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_25_LC_22_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_25_LC_22_7_5  (
            .in0(_gnd_net_),
            .in1(N__33359),
            .in2(_gnd_net_),
            .in3(N__35626),
            .lcout(M_this_oam_ram_write_data_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_17_LC_22_7_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_17_LC_22_7_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_17_LC_22_7_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a4_17_LC_22_7_6  (
            .in0(N__35628),
            .in1(_gnd_net_),
            .in2(N__29163),
            .in3(_gnd_net_),
            .lcout(M_this_oam_ram_write_data_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc1_LC_22_7_7 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc1_LC_22_7_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc1_LC_22_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_oam_data_axbxc1_LC_22_7_7  (
            .in0(_gnd_net_),
            .in1(N__32099),
            .in2(_gnd_net_),
            .in3(N__32065),
            .lcout(\this_ppu.un1_M_vaddress_q_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_22_LC_22_8_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_22_LC_22_8_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_22_LC_22_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_22_LC_22_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34440),
            .lcout(M_this_data_tmp_qZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36858),
            .ce(N__34018),
            .sr(N__36022));
    defparam M_this_data_tmp_q_esr_21_LC_22_8_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_21_LC_22_8_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_21_LC_22_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_21_LC_22_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36252),
            .lcout(M_this_data_tmp_qZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36858),
            .ce(N__34018),
            .sr(N__36022));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_24_LC_22_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_24_LC_22_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_24_LC_22_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_24_LC_22_9_7  (
            .in0(_gnd_net_),
            .in1(N__31351),
            .in2(_gnd_net_),
            .in3(N__35625),
            .lcout(M_this_oam_ram_write_data_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_22_11_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_22_11_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_22_11_4.LUT_INIT=16'b1111111101000000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_0_1_LC_22_11_4 (
            .in0(N__30556),
            .in1(N__30669),
            .in2(N__30845),
            .in3(N__36101),
            .lcout(N_1404_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_1_LC_22_14_1.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_22_14_1.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_22_14_1.LUT_INIT=16'b1111111100100000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_LC_22_14_1 (
            .in0(N__30552),
            .in1(N__30668),
            .in2(N__30852),
            .in3(N__36100),
            .lcout(N_1396_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_1_LC_22_16_1.C_ON=1'b0;
    defparam M_this_oam_address_q_1_LC_22_16_1.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_1_LC_22_16_1.LUT_INIT=16'b0000000001101010;
    LogicCell40 M_this_oam_address_q_1_LC_22_16_1 (
            .in0(N__30547),
            .in1(N__30666),
            .in2(N__30855),
            .in3(N__33250),
            .lcout(M_this_oam_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36915),
            .ce(),
            .sr(N__32213));
    defparam M_this_state_q_12_LC_22_17_7.C_ON=1'b0;
    defparam M_this_state_q_12_LC_22_17_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_22_17_7.LUT_INIT=16'b1111111011111010;
    LogicCell40 M_this_state_q_12_LC_22_17_7 (
            .in0(N__33227),
            .in1(N__29406),
            .in2(N__30854),
            .in3(N__30489),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36925),
            .ce(),
            .sr(N__36005));
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_o2_LC_22_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_o2_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_o2_LC_22_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.un1_M_this_substate_q4_1_i_0_251_i_0_o2_LC_22_19_1  (
            .in0(_gnd_net_),
            .in1(N__30604),
            .in2(_gnd_net_),
            .in3(N__29375),
            .lcout(),
            .ltout(\this_vga_signals.N_469_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_m2_LC_22_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_m2_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_m2_LC_22_19_2 .LUT_INIT=16'b0001000010111111;
    LogicCell40 \this_vga_signals.M_this_external_address_qlde_i_0_m2_LC_22_19_2  (
            .in0(N__31214),
            .in1(N__30444),
            .in2(N__29340),
            .in3(N__31118),
            .lcout(),
            .ltout(\this_vga_signals.N_506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_i_LC_22_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_i_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_i_LC_22_19_3 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \this_vga_signals.M_this_external_address_qlde_i_0_i_LC_22_19_3  (
            .in0(N__29727),
            .in1(N__36099),
            .in2(N__29337),
            .in3(N__29330),
            .lcout(N_47),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_1_LC_22_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_1_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_o2_1_LC_22_19_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_o2_1_LC_22_19_4  (
            .in0(N__30280),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31538),
            .lcout(\this_vga_signals.N_461_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNI60TF_15_LC_22_20_3.C_ON=1'b0;
    defparam M_this_data_count_q_RNI60TF_15_LC_22_20_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNI60TF_15_LC_22_20_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNI60TF_15_LC_22_20_3 (
            .in0(N__29831),
            .in1(N__29815),
            .in2(N__29798),
            .in3(N__29774),
            .lcout(M_this_state_d62_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_a2_LC_22_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_a2_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_qlde_i_0_a2_LC_22_20_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \this_vga_signals.M_this_external_address_qlde_i_0_a2_LC_22_20_4  (
            .in0(N__35164),
            .in1(N__36324),
            .in2(_gnd_net_),
            .in3(N__29761),
            .lcout(\this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2 ),
            .ltout(\this_vga_signals.M_this_external_address_qlde_i_0_aZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_data_count_qlde_i_i_LC_22_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_data_count_qlde_i_i_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_data_count_qlde_i_i_LC_22_20_5 .LUT_INIT=16'b1101110011111111;
    LogicCell40 \this_vga_signals.M_this_data_count_qlde_i_i_LC_22_20_5  (
            .in0(N__29721),
            .in1(N__29710),
            .in2(N__29610),
            .in3(N__29607),
            .lcout(N_364),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIQ9QL_0_LC_22_21_0.C_ON=1'b0;
    defparam M_this_data_count_q_RNIQ9QL_0_LC_22_21_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIQ9QL_0_LC_22_21_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIQ9QL_0_LC_22_21_0 (
            .in0(N__29597),
            .in1(N__30025),
            .in2(N__29999),
            .in3(N__29584),
            .lcout(),
            .ltout(M_this_state_d62_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNII1EE2_10_LC_22_21_1.C_ON=1'b0;
    defparam M_this_data_count_q_RNII1EE2_10_LC_22_21_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNII1EE2_10_LC_22_21_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_data_count_q_RNII1EE2_10_LC_22_21_1 (
            .in0(N__29568),
            .in1(N__29442),
            .in2(N__29559),
            .in3(N__29436),
            .lcout(M_this_state_d62),
            .ltout(M_this_state_d62_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_716_i_LC_22_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.N_716_i_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_716_i_LC_22_21_2 .LUT_INIT=16'b1111111111110011;
    LogicCell40 \this_vga_signals.N_716_i_LC_22_21_2  (
            .in0(_gnd_net_),
            .in1(N__29556),
            .in2(N__29529),
            .in3(N__36096),
            .lcout(N_716_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNI8TRI_10_LC_22_21_3.C_ON=1'b0;
    defparam M_this_data_count_q_RNI8TRI_10_LC_22_21_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNI8TRI_10_LC_22_21_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNI8TRI_10_LC_22_21_3 (
            .in0(N__29519),
            .in1(N__29492),
            .in2(N__29481),
            .in3(N__29453),
            .lcout(M_this_state_d62_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIAQQL_4_LC_22_21_4.C_ON=1'b0;
    defparam M_this_data_count_q_RNIAQQL_4_LC_22_21_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIAQQL_4_LC_22_21_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIAQQL_4_LC_22_21_4 (
            .in0(N__29919),
            .in1(N__29941),
            .in2(N__31427),
            .in3(N__29968),
            .lcout(M_this_state_d62_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_22_22_0.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_22_22_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_22_22_0.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_1_LC_22_22_0 (
            .in0(N__30036),
            .in1(N__31489),
            .in2(_gnd_net_),
            .in3(N__30029),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36947),
            .ce(N__31393),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_22_22_1.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_22_22_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_22_22_1.LUT_INIT=16'b0101000000000101;
    LogicCell40 M_this_data_count_q_3_LC_22_22_1 (
            .in0(N__31490),
            .in1(_gnd_net_),
            .in2(N__30009),
            .in3(N__29998),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36947),
            .ce(N__31393),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_22_22_2.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_22_22_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_22_22_2.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_4_LC_22_22_2 (
            .in0(N__29976),
            .in1(N__31491),
            .in2(_gnd_net_),
            .in3(N__29970),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36947),
            .ce(N__31393),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_22_22_3.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_22_22_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_22_22_3.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_5_LC_22_22_3 (
            .in0(N__31492),
            .in1(N__29952),
            .in2(_gnd_net_),
            .in3(N__29945),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36947),
            .ce(N__31393),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_22_22_4.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_22_22_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_22_22_4.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_6_LC_22_22_4 (
            .in0(N__29925),
            .in1(N__31493),
            .in2(_gnd_net_),
            .in3(N__29918),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36947),
            .ce(N__31393),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_4_LC_23_5_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_4_LC_23_5_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_4_LC_23_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_4_LC_23_5_0  (
            .in0(_gnd_net_),
            .in1(N__30249),
            .in2(_gnd_net_),
            .in3(N__35699),
            .lcout(M_this_oam_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_7_LC_23_5_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_7_LC_23_5_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_7_LC_23_5_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_7_LC_23_5_2  (
            .in0(_gnd_net_),
            .in1(N__29886),
            .in2(_gnd_net_),
            .in3(N__35700),
            .lcout(M_this_oam_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_8_LC_23_5_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_8_LC_23_5_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_8_LC_23_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a4_8_LC_23_5_4  (
            .in0(_gnd_net_),
            .in1(N__30867),
            .in2(_gnd_net_),
            .in3(N__35701),
            .lcout(M_this_oam_ram_write_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_0_LC_23_5_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_0_LC_23_5_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_0_LC_23_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_0_LC_23_5_6  (
            .in0(_gnd_net_),
            .in1(N__30243),
            .in2(_gnd_net_),
            .in3(N__35698),
            .lcout(M_this_oam_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_4_LC_23_6_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_4_LC_23_6_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_4_LC_23_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_4_LC_23_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32448),
            .lcout(M_this_data_tmp_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36855),
            .ce(N__30237),
            .sr(N__36026));
    defparam M_this_data_tmp_q_esr_0_LC_23_6_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_0_LC_23_6_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_0_LC_23_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_0_LC_23_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31361),
            .lcout(M_this_data_tmp_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36855),
            .ce(N__30237),
            .sr(N__36026));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_3_LC_23_7_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_3_LC_23_7_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_3_LC_23_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_3_LC_23_7_3  (
            .in0(N__35630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30174),
            .lcout(M_this_oam_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_10_LC_23_7_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_10_LC_23_7_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_10_LC_23_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_10_LC_23_7_4  (
            .in0(_gnd_net_),
            .in1(N__30138),
            .in2(_gnd_net_),
            .in3(N__35629),
            .lcout(M_this_oam_ram_write_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_10_LC_23_8_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_10_LC_23_8_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_10_LC_23_8_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_10_LC_23_8_1 (
            .in0(N__35203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36867),
            .ce(N__36143),
            .sr(N__36021));
    defparam M_this_data_tmp_q_esr_12_LC_23_8_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_12_LC_23_8_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_12_LC_23_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_12_LC_23_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32444),
            .lcout(M_this_data_tmp_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36867),
            .ce(N__36143),
            .sr(N__36021));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_11_LC_23_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_11_LC_23_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_11_LC_23_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a4_11_LC_23_9_5  (
            .in0(_gnd_net_),
            .in1(N__30042),
            .in2(_gnd_net_),
            .in3(N__35642),
            .lcout(M_this_oam_ram_write_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNIOKR51_5_LC_23_9_7.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIOKR51_5_LC_23_9_7.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIOKR51_5_LC_23_9_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_this_oam_address_q_RNIOKR51_5_LC_23_9_7 (
            .in0(N__30110),
            .in1(N__30077),
            .in2(_gnd_net_),
            .in3(N__30764),
            .lcout(un1_M_this_oam_address_q_c6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_11_LC_23_10_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_11_LC_23_10_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_11_LC_23_10_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_11_LC_23_10_6 (
            .in0(N__35864),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36880),
            .ce(N__36141),
            .sr(N__36013));
    defparam M_this_data_tmp_q_esr_8_LC_23_11_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_8_LC_23_11_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_8_LC_23_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_8_LC_23_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31303),
            .lcout(M_this_data_tmp_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36888),
            .ce(N__36128),
            .sr(N__36010));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_0_a2_1_a2_LC_23_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_0_a2_1_a2_LC_23_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_0_a2_1_a2_LC_23_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_0_a2_1_a2_LC_23_12_6  (
            .in0(N__30811),
            .in1(N__30557),
            .in2(_gnd_net_),
            .in3(N__30667),
            .lcout(M_this_oam_ram_write_data_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNILNG41_3_LC_23_13_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNILNG41_3_LC_23_13_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNILNG41_3_LC_23_13_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_this_oam_address_q_RNILNG41_3_LC_23_13_4 (
            .in0(N__30727),
            .in1(N__30690),
            .in2(_gnd_net_),
            .in3(N__30505),
            .lcout(un1_M_this_oam_address_q_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_3_LC_23_14_4.C_ON=1'b0;
    defparam M_this_oam_address_q_3_LC_23_14_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_3_LC_23_14_4.LUT_INIT=16'b0000011000001100;
    LogicCell40 M_this_oam_address_q_3_LC_23_14_4 (
            .in0(N__30507),
            .in1(N__30728),
            .in2(N__33251),
            .in3(N__30692),
            .lcout(M_this_oam_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36908),
            .ce(),
            .sr(N__32215));
    defparam M_this_oam_address_q_2_LC_23_14_5.C_ON=1'b0;
    defparam M_this_oam_address_q_2_LC_23_14_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_2_LC_23_14_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_2_LC_23_14_5 (
            .in0(N__30691),
            .in1(N__33240),
            .in2(_gnd_net_),
            .in3(N__30506),
            .lcout(M_this_oam_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36908),
            .ce(),
            .sr(N__32215));
    defparam M_this_oam_address_q_RNIMU531_1_LC_23_16_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIMU531_1_LC_23_16_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIMU531_1_LC_23_16_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNIMU531_1_LC_23_16_4 (
            .in0(N__30665),
            .in1(N__30606),
            .in2(N__30548),
            .in3(N__31106),
            .lcout(un1_M_this_oam_address_q_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_23_19_2.C_ON=1'b0;
    defparam M_this_state_q_7_LC_23_19_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_23_19_2.LUT_INIT=16'b1111111111111000;
    LogicCell40 M_this_state_q_7_LC_23_19_2 (
            .in0(N__30374),
            .in1(N__30481),
            .in2(N__30459),
            .in3(N__30443),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36938),
            .ce(),
            .sr(N__36006));
    defparam M_this_state_q_0_LC_23_19_6.C_ON=1'b0;
    defparam M_this_state_q_0_LC_23_19_6.SEQ_MODE=4'b1001;
    defparam M_this_state_q_0_LC_23_19_6.LUT_INIT=16'b0101011100000011;
    LogicCell40 M_this_state_q_0_LC_23_19_6 (
            .in0(N__30327),
            .in1(N__30312),
            .in2(N__30300),
            .in3(N__30284),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36938),
            .ce(),
            .sr(N__36006));
    defparam \this_vga_signals.M_this_external_address_q_3_i_i_14_LC_23_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_i_i_14_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_i_i_14_LC_23_20_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_i_i_14_LC_23_20_1  (
            .in0(N__31677),
            .in1(N__35038),
            .in2(N__34424),
            .in3(N__31707),
            .lcout(N_312_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0_12_LC_23_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0_12_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0_12_LC_23_20_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0_12_LC_23_20_2  (
            .in0(N__36284),
            .in1(N__31209),
            .in2(_gnd_net_),
            .in3(N__36093),
            .lcout(\this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12 ),
            .ltout(\this_vga_signals.M_this_external_address_q_3_0_0_a4_0_0Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_12_LC_23_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_12_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_12_LC_23_20_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_0_0_12_LC_23_20_3  (
            .in0(N__32406),
            .in1(N__31671),
            .in2(N__31656),
            .in3(N__35040),
            .lcout(M_this_external_address_q_3_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3L4_LC_23_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3L4_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3L4_LC_23_20_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3L4_LC_23_20_6  (
            .in0(N__31589),
            .in1(N__31562),
            .in2(_gnd_net_),
            .in3(N__31531),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_3LZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_3_i_0_0_15_LC_23_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_i_0_0_15_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_i_0_0_15_LC_23_20_7 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_i_0_0_15_LC_23_20_7  (
            .in0(N__36094),
            .in1(N__34552),
            .in2(N__31215),
            .in3(N__31119),
            .lcout(this_vga_signals_M_this_external_address_q_3_i_0_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_23_21_5.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_23_21_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_23_21_5.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_7_LC_23_21_5 (
            .in0(N__31506),
            .in1(N__31494),
            .in2(_gnd_net_),
            .in3(N__31420),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36948),
            .ce(N__31401),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_8_LC_23_22_4.C_ON=1'b0;
    defparam M_this_external_address_q_8_LC_23_22_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_23_22_4.LUT_INIT=16'b1110001000100010;
    LogicCell40 M_this_external_address_q_8_LC_23_22_4 (
            .in0(N__36495),
            .in1(N__37107),
            .in2(N__31360),
            .in3(N__35035),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36951),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_a2_12_LC_23_22_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_a2_12_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_a2_12_LC_23_22_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_0_0_a2_12_LC_23_22_5  (
            .in0(N__31184),
            .in1(N__36091),
            .in2(_gnd_net_),
            .in3(N__31107),
            .lcout(N_760),
            .ltout(N_760_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_11_LC_23_22_6.C_ON=1'b0;
    defparam M_this_external_address_q_11_LC_23_22_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_23_22_6.LUT_INIT=16'b1011001110000000;
    LogicCell40 M_this_external_address_q_11_LC_23_22_6 (
            .in0(N__35839),
            .in1(N__37106),
            .in2(N__30870),
            .in3(N__36372),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36951),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_12_LC_23_22_7.C_ON=1'b0;
    defparam M_this_external_address_q_12_LC_23_22_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_23_22_7.LUT_INIT=16'b0001010010111110;
    LogicCell40 M_this_external_address_q_12_LC_23_22_7 (
            .in0(N__37105),
            .in1(N__37317),
            .in2(N__37343),
            .in3(N__31938),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36951),
            .ce(N__36561),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_23_25_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_23_25_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_23_25_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_5_0_wclke_3_LC_23_25_7  (
            .in0(N__34993),
            .in1(N__34910),
            .in2(N__34830),
            .in3(N__34682),
            .lcout(\this_sprites_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_24_5_0 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_24_5_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc2_LC_24_5_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc2_LC_24_5_0  (
            .in0(N__31737),
            .in1(N__31831),
            .in2(_gnd_net_),
            .in3(N__31797),
            .lcout(\this_ppu.un1_M_haddress_q_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_13_LC_24_5_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_13_LC_24_5_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_13_LC_24_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_13_LC_24_5_3  (
            .in0(N__36159),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35705),
            .lcout(M_this_oam_ram_write_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_15_LC_24_5_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_15_LC_24_5_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_15_LC_24_5_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_15_LC_24_5_4  (
            .in0(N__35706),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34467),
            .lcout(M_this_oam_ram_write_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_24_5_5 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_24_5_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc4_LC_24_5_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc4_LC_24_5_5  (
            .in0(N__31763),
            .in1(N__31739),
            .in2(N__31871),
            .in3(N__31776),
            .lcout(\this_ppu.un1_M_haddress_q_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_24_5_6 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_24_5_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_ac0_1_LC_24_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_ac0_1_LC_24_5_6  (
            .in0(_gnd_net_),
            .in1(N__31830),
            .in2(_gnd_net_),
            .in3(N__31796),
            .lcout(\this_ppu.un1_oam_data_1_c2 ),
            .ltout(\this_ppu.un1_oam_data_1_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_5_7 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_5_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_axbxc3_LC_24_5_7 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \this_ppu.un1_oam_data_1_axbxc3_LC_24_5_7  (
            .in0(_gnd_net_),
            .in1(N__31762),
            .in2(N__31746),
            .in3(N__31738),
            .lcout(\this_ppu.un1_M_haddress_q_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_12_LC_24_6_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_12_LC_24_6_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_12_LC_24_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_12_LC_24_6_3  (
            .in0(_gnd_net_),
            .in1(N__32157),
            .in2(_gnd_net_),
            .in3(N__35702),
            .lcout(M_this_oam_ram_write_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_6_4 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_6_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_axbxc2_LC_24_6_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.un1_oam_data_axbxc2_LC_24_6_4  (
            .in0(N__32128),
            .in1(N__32097),
            .in2(_gnd_net_),
            .in3(N__32063),
            .lcout(\this_ppu.un1_M_vaddress_q_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_5_LC_24_6_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_5_LC_24_6_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_5_LC_24_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_5_LC_24_6_5  (
            .in0(_gnd_net_),
            .in1(N__32022),
            .in2(_gnd_net_),
            .in3(N__35703),
            .lcout(M_this_oam_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_6_6 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_6_6 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31984),
            .lcout(M_this_oam_ram_read_data_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_9_LC_24_6_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_9_LC_24_6_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_9_LC_24_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a4_9_LC_24_6_7  (
            .in0(_gnd_net_),
            .in1(N__32166),
            .in2(_gnd_net_),
            .in3(N__35704),
            .lcout(M_this_oam_ram_write_data_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_18_LC_24_7_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_18_LC_24_7_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_18_LC_24_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_18_LC_24_7_0  (
            .in0(_gnd_net_),
            .in1(N__32460),
            .in2(_gnd_net_),
            .in3(N__35695),
            .lcout(M_this_oam_ram_write_data_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_20_LC_24_7_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_20_LC_24_7_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_20_LC_24_7_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_20_LC_24_7_1  (
            .in0(N__35696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32454),
            .lcout(M_this_oam_ram_write_data_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_29_LC_24_7_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_29_LC_24_7_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_29_LC_24_7_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_29_LC_24_7_2  (
            .in0(N__36301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35692),
            .lcout(M_this_oam_ram_write_data_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_30_LC_24_7_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_30_LC_24_7_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_30_LC_24_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_30_LC_24_7_3  (
            .in0(N__35693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34417),
            .lcout(M_this_oam_ram_write_data_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_22_LC_24_7_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_22_LC_24_7_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_22_LC_24_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_22_LC_24_7_4  (
            .in0(_gnd_net_),
            .in1(N__32487),
            .in2(_gnd_net_),
            .in3(N__35697),
            .lcout(M_this_oam_ram_write_data_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_31_LC_24_7_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_31_LC_24_7_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_31_LC_24_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_31_LC_24_7_7  (
            .in0(N__35694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34529),
            .lcout(M_this_oam_ram_write_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_18_LC_24_8_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_18_LC_24_8_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_18_LC_24_8_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_18_LC_24_8_1 (
            .in0(N__35234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36873),
            .ce(N__34020),
            .sr(N__36017));
    defparam M_this_data_tmp_q_esr_20_LC_24_8_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_20_LC_24_8_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_20_LC_24_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_20_LC_24_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32442),
            .lcout(M_this_data_tmp_qZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36873),
            .ce(N__34020),
            .sr(N__36017));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_28_LC_24_8_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_28_LC_24_8_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_28_LC_24_8_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_28_LC_24_8_6  (
            .in0(N__32443),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35643),
            .lcout(M_this_oam_ram_write_data_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_21_LC_24_8_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_21_LC_24_8_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_21_LC_24_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_21_LC_24_8_7  (
            .in0(N__35644),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32289),
            .lcout(M_this_oam_ram_write_data_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_6_LC_24_9_0.C_ON=1'b0;
    defparam M_this_oam_address_q_6_LC_24_9_0.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_6_LC_24_9_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_6_LC_24_9_0 (
            .in0(N__32266),
            .in1(N__33245),
            .in2(_gnd_net_),
            .in3(N__32249),
            .lcout(M_this_oam_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36881),
            .ce(),
            .sr(N__32216));
    defparam M_this_oam_address_q_7_LC_24_9_2.C_ON=1'b0;
    defparam M_this_oam_address_q_7_LC_24_9_2.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_7_LC_24_9_2.LUT_INIT=16'b0001001000110000;
    LogicCell40 M_this_oam_address_q_7_LC_24_9_2 (
            .in0(N__32267),
            .in1(N__33246),
            .in2(N__32237),
            .in3(N__32250),
            .lcout(M_this_oam_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36881),
            .ce(),
            .sr(N__32216));
    defparam M_this_data_tmp_q_esr_9_LC_24_10_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_9_LC_24_10_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_9_LC_24_10_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_9_LC_24_10_6 (
            .in0(N__33371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36889),
            .ce(N__36142),
            .sr(N__36011));
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_11_0 .C_ON=1'b1;
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_11_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_11_0  (
            .in0(_gnd_net_),
            .in1(N__33153),
            .in2(N__34307),
            .in3(N__32793),
            .lcout(\this_ppu.M_this_oam_ram_read_data_iZ0Z_8 ),
            .ltout(),
            .carryin(bfn_24_11_0_),
            .carryout(\this_ppu.un2_hscroll_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_11_1 .C_ON=1'b1;
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_11_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(N__33147),
            .in2(N__33066),
            .in3(N__33138),
            .lcout(\this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0 ),
            .ltout(),
            .carryin(\this_ppu.un2_hscroll_cry_0 ),
            .carryout(\this_ppu.un2_hscroll_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_11_2 .C_ON=1'b0;
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_11_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_11_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_11_2  (
            .in0(N__33131),
            .in1(N__32739),
            .in2(_gnd_net_),
            .in3(N__33093),
            .lcout(\this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_26_LC_24_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_26_LC_24_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_26_LC_24_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_26_LC_24_11_6  (
            .in0(_gnd_net_),
            .in1(N__35168),
            .in2(_gnd_net_),
            .in3(N__35540),
            .lcout(M_this_oam_ram_write_data_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_19_LC_24_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_19_LC_24_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a4_19_LC_24_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a4_19_LC_24_11_7  (
            .in0(N__35541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34029),
            .lcout(M_this_oam_ram_write_data_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI0O061_1_LC_24_12_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI0O061_1_LC_24_12_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI0O061_1_LC_24_12_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \this_ppu.M_haddress_q_RNI0O061_1_LC_24_12_1  (
            .in0(N__33790),
            .in1(N__33064),
            .in2(N__33933),
            .in3(N__32994),
            .lcout(M_this_ppu_sprites_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_24_12_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_24_12_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI88B5_0_LC_24_12_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_ppu.M_haddress_q_RNI88B5_0_LC_24_12_2  (
            .in0(N__32794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34301),
            .lcout(\this_ppu.un2_hscroll_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI3S161_2_LC_24_13_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI3S161_2_LC_24_13_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI3S161_2_LC_24_13_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \this_ppu.M_haddress_q_RNI3S161_2_LC_24_13_0  (
            .in0(N__33775),
            .in1(N__33917),
            .in2(N__32747),
            .in3(N__32670),
            .lcout(M_this_ppu_sprites_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIRG7O_0_LC_24_13_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIRG7O_0_LC_24_13_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIRG7O_0_LC_24_13_5 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \this_ppu.M_haddress_q_RNIRG7O_0_LC_24_13_5  (
            .in0(N__34320),
            .in1(N__33774),
            .in2(N__33932),
            .in3(N__34302),
            .lcout(M_this_ppu_sprites_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_19_LC_24_14_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_19_LC_24_14_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_19_LC_24_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_19_LC_24_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35848),
            .lcout(M_this_data_tmp_qZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36916),
            .ce(N__34005),
            .sr(N__36007));
    defparam \this_ppu.M_state_q_RNI0VTU_2_4_LC_24_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI0VTU_2_4_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI0VTU_2_4_LC_24_15_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \this_ppu.M_state_q_RNI0VTU_2_4_LC_24_15_6  (
            .in0(N__33975),
            .in1(N__33960),
            .in2(N__33931),
            .in3(N__33791),
            .lcout(M_this_ppu_sprites_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_17_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_17_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_17_3  (
            .in0(N__34996),
            .in1(N__34905),
            .in2(N__34832),
            .in3(N__34709),
            .lcout(\this_sprites_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_17_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_17_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_17_4  (
            .in0(N__34710),
            .in1(N__34821),
            .in2(N__34913),
            .in3(N__34997),
            .lcout(\this_sprites_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_18_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_18_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_18_7  (
            .in0(N__34998),
            .in1(N__34889),
            .in2(N__34833),
            .in3(N__34708),
            .lcout(\this_sprites_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_9_LC_24_19_3.C_ON=1'b0;
    defparam M_this_external_address_q_9_LC_24_19_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_24_19_3.LUT_INIT=16'b1010000011001100;
    LogicCell40 M_this_external_address_q_9_LC_24_19_3 (
            .in0(N__35039),
            .in1(N__36453),
            .in2(N__33400),
            .in3(N__37116),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36944),
            .ce(N__36560),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_15_LC_24_19_6.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_24_19_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_24_19_6.LUT_INIT=16'b0101000011011000;
    LogicCell40 M_this_external_address_q_15_LC_24_19_6 (
            .in0(N__37115),
            .in1(N__33267),
            .in2(N__37176),
            .in3(N__33244),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36944),
            .ce(N__36560),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_20_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_20_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_20_5  (
            .in0(N__34906),
            .in1(N__34991),
            .in2(N__34828),
            .in3(N__34693),
            .lcout(\this_sprites_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_13_LC_24_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_13_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_external_address_q_3_0_0_13_LC_24_20_7 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \this_vga_signals.M_this_external_address_q_3_0_0_13_LC_24_20_7  (
            .in0(N__36259),
            .in1(N__35037),
            .in2(_gnd_net_),
            .in3(N__35361),
            .lcout(M_this_external_address_q_3_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4L6_LC_24_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4L6_LC_24_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4L6_LC_24_21_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4L6_LC_24_21_1  (
            .in0(N__35285),
            .in1(N__35270),
            .in2(N__35307),
            .in3(N__35352),
            .lcout(\this_vga_signals.M_this_state_q_ns_0_i_0_0_a4_0_N_4LZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_4_LC_24_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_4_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_this_state_q_19_i_0_o2_4_LC_24_21_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.un1_M_this_state_q_19_i_0_o2_4_LC_24_21_5  (
            .in0(N__35327),
            .in1(N__35306),
            .in2(N__35289),
            .in3(N__35271),
            .lcout(\this_vga_signals.un1_M_this_state_q_19_i_0_o2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_10_LC_24_22_3.C_ON=1'b0;
    defparam M_this_external_address_q_10_LC_24_22_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_24_22_3.LUT_INIT=16'b1110010001000100;
    LogicCell40 M_this_external_address_q_10_LC_24_22_3 (
            .in0(N__37114),
            .in1(N__36411),
            .in2(N__35172),
            .in3(N__35036),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36954),
            .ce(N__36576),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_25_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_25_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_25_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_25_5  (
            .in0(N__34992),
            .in1(N__34911),
            .in2(N__34829),
            .in3(N__34683),
            .lcout(\this_sprites_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_14_LC_26_5_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_14_LC_26_5_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_14_LC_26_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_14_LC_26_5_3  (
            .in0(_gnd_net_),
            .in1(N__34329),
            .in2(_gnd_net_),
            .in3(N__35691),
            .lcout(M_this_oam_ram_write_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_15_LC_26_7_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_15_LC_26_7_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_15_LC_26_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_15_LC_26_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34513),
            .lcout(M_this_data_tmp_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36882),
            .ce(N__36147),
            .sr(N__36014));
    defparam M_this_data_tmp_q_esr_14_LC_26_7_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_14_LC_26_7_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_14_LC_26_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_14_LC_26_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34391),
            .lcout(M_this_data_tmp_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36882),
            .ce(N__36147),
            .sr(N__36014));
    defparam M_this_data_tmp_q_esr_13_LC_26_7_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_13_LC_26_7_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_13_LC_26_7_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_13_LC_26_7_5 (
            .in0(N__36300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36882),
            .ce(N__36147),
            .sr(N__36014));
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_27_LC_26_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_27_LC_26_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_27_LC_26_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_oam_ram_write_data_0_a3_0_a4_27_LC_26_9_2  (
            .in0(_gnd_net_),
            .in1(N__35838),
            .in2(_gnd_net_),
            .in3(N__35641),
            .lcout(M_this_oam_ram_write_data_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_13_LC_26_20_5.C_ON=1'b0;
    defparam M_this_external_address_q_13_LC_26_20_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_26_20_5.LUT_INIT=16'b0001010010111110;
    LogicCell40 M_this_external_address_q_13_LC_26_20_5 (
            .in0(N__37113),
            .in1(N__37272),
            .in2(N__37298),
            .in3(N__35502),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36957),
            .ce(N__36574),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_14_LC_26_20_7.C_ON=1'b0;
    defparam M_this_external_address_q_14_LC_26_20_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_26_20_7.LUT_INIT=16'b0001010010111110;
    LogicCell40 M_this_external_address_q_14_LC_26_20_7 (
            .in0(N__37112),
            .in1(N__37227),
            .in2(N__37253),
            .in3(N__35493),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36957),
            .ce(N__36574),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_0_LC_26_21_0.C_ON=1'b1;
    defparam M_this_external_address_q_0_LC_26_21_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_26_21_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_0_LC_26_21_0 (
            .in0(N__37108),
            .in1(N__35471),
            .in2(_gnd_net_),
            .in3(N__35460),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_26_21_0_),
            .carryout(M_this_external_address_q_cry_0),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_1_LC_26_21_1.C_ON=1'b1;
    defparam M_this_external_address_q_1_LC_26_21_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_26_21_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_1_LC_26_21_1 (
            .in0(N__37079),
            .in1(N__35450),
            .in2(_gnd_net_),
            .in3(N__35439),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(M_this_external_address_q_cry_0),
            .carryout(M_this_external_address_q_cry_1),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_2_LC_26_21_2.C_ON=1'b1;
    defparam M_this_external_address_q_2_LC_26_21_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_26_21_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_2_LC_26_21_2 (
            .in0(N__37109),
            .in1(N__35423),
            .in2(_gnd_net_),
            .in3(N__35412),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(M_this_external_address_q_cry_1),
            .carryout(M_this_external_address_q_cry_2),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_3_LC_26_21_3.C_ON=1'b1;
    defparam M_this_external_address_q_3_LC_26_21_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_26_21_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_3_LC_26_21_3 (
            .in0(N__37080),
            .in1(N__35396),
            .in2(_gnd_net_),
            .in3(N__35385),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(M_this_external_address_q_cry_2),
            .carryout(M_this_external_address_q_cry_3),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_4_LC_26_21_4.C_ON=1'b1;
    defparam M_this_external_address_q_4_LC_26_21_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_26_21_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_4_LC_26_21_4 (
            .in0(N__37110),
            .in1(N__35372),
            .in2(_gnd_net_),
            .in3(N__37161),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(M_this_external_address_q_cry_3),
            .carryout(M_this_external_address_q_cry_4),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_5_LC_26_21_5.C_ON=1'b1;
    defparam M_this_external_address_q_5_LC_26_21_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_26_21_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_5_LC_26_21_5 (
            .in0(N__37081),
            .in1(N__37154),
            .in2(_gnd_net_),
            .in3(N__37143),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(M_this_external_address_q_cry_4),
            .carryout(M_this_external_address_q_cry_5),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_6_LC_26_21_6.C_ON=1'b1;
    defparam M_this_external_address_q_6_LC_26_21_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_26_21_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_6_LC_26_21_6 (
            .in0(N__37111),
            .in1(N__37130),
            .in2(_gnd_net_),
            .in3(N__37119),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(M_this_external_address_q_cry_5),
            .carryout(M_this_external_address_q_cry_6),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_7_LC_26_21_7.C_ON=1'b1;
    defparam M_this_external_address_q_7_LC_26_21_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_26_21_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_7_LC_26_21_7 (
            .in0(N__37082),
            .in1(N__36992),
            .in2(_gnd_net_),
            .in3(N__36981),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(M_this_external_address_q_cry_6),
            .carryout(M_this_external_address_q_cry_7),
            .clk(N__36958),
            .ce(N__36575),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_8_LC_26_22_0.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_8_LC_26_22_0.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_8_LC_26_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_8_LC_26_22_0 (
            .in0(_gnd_net_),
            .in1(N__36512),
            .in2(_gnd_net_),
            .in3(N__36486),
            .lcout(M_this_external_address_q_s_8),
            .ltout(),
            .carryin(bfn_26_22_0_),
            .carryout(M_this_external_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_9_LC_26_22_1.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_9_LC_26_22_1.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_9_LC_26_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_9_LC_26_22_1 (
            .in0(_gnd_net_),
            .in1(N__36476),
            .in2(_gnd_net_),
            .in3(N__36441),
            .lcout(M_this_external_address_q_s_9),
            .ltout(),
            .carryin(M_this_external_address_q_cry_8),
            .carryout(M_this_external_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_10_LC_26_22_2.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_10_LC_26_22_2.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_10_LC_26_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_10_LC_26_22_2 (
            .in0(_gnd_net_),
            .in1(N__36428),
            .in2(_gnd_net_),
            .in3(N__36402),
            .lcout(M_this_external_address_q_s_10),
            .ltout(),
            .carryin(M_this_external_address_q_cry_9),
            .carryout(M_this_external_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_11_LC_26_22_3.C_ON=1'b1;
    defparam M_this_external_address_q_RNO_0_11_LC_26_22_3.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_11_LC_26_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_external_address_q_RNO_0_11_LC_26_22_3 (
            .in0(_gnd_net_),
            .in1(N__36386),
            .in2(_gnd_net_),
            .in3(N__36363),
            .lcout(M_this_external_address_q_s_11),
            .ltout(),
            .carryin(M_this_external_address_q_cry_10),
            .carryout(M_this_external_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_22_4.C_ON=1'b1;
    defparam M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_22_4.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_22_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_external_address_q_cry_11_THRU_LUT4_0_LC_26_22_4 (
            .in0(_gnd_net_),
            .in1(N__37342),
            .in2(_gnd_net_),
            .in3(N__37308),
            .lcout(M_this_external_address_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(M_this_external_address_q_cry_11),
            .carryout(M_this_external_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_22_5.C_ON=1'b1;
    defparam M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_22_5.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_22_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_external_address_q_cry_12_THRU_LUT4_0_LC_26_22_5 (
            .in0(_gnd_net_),
            .in1(N__37297),
            .in2(_gnd_net_),
            .in3(N__37263),
            .lcout(M_this_external_address_q_cry_12_THRU_CO),
            .ltout(),
            .carryin(M_this_external_address_q_cry_12),
            .carryout(M_this_external_address_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_22_6.C_ON=1'b1;
    defparam M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_22_6.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_22_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_external_address_q_cry_13_THRU_LUT4_0_LC_26_22_6 (
            .in0(_gnd_net_),
            .in1(N__37252),
            .in2(_gnd_net_),
            .in3(N__37218),
            .lcout(M_this_external_address_q_cry_13_THRU_CO),
            .ltout(),
            .carryin(M_this_external_address_q_cry_13),
            .carryout(M_this_external_address_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_RNO_0_15_LC_26_22_7.C_ON=1'b0;
    defparam M_this_external_address_q_RNO_0_15_LC_26_22_7.SEQ_MODE=4'b0000;
    defparam M_this_external_address_q_RNO_0_15_LC_26_22_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_this_external_address_q_RNO_0_15_LC_26_22_7 (
            .in0(_gnd_net_),
            .in1(N__37202),
            .in2(_gnd_net_),
            .in3(N__37179),
            .lcout(M_this_external_address_q_s_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
