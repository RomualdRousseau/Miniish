-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 3 2022 11:35:56

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : in std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : in std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    debug : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_rw_c_i : std_logic;
signal port_nmib_c_i : std_logic;
signal \this_vga_signals.N_29_cascade_\ : std_logic;
signal \this_vga_signals.N_40_cascade_\ : std_logic;
signal \this_vga_signals.N_20\ : std_logic;
signal \this_vga_signals.N_18_cascade_\ : std_logic;
signal \this_vga_signals_N_274_i\ : std_logic;
signal \this_vga_signals.hvisible_i_a2_0_3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_1\ : std_logic;
signal \this_vga_signals.N_49_cascade_\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_vga_signals.N_32\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_0\ : std_logic;
signal \this_vga_signals.N_26\ : std_logic;
signal \this_vga_signals.N_26_cascade_\ : std_logic;
signal \this_vga_signals.N_51\ : std_logic;
signal \this_vga_signals.N_273\ : std_logic;
signal \this_vga_signals.N_2_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.N_70_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.m44_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNIQE2J1Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_RNI3BJLZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_2_cascade_\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_7\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_9\ : std_logic;
signal \this_vga_signals.M_hstate_d_0_sqmuxa\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_10\ : std_logic;
signal \this_vga_signals.g1_0_0_a2_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_11_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KANZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.N_2\ : std_logic;
signal \this_vga_signals.i9_mux_cascade_\ : std_logic;
signal \this_vga_signals.i9_mux\ : std_logic;
signal \this_vga_signals.address_1_c5_i\ : std_logic;
signal port_nmib_c : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCNZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_vga_signals.address_1_c4_cascade_\ : std_logic;
signal \this_vga_signals.N_70\ : std_logic;
signal \this_vga_signals.SUM_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_c\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axbxc1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.N_13_0\ : std_logic;
signal \this_vga_signals.if_i1_mux\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNO_0Z0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.address_m24_ns_1Z0Z_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNO_0Z0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.un12_address_cry_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un12_address_cry_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un12_address_cry_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un12_address_cry_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un12_address_cry_4\ : std_logic;
signal \this_vga_signals.un12_address_cry_5\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.un12_address_cry_6\ : std_logic;
signal \this_vga_signals.un12_address_cry_7\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \this_vga_signals.un12_address_cry_8\ : std_logic;
signal \this_vga_signals.un12_address_cry_9\ : std_logic;
signal \this_vga_signals.un12_address_cry_10\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.N_49\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_11\ : std_logic;
signal \N_16\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_7_0_3_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_7_0_3_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.N_27\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.hvisible_i_a2_2_0\ : std_logic;
signal rgb_c_4 : std_logic;
signal \this_vga_signals.m30_3\ : std_logic;
signal \this_vga_signals.m30_4_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.N_3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal rgb_c_0 : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.address_m1_1_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2\ : std_logic;
signal \this_vga_signals.address_i3_mux_i\ : std_logic;
signal \this_vga_signals.address_m27_ns_1_cascade_\ : std_logic;
signal \this_vga_signals.address_i2_mux_3_cascade_\ : std_logic;
signal \this_vga_signals.address_i2_mux_2\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNO_0Z0Z_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_8_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_10\ : std_logic;
signal \this_vga_signals.M_hcounter_q_i_11\ : std_logic;
signal \this_vga_signals.un12_address_cry_9_THRU_CO\ : std_logic;
signal \this_vga_signals.un12_address_cry_9_c_RNIVF1R\ : std_logic;
signal \this_vga_signals.un12_address_cry_10_c_RNINP5K\ : std_logic;
signal \this_vga_signals.un12_address_cry_9_c_RNIVF1R_cascade_\ : std_logic;
signal \this_vga_signals.un12_address_cry_9_c_RNIEJOE\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb3_x1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb3_cascade_\ : std_logic;
signal \this_vga_signals.if_m5_sn\ : std_logic;
signal \this_vga_signals.if_m5_rn_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c5_cascade_\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_7_0_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_7_0_4_cascade_\ : std_logic;
signal \this_vga_signals.if_m4_0_1_cascade_\ : std_logic;
signal \this_vga_signals.G_12_0_x3_0_cascade_\ : std_logic;
signal vsync_c : std_logic;
signal \this_vga_signals.N_52_cascade_\ : std_logic;
signal \this_vga_signals.N_76_mux\ : std_logic;
signal \this_vga_signals.N_76_mux_cascade_\ : std_logic;
signal \this_vga_signals.N_72_mux\ : std_logic;
signal \this_vga_signals.N_55_cascade_\ : std_logic;
signal \this_vga_signals.M_vstate_q_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vstate_q_RNO_2Z0Z_0\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_1\ : std_logic;
signal \this_vga_signals.m35_e_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c2\ : std_logic;
signal \this_vga_signals.address_N_9_0_cascade_\ : std_logic;
signal \this_vga_signals.address_N_10_0\ : std_logic;
signal \this_vga_signals.address_N_3\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNI8OSG6BZ0Z_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3\ : std_logic;
signal \this_vga_signals.address_m35_1\ : std_logic;
signal \this_vga_signals.N_75_mux\ : std_logic;
signal \this_vga_signals.N_84\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNO_0Z0Z_2\ : std_logic;
signal \this_vga_signals.address_m31_1\ : std_logic;
signal \this_vga_signals.address_i2_mux_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0\ : std_logic;
signal \this_vga_signals.address_N_9_0\ : std_logic;
signal \this_vga_signals.address_N_33_cascade_\ : std_logic;
signal \this_vga_signals.address_N_34\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb3_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_4_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb3_out\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb4\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c5\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb4_x0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_7_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb4_x1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb4_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb4_i\ : std_logic;
signal \this_vga_signals.g0_6_0_0_1\ : std_logic;
signal \this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb3\ : std_logic;
signal \this_vga_signals.if_m4_0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc5\ : std_logic;
signal \this_vga_signals.un12_address_cry_7_c_RNI32HB\ : std_logic;
signal \this_vga_signals.if_m2_3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb3_1\ : std_logic;
signal \this_vga_signals.G_12_0_3_1\ : std_logic;
signal \this_vga_signals.N_9_cascade_\ : std_logic;
signal \this_vga_signals.G_12_0_3_cascade_\ : std_logic;
signal \this_vga_signals.if_m4_0_1\ : std_logic;
signal \this_vga_signals_un17_address_if_N_8_mux_cascade_\ : std_logic;
signal \this_vga_signals.N_10_0\ : std_logic;
signal \N_6_i_cascade_\ : std_logic;
signal \this_vga_signals.N_18_0\ : std_logic;
signal \this_vga_signals.g0_6_1\ : std_logic;
signal \this_vga_signals.G_12_0_x3_0\ : std_logic;
signal \N_11_0_cascade_\ : std_logic;
signal \this_vga_signals.N_5_i\ : std_logic;
signal \this_vga_signals.G_12_0_1\ : std_logic;
signal \this_vga_signals.N_25\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.N_275\ : std_logic;
signal \this_vga_signals.if_N_9_i_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_\ : std_logic;
signal \M_this_vga_signals_address_8\ : std_logic;
signal \this_vga_signals.address_m6_0_1_cascade_\ : std_logic;
signal \this_vga_signals.address_mZ0Z1\ : std_logic;
signal \this_vga_signals.address_i2_mux_cascade_\ : std_logic;
signal \this_vga_signals.address_N_11\ : std_logic;
signal \this_vga_signals.address_i2_mux_0\ : std_logic;
signal \this_vga_signals.address_m21_ns_1_cascade_\ : std_logic;
signal \this_vga_signals.address_i2_mux_1\ : std_logic;
signal \this_vga_signals.address_N_22_cascade_\ : std_logic;
signal \this_vga_signals.address_N_36\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_0\ : std_logic;
signal \this_vga_signals.if_m16_0_o4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.address_N_40\ : std_logic;
signal \this_vga_signals.if_m4_0_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_3L3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_2L1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5_cascade_\ : std_logic;
signal \this_vga_signals.N_21_0\ : std_logic;
signal \this_vga_signals.g0_6_0_0_2\ : std_logic;
signal \this_vga_signals.if_N_8_mux_2_2\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axb3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_4\ : std_logic;
signal \this_vga_signals.g0_i_x4_4_a3_1\ : std_logic;
signal \this_vga_signals.if_m1_0\ : std_logic;
signal \this_vga_signals.if_N_3_3_i\ : std_logic;
signal \this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5_cascade_\ : std_logic;
signal \this_vga_signals.if_N_3_2_i_cascade_\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_7_0_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_5\ : std_logic;
signal \this_vga_signals.N_12\ : std_logic;
signal \this_vga_signals.g0_0_0_a2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_3_2_i_3_1_cascade_\ : std_logic;
signal \this_vga_signals.N_31\ : std_logic;
signal \this_vga_signals.N_20_i_i\ : std_logic;
signal \this_vga_signals.N_20_i_i_cascade_\ : std_logic;
signal \this_vga_signals.N_26_i_i\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0\ : std_logic;
signal \M_this_vga_signals_address_9\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_7\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_8\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vga_signals.N_4\ : std_logic;
signal \this_vram.M_this_vram_read_data_1_cascade_\ : std_logic;
signal rgb_c_2 : std_logic;
signal \this_vga_signals.g0_4\ : std_logic;
signal \this_vga_signals.if_N_8_mux_2_2_1\ : std_logic;
signal \this_vga_signals.N_3_1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_2_0_0\ : std_logic;
signal \this_vga_signals.g0_0_0_0\ : std_logic;
signal \this_vga_signals.if_m1_0_0\ : std_logic;
signal \this_vga_signals.N_21\ : std_logic;
signal \this_vga_signals.g0_3\ : std_logic;
signal \this_vga_signals.N_20_i_i_0\ : std_logic;
signal \this_vga_signals.g0_0_a3_3\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_7_0_1_0\ : std_logic;
signal \this_vga_signals.N_11_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_a3_2\ : std_logic;
signal \this_vga_signals.g0_0_a3_5_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_4_a3\ : std_logic;
signal \this_vga_signals.N_3_3_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_1\ : std_logic;
signal \this_vga_signals.g0_0_1_0\ : std_logic;
signal \this_vga_signals.g1_5_0_0_cascade_\ : std_logic;
signal \this_vga_signals.r_N_2_0_0_0\ : std_logic;
signal \this_vga_signals.g0_1_0\ : std_logic;
signal \this_vga_signals.g0_1_2_cascade_\ : std_logic;
signal \this_vga_signals_un17_address_if_N_8_mux\ : std_logic;
signal \this_vga_signals.g0_3_0_a2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_7_0_1_2\ : std_logic;
signal \this_vga_signals.if_N_8_mux_2_0\ : std_logic;
signal this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5 : std_logic;
signal \this_vga_signals.if_N_3_2_i\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0 : std_logic;
signal \this_vga_signals.g0_6_0\ : std_logic;
signal \this_vga_signals.g1_2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5\ : std_logic;
signal \this_vga_signals.g1_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb3\ : std_logic;
signal \this_vga_signals.g0_0_1_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_2_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0_0\ : std_logic;
signal \this_vga_signals.g0_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_7_0_1_4\ : std_logic;
signal \this_vga_signals.g0_6\ : std_logic;
signal \this_vga_signals.g0_13\ : std_logic;
signal \this_vga_signals.if_N_3_2_i_0\ : std_logic;
signal \this_vga_signals.g0_0_0_a2_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_0\ : std_logic;
signal \this_vga_signals.g1_2_cascade_\ : std_logic;
signal \this_vga_signals.r_N_2_0_0_2_cascade_\ : std_logic;
signal \this_vga_signals.N_3_1_1\ : std_logic;
signal \this_vga_signals.g0_3_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c5\ : std_logic;
signal \this_vga_signals.un12_address_cry_3_c_RNIRLCB\ : std_logic;
signal \this_vga_signals.g0_5_3_cascade_\ : std_logic;
signal \this_vga_signals.un12_address_cry_2_c_RNIPIBB\ : std_logic;
signal \this_vga_signals.un12_address_cry_1_c_RNINFAB\ : std_logic;
signal \this_vga_signals.mult1_un96_sum_c5_0_1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.N_3_1_2\ : std_logic;
signal \this_vga_signals.g1_0_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un96_sum_c5_cascade_\ : std_logic;
signal \this_vga_signals.g2_0\ : std_logic;
signal \this_vga_signals.mult1_un96_sum_axbxc5_2\ : std_logic;
signal \this_vga_signals.g1_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c5_0_0_0_0\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.if_N_3_2_i_1\ : std_logic;
signal \this_vga_signals.un12_address_cry_4_c_RNITODB\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc5\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_ac0_7_0_1_3\ : std_logic;
signal \this_vga_signals.un12_address_cry_5_c_RNIVREB\ : std_logic;
signal this_vga_signals_un17_address_if_m2_2_0 : std_logic;
signal \this_vga_signals.g0_38\ : std_logic;
signal \this_vga_signals.N_4_0_1\ : std_logic;
signal \this_vga_signals.if_N_3_2_i_2_0\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_0\ : std_logic;
signal port_clk_c : std_logic;
signal \this_start_data_delay_this_edge_detector_M_last_q\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_0\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_3\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_1\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_2\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_5\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_1\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_2\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_3\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_4\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_10\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_9\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_6\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_4\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1\ : std_logic;
signal \M_this_vga_signals_address_10\ : std_logic;
signal \this_vram.M_this_vram_read_data_0\ : std_logic;
signal \this_vram.N_17_0\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_11\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_12\ : std_logic;
signal debug_d : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_13\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_14\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_15\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_16\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_17\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_18\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_7\ : std_logic;
signal \this_start_data_delay.this_delay.M_pipe_qZ0Z_8\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_215\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_212\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_219\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_8\ : std_logic;
signal port_data_c_5 : std_logic;
signal \this_start_data_delay.this_edge_detector.N_222\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_6\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_7\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_9\ : std_logic;
signal \bfn_19_23_0_\ : std_logic;
signal \un1_M_current_address_q_cry_0\ : std_logic;
signal \M_current_address_qZ0Z_2\ : std_logic;
signal \un1_M_current_address_q_cry_1_c_RNI4TBNZ0\ : std_logic;
signal \un1_M_current_address_q_cry_1\ : std_logic;
signal \un1_M_current_address_q_cry_2\ : std_logic;
signal \un1_M_current_address_q_cry_3_c_RNI83ENZ0\ : std_logic;
signal \un1_M_current_address_q_cry_3\ : std_logic;
signal \M_current_address_qZ0Z_5\ : std_logic;
signal \un1_M_current_address_q_cry_4_c_RNIA6FNZ0\ : std_logic;
signal \un1_M_current_address_q_cry_4\ : std_logic;
signal \un1_M_current_address_q_cry_5\ : std_logic;
signal \un1_M_current_address_q_cry_6\ : std_logic;
signal \un1_M_current_address_q_cry_7\ : std_logic;
signal \un1_M_current_address_q_cry_7_c_RNIGFINZ0\ : std_logic;
signal \bfn_19_24_0_\ : std_logic;
signal \M_current_address_qZ0Z_9\ : std_logic;
signal \un1_M_current_address_q_cry_8_c_RNIIIJNZ0\ : std_logic;
signal \un1_M_current_address_q_cry_8\ : std_logic;
signal \un1_M_current_address_q_cry_9\ : std_logic;
signal \un1_M_current_address_q_cry_10\ : std_logic;
signal \un1_M_current_address_q_cry_11_c_RNI6NLHZ0\ : std_logic;
signal \un1_M_current_address_q_cry_11\ : std_logic;
signal \un1_M_current_address_q_cry_12\ : std_logic;
signal \N_177_0\ : std_logic;
signal \un1_M_current_address_q_cry_9_c_RNIRDIMZ0\ : std_logic;
signal \un1_M_current_address_q_cry_0_c_RNI2QANZ0\ : std_logic;
signal \un1_M_current_address_q_cry_12_c_RNI8QMHZ0\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_12\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_10\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_11\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_13\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_14\ : std_logic;
signal \M_current_address_q_RNIHDTUZ0Z_0\ : std_logic;
signal \un1_M_current_address_q_cry_5_c_RNIC9GNZ0\ : std_logic;
signal \un1_M_current_address_q_cry_6_c_RNIECHNZ0\ : std_logic;
signal \un1_M_current_address_q_cry_10_c_RNI4KKHZ0\ : std_logic;
signal \un1_M_current_address_q_cry_2_c_RNI60DNZ0\ : std_logic;
signal \N_339_g\ : std_logic;
signal \M_current_address_qZ0Z_6\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_216\ : std_logic;
signal \M_current_address_qZ0Z_3\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_213\ : std_logic;
signal \M_current_address_qZ0Z_8\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_218\ : std_logic;
signal \M_current_address_qZ0Z_10\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_220\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_221\ : std_logic;
signal port_data_c_6 : std_logic;
signal \this_start_data_delay.this_edge_detector.N_223\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_15\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_16\ : std_logic;
signal \M_current_address_qZ0Z_7\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_217\ : std_logic;
signal \M_current_address_qZ0Z_0\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_210\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_17\ : std_logic;
signal \this_start_address_delay.this_delay.M_pipe_qZ0Z_18\ : std_logic;
signal \M_this_start_address_delay_out_0\ : std_logic;
signal \M_state_q_ns_1_0__N_24_mux_cascade_\ : std_logic;
signal \M_state_q_ns_1_0__N_10_cascade_\ : std_logic;
signal \M_current_address_qZ0Z_1\ : std_logic;
signal \this_start_data_delay.this_edge_detector.N_211\ : std_logic;
signal \M_current_address_qZ0Z_4\ : std_logic;
signal port_data_c_4 : std_logic;
signal \this_start_data_delay.this_edge_detector.N_214\ : std_logic;
signal \M_state_qZ0Z_0\ : std_logic;
signal port_address_c_1 : std_logic;
signal \M_state_q_ns_1_0__N_24_mux\ : std_logic;
signal port_address_c_0 : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \M_this_start_data_delay_out_0\ : std_logic;
signal \M_state_q_ns_1_0__i12_mux_cascade_\ : std_logic;
signal \M_state_qZ0Z_1\ : std_logic;
signal clk_c_g : std_logic;
signal port_data_c_0 : std_logic;
signal \M_this_vram_write_data_0\ : std_logic;
signal \this_vram.mem_WE_8\ : std_logic;
signal \this_vram.mem_N_91\ : std_logic;
signal \this_vram.mem_N_88\ : std_logic;
signal \N_16_0\ : std_logic;
signal port_address_c_4 : std_logic;
signal port_address_c_7 : std_logic;
signal port_enb_c : std_logic;
signal port_address_c_2 : std_logic;
signal \M_state_q_ns_1_0__m7Z0Z_5\ : std_logic;
signal port_data_c_1 : std_logic;
signal \M_this_vram_write_data_1\ : std_logic;
signal \this_vram.mem_out_bus2_1\ : std_logic;
signal \this_vram.mem_out_bus6_1\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\ : std_logic;
signal \this_vram.mem_WE_14\ : std_logic;
signal \this_vram.mem_WE_10\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vram.mem_out_bus4_1\ : std_logic;
signal \this_vram.mem_out_bus0_1\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus7_3\ : std_logic;
signal \this_vram.mem_out_bus3_3\ : std_logic;
signal \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_102\ : std_logic;
signal \this_vram.mem_radregZ0Z_11\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \this_vram.mem_WE_12\ : std_logic;
signal \this_vram.mem_N_109\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc5\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \this_vram.mem_out_bus1_2\ : std_logic;
signal \this_vram.mem_out_bus5_2\ : std_logic;
signal \this_vram.mem_out_bus1_1\ : std_logic;
signal \this_vram.mem_out_bus5_1\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus6_0\ : std_logic;
signal \this_vram.mem_out_bus2_0\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0NZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_N_112\ : std_logic;
signal \this_vram.mem_out_bus4_0\ : std_logic;
signal \this_vram.mem_out_bus0_0\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOIZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus3_2\ : std_logic;
signal \this_vram.mem_out_bus7_2\ : std_logic;
signal \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_mem_1_1_RNIUSKZ0Z11\ : std_logic;
signal \this_vram.mem_N_95\ : std_logic;
signal \this_vram.mem_out_bus5_3\ : std_logic;
signal \this_vram.mem_out_bus1_3\ : std_logic;
signal \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus3_0\ : std_logic;
signal \this_vram.mem_out_bus7_0\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05PZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus6_3\ : std_logic;
signal \this_vram.mem_out_bus2_3\ : std_logic;
signal \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_105\ : std_logic;
signal \this_vram.mem_out_bus0_3\ : std_logic;
signal \this_vram.mem_out_bus4_3\ : std_logic;
signal \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus2_2\ : std_logic;
signal \this_vram.mem_out_bus6_2\ : std_logic;
signal \this_vram.mem_out_bus0_2\ : std_logic;
signal \this_vram.mem_out_bus4_2\ : std_logic;
signal \this_vram.mem_mem_2_1_RNI01NZ0Z11\ : std_logic;
signal \this_vram.mem_mem_0_1_RNISOIZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_radregZ0Z_12\ : std_logic;
signal \this_vram.mem_N_98\ : std_logic;
signal \this_vram.mem_out_bus1_0\ : std_logic;
signal \this_vram.mem_out_bus5_0\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSKZ0Z11\ : std_logic;
signal \this_vram.mem_radregZ0Z_13\ : std_logic;
signal \this_vram.mem_out_bus7_1\ : std_logic;
signal \this_vram.mem_out_bus3_1\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\ : std_logic;
signal \this_vram.mem_WE_6\ : std_logic;
signal \this_vram.mem_WE_4\ : std_logic;
signal \this_vram.mem_WE_2\ : std_logic;
signal \M_current_address_qZ0Z_12\ : std_logic;
signal \M_current_address_qZ0Z_11\ : std_logic;
signal \M_current_address_qZ0Z_13\ : std_logic;
signal \this_vram.mem_WE_0\ : std_logic;
signal port_data_c_2 : std_logic;
signal \M_this_vram_write_data_2\ : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_vram_write_en_0_sqmuxa\ : std_logic;
signal \M_this_vram_write_data_3\ : std_logic;
signal \this_vga_signals.g0_7\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c5\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.rgb72\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c5\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc5_1_i\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal port_rw_c : std_logic;
signal port_address_c_6 : std_logic;
signal port_address_c_5 : std_logic;
signal port_address_c_3 : std_logic;
signal \M_state_q_ns_1_0__m7Z0Z_4\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic;
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal port_address_wire : std_logic_vector(15 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal port_rw_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    port_address_wire <= port_address;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    port_rw_wire <= port_rw;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \this_vram.mem_out_bus0_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= \N__14252\&\N__11510\&\N__10451\&\N__11156\&\N__12218\&\N__18278\&\N__9338\&\N__11342\&\N__19814\&\N__20120\&\N__13949\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= \N__16013\&\N__14900\&\N__16145\&\N__15821\&\N__15386\&\N__15050\&\N__16529\&\N__15263\&\N__14687\&\N__16661\&\N__15686\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16793\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17111\&'0'&'0'&'0';
    \this_vram.mem_out_bus0_3\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_2\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_1_physical_RADDR_wire\ <= \N__14246\&\N__11504\&\N__10445\&\N__11150\&\N__12212\&\N__18272\&\N__9332\&\N__11336\&\N__19808\&\N__20114\&\N__13943\;
    \this_vram.mem_mem_0_1_physical_WADDR_wire\ <= \N__16007\&\N__14894\&\N__16139\&\N__15815\&\N__15380\&\N__15044\&\N__16523\&\N__15257\&\N__14681\&\N__16655\&\N__15680\;
    \this_vram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20228\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18996\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_1\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_0\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_0_physical_RADDR_wire\ <= \N__14240\&\N__11498\&\N__10439\&\N__11144\&\N__12206\&\N__18266\&\N__9326\&\N__11330\&\N__19802\&\N__20108\&\N__13937\;
    \this_vram.mem_mem_1_0_physical_WADDR_wire\ <= \N__16001\&\N__14888\&\N__16133\&\N__15809\&\N__15374\&\N__15038\&\N__16517\&\N__15251\&\N__14675\&\N__16649\&\N__15674\;
    \this_vram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16789\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17107\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_3\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_2\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_1_physical_RADDR_wire\ <= \N__14234\&\N__11492\&\N__10433\&\N__11138\&\N__12200\&\N__18260\&\N__9320\&\N__11324\&\N__19796\&\N__20102\&\N__13931\;
    \this_vram.mem_mem_1_1_physical_WADDR_wire\ <= \N__15995\&\N__14882\&\N__16127\&\N__15803\&\N__15368\&\N__15032\&\N__16511\&\N__15245\&\N__14669\&\N__16643\&\N__15668\;
    \this_vram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20224\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19001\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_1\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_0\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_0_physical_RADDR_wire\ <= \N__14228\&\N__11486\&\N__10427\&\N__11132\&\N__12194\&\N__18254\&\N__9314\&\N__11318\&\N__19790\&\N__20096\&\N__13925\;
    \this_vram.mem_mem_2_0_physical_WADDR_wire\ <= \N__15989\&\N__14876\&\N__16121\&\N__15797\&\N__15362\&\N__15026\&\N__16505\&\N__15239\&\N__14663\&\N__16637\&\N__15662\;
    \this_vram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16782\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17100\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_3\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_2\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_1_physical_RADDR_wire\ <= \N__14222\&\N__11480\&\N__10421\&\N__11126\&\N__12188\&\N__18248\&\N__9308\&\N__11312\&\N__19784\&\N__20090\&\N__13919\;
    \this_vram.mem_mem_2_1_physical_WADDR_wire\ <= \N__15983\&\N__14870\&\N__16115\&\N__15791\&\N__15356\&\N__15020\&\N__16499\&\N__15233\&\N__14657\&\N__16631\&\N__15656\;
    \this_vram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20217\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18997\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_1\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_0\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_0_physical_RADDR_wire\ <= \N__14216\&\N__11474\&\N__10415\&\N__11120\&\N__12182\&\N__18242\&\N__9302\&\N__11306\&\N__19778\&\N__20084\&\N__13913\;
    \this_vram.mem_mem_3_0_physical_WADDR_wire\ <= \N__15977\&\N__14864\&\N__16109\&\N__15785\&\N__15350\&\N__15014\&\N__16493\&\N__15227\&\N__14651\&\N__16625\&\N__15650\;
    \this_vram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16772\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17091\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_3\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_2\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_1_physical_RADDR_wire\ <= \N__14210\&\N__11468\&\N__10409\&\N__11114\&\N__12176\&\N__18236\&\N__9296\&\N__11300\&\N__19772\&\N__20078\&\N__13907\;
    \this_vram.mem_mem_3_1_physical_WADDR_wire\ <= \N__15971\&\N__14858\&\N__16103\&\N__15779\&\N__15344\&\N__15008\&\N__16487\&\N__15221\&\N__14645\&\N__16619\&\N__15644\;
    \this_vram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20208\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18989\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_1\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_0\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_0_physical_RADDR_wire\ <= \N__14204\&\N__11462\&\N__10403\&\N__11108\&\N__12170\&\N__18230\&\N__9290\&\N__11294\&\N__19766\&\N__20072\&\N__13901\;
    \this_vram.mem_mem_4_0_physical_WADDR_wire\ <= \N__15965\&\N__14852\&\N__16097\&\N__15773\&\N__15338\&\N__15002\&\N__16481\&\N__15215\&\N__14639\&\N__16613\&\N__15638\;
    \this_vram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16760\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17082\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_3\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_2\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_1_physical_RADDR_wire\ <= \N__14198\&\N__11456\&\N__10397\&\N__11102\&\N__12164\&\N__18224\&\N__9284\&\N__11288\&\N__19760\&\N__20066\&\N__13895\;
    \this_vram.mem_mem_4_1_physical_WADDR_wire\ <= \N__15959\&\N__14846\&\N__16091\&\N__15767\&\N__15332\&\N__14996\&\N__16475\&\N__15209\&\N__14633\&\N__16607\&\N__15632\;
    \this_vram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20199\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18977\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_1\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_0\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_0_physical_RADDR_wire\ <= \N__14192\&\N__11450\&\N__10391\&\N__11096\&\N__12158\&\N__18218\&\N__9278\&\N__11282\&\N__19754\&\N__20060\&\N__13889\;
    \this_vram.mem_mem_5_0_physical_WADDR_wire\ <= \N__15953\&\N__14840\&\N__16085\&\N__15761\&\N__15326\&\N__14990\&\N__16469\&\N__15203\&\N__14627\&\N__16601\&\N__15626\;
    \this_vram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16748\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17073\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_3\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_2\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_1_physical_RADDR_wire\ <= \N__14186\&\N__11444\&\N__10385\&\N__11090\&\N__12152\&\N__18212\&\N__9272\&\N__11276\&\N__19748\&\N__20054\&\N__13883\;
    \this_vram.mem_mem_5_1_physical_WADDR_wire\ <= \N__15947\&\N__14834\&\N__16079\&\N__15755\&\N__15320\&\N__14984\&\N__16463\&\N__15197\&\N__14621\&\N__16595\&\N__15620\;
    \this_vram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20189\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18964\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_1\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_0\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_0_physical_RADDR_wire\ <= \N__14180\&\N__11438\&\N__10379\&\N__11084\&\N__12146\&\N__18206\&\N__9266\&\N__11270\&\N__19742\&\N__20048\&\N__13877\;
    \this_vram.mem_mem_6_0_physical_WADDR_wire\ <= \N__15941\&\N__14828\&\N__16073\&\N__15749\&\N__15314\&\N__14978\&\N__16457\&\N__15191\&\N__14615\&\N__16589\&\N__15614\;
    \this_vram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16732\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17063\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_3\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_2\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_1_physical_RADDR_wire\ <= \N__14174\&\N__11432\&\N__10373\&\N__11078\&\N__12140\&\N__18200\&\N__9260\&\N__11264\&\N__19736\&\N__20042\&\N__13871\;
    \this_vram.mem_mem_6_1_physical_WADDR_wire\ <= \N__15935\&\N__14822\&\N__16067\&\N__15743\&\N__15308\&\N__14972\&\N__16451\&\N__15185\&\N__14609\&\N__16583\&\N__15608\;
    \this_vram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20168\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18960\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_1\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_0\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_0_physical_RADDR_wire\ <= \N__14168\&\N__11426\&\N__10367\&\N__11072\&\N__12134\&\N__18194\&\N__9254\&\N__11258\&\N__19730\&\N__20036\&\N__13865\;
    \this_vram.mem_mem_7_0_physical_WADDR_wire\ <= \N__15929\&\N__14816\&\N__16061\&\N__15737\&\N__15302\&\N__14966\&\N__16445\&\N__15179\&\N__14603\&\N__16577\&\N__15602\;
    \this_vram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16747\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17072\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_3\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_2\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_1_physical_RADDR_wire\ <= \N__14162\&\N__11420\&\N__10361\&\N__11066\&\N__12128\&\N__18188\&\N__9248\&\N__11252\&\N__19724\&\N__20030\&\N__13859\;
    \this_vram.mem_mem_7_1_physical_WADDR_wire\ <= \N__15923\&\N__14810\&\N__16055\&\N__15731\&\N__15296\&\N__14960\&\N__16439\&\N__15173\&\N__14597\&\N__16571\&\N__15596\;
    \this_vram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__20190\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18976\&'0'&'0'&'0';

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17302\,
            RE => \N__18695\,
            WCLKE => \N__17984\,
            WCLK => \N__17303\,
            WE => \N__18610\
        );

    \this_vram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17304\,
            RE => \N__18691\,
            WCLKE => \N__17980\,
            WCLK => \N__17305\,
            WE => \N__18688\
        );

    \this_vram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17306\,
            RE => \N__18690\,
            WCLKE => \N__17771\,
            WCLK => \N__17307\,
            WE => \N__18687\
        );

    \this_vram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17308\,
            RE => \N__18666\,
            WCLKE => \N__17767\,
            WCLK => \N__17309\,
            WE => \N__18677\
        );

    \this_vram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17311\,
            RE => \N__18665\,
            WCLKE => \N__17951\,
            WCLK => \N__17310\,
            WE => \N__18609\
        );

    \this_vram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17313\,
            RE => \N__18634\,
            WCLKE => \N__17947\,
            WCLK => \N__17314\,
            WE => \N__18654\
        );

    \this_vram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17321\,
            RE => \N__18633\,
            WCLKE => \N__17036\,
            WCLK => \N__17322\,
            WE => \N__18563\
        );

    \this_vram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17334\,
            RE => \N__18595\,
            WCLKE => \N__17032\,
            WCLK => \N__17335\,
            WE => \N__18624\
        );

    \this_vram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17344\,
            RE => \N__18594\,
            WCLKE => \N__19403\,
            WCLK => \N__17345\,
            WE => \N__18575\
        );

    \this_vram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17355\,
            RE => \N__18515\,
            WCLKE => \N__19399\,
            WCLK => \N__17356\,
            WE => \N__18562\
        );

    \this_vram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17366\,
            RE => \N__18514\,
            WCLKE => \N__19376\,
            WCLK => \N__17367\,
            WE => \N__18495\
        );

    \this_vram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17369\,
            RE => \N__18519\,
            WCLKE => \N__19372\,
            WCLK => \N__17370\,
            WE => \N__18521\
        );

    \this_vram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17371\,
            RE => \N__18520\,
            WCLKE => \N__19348\,
            WCLK => \N__17372\,
            WE => \N__18522\
        );

    \this_vram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17373\,
            RE => \N__18576\,
            WCLKE => \N__19349\,
            WCLK => \N__17374\,
            WE => \N__18581\
        );

    \this_vram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17375\,
            RE => \N__18577\,
            WCLKE => \N__19057\,
            WCLK => \N__17376\,
            WE => \N__18582\
        );

    \this_vram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__17377\,
            RE => \N__18623\,
            WCLKE => \N__19058\,
            WCLK => \N__17378\,
            WE => \N__18622\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__20688\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20690\,
            DIN => \N__20689\,
            DOUT => \N__20688\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20690\,
            PADOUT => \N__20689\,
            PADIN => \N__20688\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20679\,
            DIN => \N__20678\,
            DOUT => \N__20677\,
            PACKAGEPIN => debug_wire
        );

    \debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20679\,
            PADOUT => \N__20678\,
            PADIN => \N__20677\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14453\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20670\,
            DIN => \N__20669\,
            DOUT => \N__20668\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20670\,
            PADOUT => \N__20669\,
            PADIN => \N__20668\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8300\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20661\,
            DIN => \N__20660\,
            DOUT => \N__20659\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20661\,
            PADOUT => \N__20660\,
            PADIN => \N__20659\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7298\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20652\,
            DIN => \N__20651\,
            DOUT => \N__20650\,
            PACKAGEPIN => port_address_wire(0)
        );

    \port_address_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20652\,
            PADOUT => \N__20651\,
            PADIN => \N__20650\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20643\,
            DIN => \N__20642\,
            DOUT => \N__20641\,
            PACKAGEPIN => port_address_wire(1)
        );

    \port_address_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20643\,
            PADOUT => \N__20642\,
            PADIN => \N__20641\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20634\,
            DIN => \N__20633\,
            DOUT => \N__20632\,
            PACKAGEPIN => port_address_wire(2)
        );

    \port_address_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20634\,
            PADOUT => \N__20633\,
            PADIN => \N__20632\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20625\,
            DIN => \N__20624\,
            DOUT => \N__20623\,
            PACKAGEPIN => port_address_wire(3)
        );

    \port_address_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20625\,
            PADOUT => \N__20624\,
            PADIN => \N__20623\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20616\,
            DIN => \N__20615\,
            DOUT => \N__20614\,
            PACKAGEPIN => port_address_wire(4)
        );

    \port_address_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20616\,
            PADOUT => \N__20615\,
            PADIN => \N__20614\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20607\,
            DIN => \N__20606\,
            DOUT => \N__20605\,
            PACKAGEPIN => port_address_wire(5)
        );

    \port_address_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20607\,
            PADOUT => \N__20606\,
            PADIN => \N__20605\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20598\,
            DIN => \N__20597\,
            DOUT => \N__20596\,
            PACKAGEPIN => port_address_wire(6)
        );

    \port_address_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20598\,
            PADOUT => \N__20597\,
            PADIN => \N__20596\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20589\,
            DIN => \N__20588\,
            DOUT => \N__20587\,
            PACKAGEPIN => port_address_wire(7)
        );

    \port_address_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20589\,
            PADOUT => \N__20588\,
            PADIN => \N__20587\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20580\,
            DIN => \N__20579\,
            DOUT => \N__20578\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20580\,
            PADOUT => \N__20579\,
            PADIN => \N__20578\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20571\,
            DIN => \N__20570\,
            DOUT => \N__20569\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20571\,
            PADOUT => \N__20570\,
            PADIN => \N__20569\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20562\,
            DIN => \N__20561\,
            DOUT => \N__20560\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20562\,
            PADOUT => \N__20561\,
            PADIN => \N__20560\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20553\,
            DIN => \N__20552\,
            DOUT => \N__20551\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20553\,
            PADOUT => \N__20552\,
            PADIN => \N__20551\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20544\,
            DIN => \N__20543\,
            DOUT => \N__20542\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20544\,
            PADOUT => \N__20543\,
            PADIN => \N__20542\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20535\,
            DIN => \N__20534\,
            DOUT => \N__20533\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20535\,
            PADOUT => \N__20534\,
            PADIN => \N__20533\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20526\,
            DIN => \N__20525\,
            DOUT => \N__20524\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20526\,
            PADOUT => \N__20525\,
            PADIN => \N__20524\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20517\,
            DIN => \N__20516\,
            DOUT => \N__20515\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20517\,
            PADOUT => \N__20516\,
            PADIN => \N__20515\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20508\,
            DIN => \N__20507\,
            DOUT => \N__20506\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20508\,
            PADOUT => \N__20507\,
            PADIN => \N__20506\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7217\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20499\,
            DIN => \N__20498\,
            DOUT => \N__20497\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20499\,
            PADOUT => \N__20498\,
            PADIN => \N__20497\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__18689\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20490\,
            DIN => \N__20489\,
            DOUT => \N__20488\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20490\,
            PADOUT => \N__20489\,
            PADIN => \N__20488\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20481\,
            DIN => \N__20480\,
            DOUT => \N__20479\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20481\,
            PADOUT => \N__20480\,
            PADIN => \N__20479\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7802\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20472\,
            DIN => \N__20471\,
            DOUT => \N__20470\,
            PACKAGEPIN => port_rw_wire
        );

    \port_rw_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20472\,
            PADOUT => \N__20471\,
            PADIN => \N__20470\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20463\,
            DIN => \N__20462\,
            DOUT => \N__20461\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20463\,
            PADOUT => \N__20462\,
            PADIN => \N__20461\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__9050\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20454\,
            DIN => \N__20453\,
            DOUT => \N__20452\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20454\,
            PADOUT => \N__20453\,
            PADIN => \N__20452\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__9040\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20445\,
            DIN => \N__20444\,
            DOUT => \N__20443\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20445\,
            PADOUT => \N__20444\,
            PADIN => \N__20443\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12088\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20436\,
            DIN => \N__20435\,
            DOUT => \N__20434\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20436\,
            PADOUT => \N__20435\,
            PADIN => \N__20434\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12098\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20427\,
            DIN => \N__20426\,
            DOUT => \N__20425\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20427\,
            PADOUT => \N__20426\,
            PADIN => \N__20425\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8707\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20418\,
            DIN => \N__20417\,
            DOUT => \N__20416\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20418\,
            PADOUT => \N__20417\,
            PADIN => \N__20416\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8714\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20409\,
            DIN => \N__20408\,
            DOUT => \N__20407\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20409\,
            PADOUT => \N__20408\,
            PADIN => \N__20407\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20400\,
            DIN => \N__20399\,
            DOUT => \N__20398\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20400\,
            PADOUT => \N__20399\,
            PADIN => \N__20398\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7211\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20391\,
            DIN => \N__20390\,
            DOUT => \N__20389\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20391\,
            PADOUT => \N__20390\,
            PADIN => \N__20389\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__9515\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__4904\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20365\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__20368\,
            I => \N__20362\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__20365\,
            I => \N__20359\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20356\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__20359\,
            I => \N__20353\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20350\
        );

    \I__4898\ : Span4Mux_v
    port map (
            O => \N__20353\,
            I => \N__20344\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__20350\,
            I => \N__20344\
        );

    \I__4896\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20341\
        );

    \I__4895\ : Sp12to4
    port map (
            O => \N__20344\,
            I => \N__20336\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__20341\,
            I => \N__20336\
        );

    \I__4893\ : Span12Mux_h
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__4892\ : Odrv12
    port map (
            O => \N__20333\,
            I => port_data_c_3
        );

    \I__4891\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20321\
        );

    \I__4890\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20321\
        );

    \I__4889\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20314\
        );

    \I__4888\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20310\
        );

    \I__4887\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20307\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__20321\,
            I => \N__20304\
        );

    \I__4885\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20301\
        );

    \I__4884\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20298\
        );

    \I__4883\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20295\
        );

    \I__4882\ : InMux
    port map (
            O => \N__20317\,
            I => \N__20292\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__20314\,
            I => \N__20289\
        );

    \I__4880\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20286\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__20310\,
            I => \N__20281\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__20307\,
            I => \N__20278\
        );

    \I__4877\ : Span4Mux_v
    port map (
            O => \N__20304\,
            I => \N__20273\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__20301\,
            I => \N__20273\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20262\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20262\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20262\
        );

    \I__4872\ : Span4Mux_v
    port map (
            O => \N__20289\,
            I => \N__20262\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__20286\,
            I => \N__20262\
        );

    \I__4870\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20259\
        );

    \I__4869\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20256\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__20281\,
            I => \N__20253\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__20278\,
            I => \N__20250\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__20273\,
            I => \N__20245\
        );

    \I__4865\ : Span4Mux_v
    port map (
            O => \N__20262\,
            I => \N__20245\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__20259\,
            I => \N__20242\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__20256\,
            I => \N__20239\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__20253\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__20250\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__20245\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4859\ : Odrv12
    port map (
            O => \N__20242\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__20239\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4857\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20221\
        );

    \I__4855\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20218\
        );

    \I__4854\ : Span4Mux_v
    port map (
            O => \N__20221\,
            I => \N__20212\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__20218\,
            I => \N__20212\
        );

    \I__4852\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20209\
        );

    \I__4851\ : Span4Mux_v
    port map (
            O => \N__20212\,
            I => \N__20203\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__20209\,
            I => \N__20203\
        );

    \I__4849\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20200\
        );

    \I__4848\ : Span4Mux_v
    port map (
            O => \N__20203\,
            I => \N__20194\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__20200\,
            I => \N__20194\
        );

    \I__4846\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20191\
        );

    \I__4845\ : Span4Mux_v
    port map (
            O => \N__20194\,
            I => \N__20184\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__20191\,
            I => \N__20184\
        );

    \I__4843\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20181\
        );

    \I__4842\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20178\
        );

    \I__4841\ : Span4Mux_v
    port map (
            O => \N__20184\,
            I => \N__20175\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20172\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20169\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__20175\,
            I => \N__20163\
        );

    \I__4837\ : Span4Mux_s2_v
    port map (
            O => \N__20172\,
            I => \N__20163\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__20169\,
            I => \N__20160\
        );

    \I__4835\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20157\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__20163\,
            I => \M_this_vram_write_data_3\
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__20160\,
            I => \M_this_vram_write_data_3\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__20157\,
            I => \M_this_vram_write_data_3\
        );

    \I__4831\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__4829\ : Span12Mux_s10_h
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__4828\ : Span12Mux_v
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__4827\ : Odrv12
    port map (
            O => \N__20138\,
            I => \this_vga_signals.g0_7\
        );

    \I__4826\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__4824\ : Span12Mux_h
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__4823\ : Span12Mux_v
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__20123\,
            I => \this_vga_signals.mult1_un89_sum_c5\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__4820\ : CascadeBuf
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__4818\ : CascadeBuf
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__4816\ : CascadeBuf
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__4815\ : CascadeMux
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__4814\ : CascadeBuf
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__4812\ : CascadeBuf
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__4811\ : CascadeMux
    port map (
            O => \N__20090\,
            I => \N__20087\
        );

    \I__4810\ : CascadeBuf
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__4809\ : CascadeMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__4808\ : CascadeBuf
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__4807\ : CascadeMux
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__4806\ : CascadeBuf
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__4804\ : CascadeBuf
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__4802\ : CascadeBuf
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__4800\ : CascadeBuf
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__4798\ : CascadeBuf
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__4796\ : CascadeBuf
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__4794\ : CascadeBuf
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__4792\ : CascadeBuf
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__4790\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__20024\,
            I => \M_this_vga_signals_address_1\
        );

    \I__4788\ : InMux
    port map (
            O => \N__20021\,
            I => \N__20016\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__20020\,
            I => \N__20013\
        );

    \I__4786\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20009\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20016\,
            I => \N__20003\
        );

    \I__4784\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20000\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__20012\,
            I => \N__19996\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__20009\,
            I => \N__19990\
        );

    \I__4781\ : InMux
    port map (
            O => \N__20008\,
            I => \N__19987\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20007\,
            I => \N__19982\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20006\,
            I => \N__19979\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__20003\,
            I => \N__19976\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20000\,
            I => \N__19973\
        );

    \I__4776\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19970\
        );

    \I__4775\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19967\
        );

    \I__4774\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19964\
        );

    \I__4773\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19961\
        );

    \I__4772\ : InMux
    port map (
            O => \N__19993\,
            I => \N__19958\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__19990\,
            I => \N__19953\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__19987\,
            I => \N__19953\
        );

    \I__4769\ : InMux
    port map (
            O => \N__19986\,
            I => \N__19950\
        );

    \I__4768\ : CascadeMux
    port map (
            O => \N__19985\,
            I => \N__19947\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19943\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__19979\,
            I => \N__19940\
        );

    \I__4765\ : Sp12to4
    port map (
            O => \N__19976\,
            I => \N__19937\
        );

    \I__4764\ : Span4Mux_h
    port map (
            O => \N__19973\,
            I => \N__19934\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19931\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__19967\,
            I => \N__19928\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__19964\,
            I => \N__19917\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__19961\,
            I => \N__19917\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19917\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__19953\,
            I => \N__19917\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__19950\,
            I => \N__19917\
        );

    \I__4756\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19914\
        );

    \I__4755\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19911\
        );

    \I__4754\ : Span12Mux_v
    port map (
            O => \N__19943\,
            I => \N__19908\
        );

    \I__4753\ : Span4Mux_v
    port map (
            O => \N__19940\,
            I => \N__19905\
        );

    \I__4752\ : Span12Mux_h
    port map (
            O => \N__19937\,
            I => \N__19902\
        );

    \I__4751\ : Sp12to4
    port map (
            O => \N__19934\,
            I => \N__19899\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__19931\,
            I => \N__19890\
        );

    \I__4749\ : Span4Mux_h
    port map (
            O => \N__19928\,
            I => \N__19890\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__19917\,
            I => \N__19890\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__19914\,
            I => \N__19890\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19887\
        );

    \I__4745\ : Span12Mux_h
    port map (
            O => \N__19908\,
            I => \N__19884\
        );

    \I__4744\ : Sp12to4
    port map (
            O => \N__19905\,
            I => \N__19877\
        );

    \I__4743\ : Span12Mux_v
    port map (
            O => \N__19902\,
            I => \N__19877\
        );

    \I__4742\ : Span12Mux_v
    port map (
            O => \N__19899\,
            I => \N__19877\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__19890\,
            I => \N__19874\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__19887\,
            I => \this_vga_signals.rgb72\
        );

    \I__4739\ : Odrv12
    port map (
            O => \N__19884\,
            I => \this_vga_signals.rgb72\
        );

    \I__4738\ : Odrv12
    port map (
            O => \N__19877\,
            I => \this_vga_signals.rgb72\
        );

    \I__4737\ : Odrv4
    port map (
            O => \N__19874\,
            I => \this_vga_signals.rgb72\
        );

    \I__4736\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19861\
        );

    \I__4735\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19858\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__19861\,
            I => \N__19855\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__19858\,
            I => \N__19852\
        );

    \I__4732\ : Span12Mux_s7_v
    port map (
            O => \N__19855\,
            I => \N__19849\
        );

    \I__4731\ : Span12Mux_h
    port map (
            O => \N__19852\,
            I => \N__19846\
        );

    \I__4730\ : Span12Mux_h
    port map (
            O => \N__19849\,
            I => \N__19843\
        );

    \I__4729\ : Span12Mux_v
    port map (
            O => \N__19846\,
            I => \N__19840\
        );

    \I__4728\ : Odrv12
    port map (
            O => \N__19843\,
            I => \this_vga_signals.mult1_un82_sum_c5\
        );

    \I__4727\ : Odrv12
    port map (
            O => \N__19840\,
            I => \this_vga_signals.mult1_un82_sum_c5\
        );

    \I__4726\ : InMux
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__4724\ : Span12Mux_s10_v
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__4723\ : Span12Mux_h
    port map (
            O => \N__19826\,
            I => \N__19822\
        );

    \I__4722\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19819\
        );

    \I__4721\ : Odrv12
    port map (
            O => \N__19822\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_i\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__19819\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_i\
        );

    \I__4719\ : CascadeMux
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__4718\ : CascadeBuf
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__4717\ : CascadeMux
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__4716\ : CascadeBuf
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__4714\ : CascadeBuf
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__4712\ : CascadeBuf
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__4711\ : CascadeMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__4710\ : CascadeBuf
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__4709\ : CascadeMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__4708\ : CascadeBuf
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__4706\ : CascadeBuf
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__4704\ : CascadeBuf
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__4702\ : CascadeBuf
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__4700\ : CascadeBuf
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__4698\ : CascadeBuf
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4696\ : CascadeBuf
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__4694\ : CascadeBuf
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__4692\ : CascadeBuf
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__4690\ : CascadeBuf
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__4688\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__19718\,
            I => \M_this_vga_signals_address_2\
        );

    \I__4686\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__4684\ : Span12Mux_s10_h
    port map (
            O => \N__19709\,
            I => \N__19706\
        );

    \I__4683\ : Span12Mux_h
    port map (
            O => \N__19706\,
            I => \N__19702\
        );

    \I__4682\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19699\
        );

    \I__4681\ : Odrv12
    port map (
            O => \N__19702\,
            I => port_rw_c
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__19699\,
            I => port_rw_c
        );

    \I__4679\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__4677\ : Span12Mux_v
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__4676\ : Odrv12
    port map (
            O => \N__19685\,
            I => port_address_c_6
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__4674\ : InMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__19676\,
            I => port_address_c_5
        );

    \I__4672\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__4670\ : Span12Mux_v
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__4669\ : Odrv12
    port map (
            O => \N__19664\,
            I => port_address_c_3
        );

    \I__4668\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__4665\ : Span4Mux_h
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4664\ : Span4Mux_h
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__19646\,
            I => \M_state_q_ns_1_0__m7Z0Z_4\
        );

    \I__4662\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__19640\,
            I => \this_vram.mem_mem_2_1_RNI01NZ0Z11\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \this_vram.mem_mem_0_1_RNISOIZ0Z11_cascade_\
        );

    \I__4659\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19629\
        );

    \I__4658\ : InMux
    port map (
            O => \N__19633\,
            I => \N__19626\
        );

    \I__4657\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19623\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__19629\,
            I => \N__19614\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__19626\,
            I => \N__19614\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19611\
        );

    \I__4653\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19607\
        );

    \I__4652\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19604\
        );

    \I__4651\ : InMux
    port map (
            O => \N__19620\,
            I => \N__19601\
        );

    \I__4650\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19598\
        );

    \I__4649\ : Span4Mux_v
    port map (
            O => \N__19614\,
            I => \N__19593\
        );

    \I__4648\ : Span4Mux_v
    port map (
            O => \N__19611\,
            I => \N__19593\
        );

    \I__4647\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19590\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__19607\,
            I => \N__19585\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__19604\,
            I => \N__19585\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__19601\,
            I => \N__19576\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19576\
        );

    \I__4642\ : Sp12to4
    port map (
            O => \N__19593\,
            I => \N__19576\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__19590\,
            I => \N__19576\
        );

    \I__4640\ : Sp12to4
    port map (
            O => \N__19585\,
            I => \N__19573\
        );

    \I__4639\ : Span12Mux_h
    port map (
            O => \N__19576\,
            I => \N__19570\
        );

    \I__4638\ : Span12Mux_v
    port map (
            O => \N__19573\,
            I => \N__19567\
        );

    \I__4637\ : Odrv12
    port map (
            O => \N__19570\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__4636\ : Odrv12
    port map (
            O => \N__19567\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__4635\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__19559\,
            I => \this_vram.mem_N_98\
        );

    \I__4633\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__4631\ : Span12Mux_h
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__4630\ : Span12Mux_v
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__4629\ : Odrv12
    port map (
            O => \N__19544\,
            I => \this_vram.mem_out_bus1_0\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__19532\,
            I => \this_vram.mem_out_bus5_0\
        );

    \I__4624\ : InMux
    port map (
            O => \N__19529\,
            I => \N__19526\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__19526\,
            I => \this_vram.mem_mem_1_0_RNISSKZ0Z11\
        );

    \I__4622\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19504\
        );

    \I__4621\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19504\
        );

    \I__4620\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19504\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19504\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19497\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19497\
        );

    \I__4616\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19497\
        );

    \I__4615\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19494\
        );

    \I__4614\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19491\
        );

    \I__4613\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19486\
        );

    \I__4612\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19486\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__19504\,
            I => \N__19475\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19475\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__19494\,
            I => \N__19475\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19475\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__19486\,
            I => \N__19475\
        );

    \I__4606\ : Span4Mux_v
    port map (
            O => \N__19475\,
            I => \N__19467\
        );

    \I__4605\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19464\
        );

    \I__4604\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19457\
        );

    \I__4603\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19457\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19457\
        );

    \I__4601\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19454\
        );

    \I__4600\ : Sp12to4
    port map (
            O => \N__19467\,
            I => \N__19445\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__19464\,
            I => \N__19445\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__19457\,
            I => \N__19445\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__19454\,
            I => \N__19445\
        );

    \I__4596\ : Span12Mux_h
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__4595\ : Odrv12
    port map (
            O => \N__19442\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__4594\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19436\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__19436\,
            I => \N__19433\
        );

    \I__4592\ : Span4Mux_v
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__4591\ : Span4Mux_v
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__19427\,
            I => \this_vram.mem_out_bus7_1\
        );

    \I__4589\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__19421\,
            I => \N__19418\
        );

    \I__4587\ : Span4Mux_v
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__19415\,
            I => \this_vram.mem_out_bus3_1\
        );

    \I__4585\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__19406\,
            I => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\
        );

    \I__4582\ : CEMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__19400\,
            I => \N__19396\
        );

    \I__4580\ : CEMux
    port map (
            O => \N__19399\,
            I => \N__19393\
        );

    \I__4579\ : Span4Mux_v
    port map (
            O => \N__19396\,
            I => \N__19390\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__19393\,
            I => \N__19387\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__19390\,
            I => \N__19384\
        );

    \I__4576\ : Span4Mux_h
    port map (
            O => \N__19387\,
            I => \N__19381\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__19384\,
            I => \this_vram.mem_WE_6\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__19381\,
            I => \this_vram.mem_WE_6\
        );

    \I__4573\ : CEMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__19373\,
            I => \N__19369\
        );

    \I__4571\ : CEMux
    port map (
            O => \N__19372\,
            I => \N__19366\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19360\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__19363\,
            I => \N__19357\
        );

    \I__4567\ : Span4Mux_h
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__19357\,
            I => \this_vram.mem_WE_4\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__19354\,
            I => \this_vram.mem_WE_4\
        );

    \I__4564\ : CEMux
    port map (
            O => \N__19349\,
            I => \N__19345\
        );

    \I__4563\ : CEMux
    port map (
            O => \N__19348\,
            I => \N__19342\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__19345\,
            I => \N__19339\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__19342\,
            I => \N__19336\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__19339\,
            I => \N__19333\
        );

    \I__4559\ : Span4Mux_h
    port map (
            O => \N__19336\,
            I => \N__19330\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__19333\,
            I => \this_vram.mem_WE_2\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__19330\,
            I => \this_vram.mem_WE_2\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19319\
        );

    \I__4555\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19319\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19312\
        );

    \I__4553\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19309\
        );

    \I__4552\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19304\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19301\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19298\
        );

    \I__4549\ : Span4Mux_h
    port map (
            O => \N__19312\,
            I => \N__19293\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__19309\,
            I => \N__19293\
        );

    \I__4547\ : InMux
    port map (
            O => \N__19308\,
            I => \N__19290\
        );

    \I__4546\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19287\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__19304\,
            I => \N__19279\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19279\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__19298\,
            I => \N__19279\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__19293\,
            I => \N__19274\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__19290\,
            I => \N__19274\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__19287\,
            I => \N__19270\
        );

    \I__4539\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19267\
        );

    \I__4538\ : Span12Mux_v
    port map (
            O => \N__19279\,
            I => \N__19264\
        );

    \I__4537\ : Span4Mux_v
    port map (
            O => \N__19274\,
            I => \N__19261\
        );

    \I__4536\ : InMux
    port map (
            O => \N__19273\,
            I => \N__19258\
        );

    \I__4535\ : Span12Mux_h
    port map (
            O => \N__19270\,
            I => \N__19253\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__19267\,
            I => \N__19253\
        );

    \I__4533\ : Odrv12
    port map (
            O => \N__19264\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__19261\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__19258\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4530\ : Odrv12
    port map (
            O => \N__19253\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4529\ : CascadeMux
    port map (
            O => \N__19244\,
            I => \N__19240\
        );

    \I__4528\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19234\
        );

    \I__4527\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19229\
        );

    \I__4526\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19229\
        );

    \I__4525\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19226\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19237\,
            I => \N__19223\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__19234\,
            I => \N__19218\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__19229\,
            I => \N__19211\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19211\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19223\,
            I => \N__19211\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19208\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19205\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__19218\,
            I => \N__19200\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__19211\,
            I => \N__19197\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__19208\,
            I => \N__19192\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19205\,
            I => \N__19192\
        );

    \I__4513\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19189\
        );

    \I__4512\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19186\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__19200\,
            I => \N__19182\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__19197\,
            I => \N__19177\
        );

    \I__4509\ : Span4Mux_v
    port map (
            O => \N__19192\,
            I => \N__19177\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19174\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__19186\,
            I => \N__19171\
        );

    \I__4506\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19168\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__19182\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__19177\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4503\ : Odrv12
    port map (
            O => \N__19174\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__19171\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19168\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__19157\,
            I => \N__19152\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__19156\,
            I => \N__19146\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__19155\,
            I => \N__19143\
        );

    \I__4497\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19139\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__19151\,
            I => \N__19136\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__19150\,
            I => \N__19133\
        );

    \I__4494\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19128\
        );

    \I__4493\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19128\
        );

    \I__4492\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19125\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__19142\,
            I => \N__19122\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__19139\,
            I => \N__19119\
        );

    \I__4489\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19116\
        );

    \I__4488\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19113\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__19128\,
            I => \N__19107\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__19125\,
            I => \N__19107\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19104\
        );

    \I__4484\ : Span4Mux_v
    port map (
            O => \N__19119\,
            I => \N__19097\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__19116\,
            I => \N__19097\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__19113\,
            I => \N__19097\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__19112\,
            I => \N__19094\
        );

    \I__4480\ : Sp12to4
    port map (
            O => \N__19107\,
            I => \N__19089\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19104\,
            I => \N__19089\
        );

    \I__4478\ : Span4Mux_v
    port map (
            O => \N__19097\,
            I => \N__19086\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19083\
        );

    \I__4476\ : Span12Mux_v
    port map (
            O => \N__19089\,
            I => \N__19078\
        );

    \I__4475\ : Sp12to4
    port map (
            O => \N__19086\,
            I => \N__19073\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__19083\,
            I => \N__19073\
        );

    \I__4473\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19070\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19067\
        );

    \I__4471\ : Odrv12
    port map (
            O => \N__19078\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__4470\ : Odrv12
    port map (
            O => \N__19073\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__19070\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19067\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__4467\ : CEMux
    port map (
            O => \N__19058\,
            I => \N__19054\
        );

    \I__4466\ : CEMux
    port map (
            O => \N__19057\,
            I => \N__19051\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19054\,
            I => \N__19046\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__19051\,
            I => \N__19046\
        );

    \I__4463\ : Span4Mux_v
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__4462\ : Span4Mux_h
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__19040\,
            I => \this_vram.mem_WE_0\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__19037\,
            I => \N__19032\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__19036\,
            I => \N__19029\
        );

    \I__4458\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19026\
        );

    \I__4457\ : InMux
    port map (
            O => \N__19032\,
            I => \N__19021\
        );

    \I__4456\ : InMux
    port map (
            O => \N__19029\,
            I => \N__19021\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__19026\,
            I => \N__19018\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__19021\,
            I => \N__19015\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__19018\,
            I => \N__19012\
        );

    \I__4452\ : Span12Mux_h
    port map (
            O => \N__19015\,
            I => \N__19009\
        );

    \I__4451\ : IoSpan4Mux
    port map (
            O => \N__19012\,
            I => \N__19006\
        );

    \I__4450\ : Odrv12
    port map (
            O => \N__19009\,
            I => port_data_c_2
        );

    \I__4449\ : Odrv4
    port map (
            O => \N__19006\,
            I => port_data_c_2
        );

    \I__4448\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__18998\,
            I => \N__18993\
        );

    \I__4446\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18990\
        );

    \I__4445\ : InMux
    port map (
            O => \N__18996\,
            I => \N__18986\
        );

    \I__4444\ : Span4Mux_v
    port map (
            O => \N__18993\,
            I => \N__18981\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__18990\,
            I => \N__18981\
        );

    \I__4442\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18978\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__18986\,
            I => \N__18973\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__18981\,
            I => \N__18968\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__18978\,
            I => \N__18968\
        );

    \I__4438\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18965\
        );

    \I__4437\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18961\
        );

    \I__4436\ : Span12Mux_v
    port map (
            O => \N__18973\,
            I => \N__18957\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__18968\,
            I => \N__18952\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__18965\,
            I => \N__18952\
        );

    \I__4433\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18949\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18946\
        );

    \I__4431\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18943\
        );

    \I__4430\ : Span12Mux_v
    port map (
            O => \N__18957\,
            I => \N__18940\
        );

    \I__4429\ : Span4Mux_v
    port map (
            O => \N__18952\,
            I => \N__18935\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__18949\,
            I => \N__18935\
        );

    \I__4427\ : Span4Mux_s3_v
    port map (
            O => \N__18946\,
            I => \N__18930\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__18943\,
            I => \N__18930\
        );

    \I__4425\ : Odrv12
    port map (
            O => \N__18940\,
            I => \M_this_vram_write_data_2\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__18935\,
            I => \M_this_vram_write_data_2\
        );

    \I__4423\ : Odrv4
    port map (
            O => \N__18930\,
            I => \M_this_vram_write_data_2\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__18923\,
            I => \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_\
        );

    \I__4421\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__18917\,
            I => \this_vram.mem_mem_1_1_RNIUSKZ0Z11\
        );

    \I__4419\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__18905\,
            I => \this_vram.mem_N_95\
        );

    \I__4415\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__4413\ : Span4Mux_v
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4412\ : Odrv4
    port map (
            O => \N__18893\,
            I => \this_vram.mem_out_bus5_3\
        );

    \I__4411\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__4409\ : Span4Mux_v
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__4408\ : Span4Mux_v
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__18878\,
            I => \this_vram.mem_out_bus1_3\
        );

    \I__4406\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__18872\,
            I => \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0\
        );

    \I__4404\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__18866\,
            I => \N__18863\
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__18863\,
            I => \this_vram.mem_out_bus3_0\
        );

    \I__4401\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__4399\ : Sp12to4
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__4398\ : Span12Mux_v
    port map (
            O => \N__18851\,
            I => \N__18848\
        );

    \I__4397\ : Odrv12
    port map (
            O => \N__18848\,
            I => \this_vram.mem_out_bus7_0\
        );

    \I__4396\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__18842\,
            I => \this_vram.mem_mem_3_0_RNI05PZ0Z11\
        );

    \I__4394\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__4392\ : Sp12to4
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__4391\ : Span12Mux_v
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__4390\ : Odrv12
    port map (
            O => \N__18827\,
            I => \this_vram.mem_out_bus6_3\
        );

    \I__4389\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__4387\ : Sp12to4
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__4386\ : Span12Mux_v
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__4385\ : Odrv12
    port map (
            O => \N__18812\,
            I => \this_vram.mem_out_bus2_3\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__18809\,
            I => \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_\
        );

    \I__4383\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__18803\,
            I => \this_vram.mem_N_105\
        );

    \I__4381\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__4379\ : Sp12to4
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__4378\ : Span12Mux_v
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__4377\ : Odrv12
    port map (
            O => \N__18788\,
            I => \this_vram.mem_out_bus0_3\
        );

    \I__4376\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__18779\,
            I => \this_vram.mem_out_bus4_3\
        );

    \I__4373\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__18773\,
            I => \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\
        );

    \I__4371\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__4369\ : Span4Mux_h
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__4368\ : Span4Mux_v
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__4367\ : Odrv4
    port map (
            O => \N__18758\,
            I => \this_vram.mem_out_bus2_2\
        );

    \I__4366\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__4363\ : Span4Mux_v
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__18743\,
            I => \this_vram.mem_out_bus6_2\
        );

    \I__4361\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__4359\ : Sp12to4
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__4358\ : Span12Mux_v
    port map (
            O => \N__18731\,
            I => \N__18728\
        );

    \I__4357\ : Odrv12
    port map (
            O => \N__18728\,
            I => \this_vram.mem_out_bus0_2\
        );

    \I__4356\ : InMux
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__18719\,
            I => \this_vram.mem_out_bus4_2\
        );

    \I__4353\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18710\
        );

    \I__4351\ : Span4Mux_v
    port map (
            O => \N__18710\,
            I => \N__18706\
        );

    \I__4350\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18703\
        );

    \I__4349\ : Sp12to4
    port map (
            O => \N__18706\,
            I => \N__18698\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__18703\,
            I => \N__18698\
        );

    \I__4347\ : Odrv12
    port map (
            O => \N__18698\,
            I => \this_vram.mem_N_109\
        );

    \I__4346\ : SRMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__18692\,
            I => \N__18684\
        );

    \I__4344\ : SRMux
    port map (
            O => \N__18691\,
            I => \N__18681\
        );

    \I__4343\ : SRMux
    port map (
            O => \N__18690\,
            I => \N__18678\
        );

    \I__4342\ : IoInMux
    port map (
            O => \N__18689\,
            I => \N__18674\
        );

    \I__4341\ : SRMux
    port map (
            O => \N__18688\,
            I => \N__18670\
        );

    \I__4340\ : SRMux
    port map (
            O => \N__18687\,
            I => \N__18667\
        );

    \I__4339\ : Span4Mux_s1_v
    port map (
            O => \N__18684\,
            I => \N__18658\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__18681\,
            I => \N__18658\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__18678\,
            I => \N__18658\
        );

    \I__4336\ : SRMux
    port map (
            O => \N__18677\,
            I => \N__18655\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18651\
        );

    \I__4334\ : CascadeMux
    port map (
            O => \N__18673\,
            I => \N__18647\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__18670\,
            I => \N__18641\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18641\
        );

    \I__4331\ : SRMux
    port map (
            O => \N__18666\,
            I => \N__18638\
        );

    \I__4330\ : SRMux
    port map (
            O => \N__18665\,
            I => \N__18635\
        );

    \I__4329\ : Span4Mux_v
    port map (
            O => \N__18658\,
            I => \N__18628\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__18655\,
            I => \N__18628\
        );

    \I__4327\ : SRMux
    port map (
            O => \N__18654\,
            I => \N__18625\
        );

    \I__4326\ : Span4Mux_s2_h
    port map (
            O => \N__18651\,
            I => \N__18619\
        );

    \I__4325\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18614\
        );

    \I__4324\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18614\
        );

    \I__4323\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18611\
        );

    \I__4322\ : Span4Mux_v
    port map (
            O => \N__18641\,
            I => \N__18602\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__18638\,
            I => \N__18602\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__18635\,
            I => \N__18602\
        );

    \I__4319\ : SRMux
    port map (
            O => \N__18634\,
            I => \N__18599\
        );

    \I__4318\ : SRMux
    port map (
            O => \N__18633\,
            I => \N__18596\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__18628\,
            I => \N__18589\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__18625\,
            I => \N__18589\
        );

    \I__4315\ : SRMux
    port map (
            O => \N__18624\,
            I => \N__18586\
        );

    \I__4314\ : SRMux
    port map (
            O => \N__18623\,
            I => \N__18583\
        );

    \I__4313\ : SRMux
    port map (
            O => \N__18622\,
            I => \N__18578\
        );

    \I__4312\ : Sp12to4
    port map (
            O => \N__18619\,
            I => \N__18572\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__18614\,
            I => \N__18567\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__18611\,
            I => \N__18567\
        );

    \I__4309\ : SRMux
    port map (
            O => \N__18610\,
            I => \N__18564\
        );

    \I__4308\ : SRMux
    port map (
            O => \N__18609\,
            I => \N__18559\
        );

    \I__4307\ : Span4Mux_v
    port map (
            O => \N__18602\,
            I => \N__18552\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__18599\,
            I => \N__18552\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__18596\,
            I => \N__18552\
        );

    \I__4304\ : SRMux
    port map (
            O => \N__18595\,
            I => \N__18549\
        );

    \I__4303\ : SRMux
    port map (
            O => \N__18594\,
            I => \N__18546\
        );

    \I__4302\ : Span4Mux_v
    port map (
            O => \N__18589\,
            I => \N__18541\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__18586\,
            I => \N__18541\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__18583\,
            I => \N__18538\
        );

    \I__4299\ : SRMux
    port map (
            O => \N__18582\,
            I => \N__18535\
        );

    \I__4298\ : SRMux
    port map (
            O => \N__18581\,
            I => \N__18532\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__18578\,
            I => \N__18529\
        );

    \I__4296\ : SRMux
    port map (
            O => \N__18577\,
            I => \N__18526\
        );

    \I__4295\ : SRMux
    port map (
            O => \N__18576\,
            I => \N__18523\
        );

    \I__4294\ : SRMux
    port map (
            O => \N__18575\,
            I => \N__18516\
        );

    \I__4293\ : Span12Mux_s9_v
    port map (
            O => \N__18572\,
            I => \N__18511\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__18567\,
            I => \N__18508\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__18564\,
            I => \N__18505\
        );

    \I__4290\ : SRMux
    port map (
            O => \N__18563\,
            I => \N__18502\
        );

    \I__4289\ : SRMux
    port map (
            O => \N__18562\,
            I => \N__18499\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__18559\,
            I => \N__18496\
        );

    \I__4287\ : Span4Mux_v
    port map (
            O => \N__18552\,
            I => \N__18488\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__18549\,
            I => \N__18488\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__18546\,
            I => \N__18488\
        );

    \I__4284\ : Span4Mux_v
    port map (
            O => \N__18541\,
            I => \N__18485\
        );

    \I__4283\ : Span4Mux_s2_v
    port map (
            O => \N__18538\,
            I => \N__18478\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__18535\,
            I => \N__18478\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__18532\,
            I => \N__18478\
        );

    \I__4280\ : Span4Mux_s2_v
    port map (
            O => \N__18529\,
            I => \N__18471\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__18526\,
            I => \N__18471\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__18523\,
            I => \N__18471\
        );

    \I__4277\ : SRMux
    port map (
            O => \N__18522\,
            I => \N__18468\
        );

    \I__4276\ : SRMux
    port map (
            O => \N__18521\,
            I => \N__18465\
        );

    \I__4275\ : SRMux
    port map (
            O => \N__18520\,
            I => \N__18462\
        );

    \I__4274\ : SRMux
    port map (
            O => \N__18519\,
            I => \N__18459\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18456\
        );

    \I__4272\ : SRMux
    port map (
            O => \N__18515\,
            I => \N__18453\
        );

    \I__4271\ : SRMux
    port map (
            O => \N__18514\,
            I => \N__18450\
        );

    \I__4270\ : Span12Mux_h
    port map (
            O => \N__18511\,
            I => \N__18447\
        );

    \I__4269\ : Span4Mux_h
    port map (
            O => \N__18508\,
            I => \N__18444\
        );

    \I__4268\ : Span12Mux_s9_h
    port map (
            O => \N__18505\,
            I => \N__18441\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__18502\,
            I => \N__18438\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__18499\,
            I => \N__18435\
        );

    \I__4265\ : Span12Mux_s9_h
    port map (
            O => \N__18496\,
            I => \N__18432\
        );

    \I__4264\ : SRMux
    port map (
            O => \N__18495\,
            I => \N__18429\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__18488\,
            I => \N__18426\
        );

    \I__4262\ : Span4Mux_v
    port map (
            O => \N__18485\,
            I => \N__18415\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__18478\,
            I => \N__18415\
        );

    \I__4260\ : Span4Mux_v
    port map (
            O => \N__18471\,
            I => \N__18415\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__18468\,
            I => \N__18415\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__18465\,
            I => \N__18415\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__18462\,
            I => \N__18410\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__18459\,
            I => \N__18410\
        );

    \I__4255\ : Span4Mux_h
    port map (
            O => \N__18456\,
            I => \N__18403\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__18453\,
            I => \N__18403\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__18450\,
            I => \N__18403\
        );

    \I__4252\ : Span12Mux_v
    port map (
            O => \N__18447\,
            I => \N__18400\
        );

    \I__4251\ : Span4Mux_h
    port map (
            O => \N__18444\,
            I => \N__18397\
        );

    \I__4250\ : Span12Mux_v
    port map (
            O => \N__18441\,
            I => \N__18392\
        );

    \I__4249\ : Span12Mux_s9_h
    port map (
            O => \N__18438\,
            I => \N__18392\
        );

    \I__4248\ : Span4Mux_h
    port map (
            O => \N__18435\,
            I => \N__18389\
        );

    \I__4247\ : Span12Mux_v
    port map (
            O => \N__18432\,
            I => \N__18384\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__18429\,
            I => \N__18384\
        );

    \I__4245\ : Span4Mux_v
    port map (
            O => \N__18426\,
            I => \N__18375\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__18415\,
            I => \N__18375\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__18410\,
            I => \N__18375\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__18403\,
            I => \N__18375\
        );

    \I__4241\ : Odrv12
    port map (
            O => \N__18400\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__18397\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4239\ : Odrv12
    port map (
            O => \N__18392\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__18389\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4237\ : Odrv12
    port map (
            O => \N__18384\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__18375\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4235\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18358\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__18361\,
            I => \N__18352\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__18358\,
            I => \N__18349\
        );

    \I__4232\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18342\
        );

    \I__4231\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18339\
        );

    \I__4230\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18334\
        );

    \I__4229\ : InMux
    port map (
            O => \N__18352\,
            I => \N__18334\
        );

    \I__4228\ : Span12Mux_h
    port map (
            O => \N__18349\,
            I => \N__18331\
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__18348\,
            I => \N__18328\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18325\
        );

    \I__4225\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18320\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18320\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18315\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18339\,
            I => \N__18315\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__18334\,
            I => \N__18312\
        );

    \I__4220\ : Span12Mux_v
    port map (
            O => \N__18331\,
            I => \N__18307\
        );

    \I__4219\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18304\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__18325\,
            I => \N__18301\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__18320\,
            I => \N__18294\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__18315\,
            I => \N__18294\
        );

    \I__4215\ : Span4Mux_v
    port map (
            O => \N__18312\,
            I => \N__18294\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18289\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18289\
        );

    \I__4212\ : Odrv12
    port map (
            O => \N__18307\,
            I => \this_vga_signals.mult1_un61_sum_axbxc5\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__18304\,
            I => \this_vga_signals.mult1_un61_sum_axbxc5\
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__18301\,
            I => \this_vga_signals.mult1_un61_sum_axbxc5\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__18294\,
            I => \this_vga_signals.mult1_un61_sum_axbxc5\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__18289\,
            I => \this_vga_signals.mult1_un61_sum_axbxc5\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__4206\ : CascadeBuf
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__4204\ : CascadeBuf
    port map (
            O => \N__18269\,
            I => \N__18266\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__18266\,
            I => \N__18263\
        );

    \I__4202\ : CascadeBuf
    port map (
            O => \N__18263\,
            I => \N__18260\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__4200\ : CascadeBuf
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__4198\ : CascadeBuf
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__18248\,
            I => \N__18245\
        );

    \I__4196\ : CascadeBuf
    port map (
            O => \N__18245\,
            I => \N__18242\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__18242\,
            I => \N__18239\
        );

    \I__4194\ : CascadeBuf
    port map (
            O => \N__18239\,
            I => \N__18236\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__4192\ : CascadeBuf
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__4190\ : CascadeBuf
    port map (
            O => \N__18227\,
            I => \N__18224\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__18224\,
            I => \N__18221\
        );

    \I__4188\ : CascadeBuf
    port map (
            O => \N__18221\,
            I => \N__18218\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__18218\,
            I => \N__18215\
        );

    \I__4186\ : CascadeBuf
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__4184\ : CascadeBuf
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__18206\,
            I => \N__18203\
        );

    \I__4182\ : CascadeBuf
    port map (
            O => \N__18203\,
            I => \N__18200\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__4180\ : CascadeBuf
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18191\
        );

    \I__4178\ : CascadeBuf
    port map (
            O => \N__18191\,
            I => \N__18188\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__18179\,
            I => \M_this_vga_signals_address_5\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__4171\ : Span4Mux_v
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__18167\,
            I => \this_vram.mem_out_bus1_2\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18164\,
            I => \N__18161\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__4167\ : Span4Mux_v
    port map (
            O => \N__18158\,
            I => \N__18155\
        );

    \I__4166\ : Span4Mux_v
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__18152\,
            I => \this_vram.mem_out_bus5_2\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__4162\ : Span4Mux_v
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__18140\,
            I => \N__18137\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__18137\,
            I => \this_vram.mem_out_bus1_1\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__4157\ : Sp12to4
    port map (
            O => \N__18128\,
            I => \N__18125\
        );

    \I__4156\ : Odrv12
    port map (
            O => \N__18125\,
            I => \this_vram.mem_out_bus5_1\
        );

    \I__4155\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__18113\,
            I => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__4149\ : Span4Mux_v
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__4148\ : Span4Mux_v
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__18098\,
            I => \this_vram.mem_out_bus6_0\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__4144\ : Span4Mux_v
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__18086\,
            I => \this_vram.mem_out_bus2_0\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__18083\,
            I => \this_vram.mem_mem_2_0_RNIU0NZ0Z11_cascade_\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18076\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18073\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18076\,
            I => \N__18068\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__18073\,
            I => \N__18068\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__4136\ : Span4Mux_h
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__18062\,
            I => \this_vram.mem_N_112\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__18053\,
            I => \this_vram.mem_out_bus4_0\
        );

    \I__4131\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__4129\ : Sp12to4
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__4128\ : Span12Mux_v
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__4127\ : Odrv12
    port map (
            O => \N__18038\,
            I => \this_vram.mem_out_bus0_0\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__18032\,
            I => \this_vram.mem_mem_0_0_RNIQOIZ0Z11\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18026\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__18026\,
            I => \this_vram.mem_out_bus3_2\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__4120\ : Sp12to4
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__4119\ : Span12Mux_v
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__4118\ : Odrv12
    port map (
            O => \N__18011\,
            I => \this_vram.mem_out_bus7_2\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__18005\,
            I => \N__18002\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__4114\ : Sp12to4
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__4113\ : Odrv12
    port map (
            O => \N__17996\,
            I => \this_vram.mem_out_bus6_1\
        );

    \I__4112\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__17987\,
            I => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\
        );

    \I__4109\ : CEMux
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__17981\,
            I => \N__17977\
        );

    \I__4107\ : CEMux
    port map (
            O => \N__17980\,
            I => \N__17974\
        );

    \I__4106\ : Span4Mux_h
    port map (
            O => \N__17977\,
            I => \N__17971\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__17974\,
            I => \N__17968\
        );

    \I__4104\ : Sp12to4
    port map (
            O => \N__17971\,
            I => \N__17965\
        );

    \I__4103\ : Span4Mux_h
    port map (
            O => \N__17968\,
            I => \N__17962\
        );

    \I__4102\ : Span12Mux_v
    port map (
            O => \N__17965\,
            I => \N__17959\
        );

    \I__4101\ : Sp12to4
    port map (
            O => \N__17962\,
            I => \N__17956\
        );

    \I__4100\ : Odrv12
    port map (
            O => \N__17959\,
            I => \this_vram.mem_WE_14\
        );

    \I__4099\ : Odrv12
    port map (
            O => \N__17956\,
            I => \this_vram.mem_WE_14\
        );

    \I__4098\ : CEMux
    port map (
            O => \N__17951\,
            I => \N__17948\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__17948\,
            I => \N__17944\
        );

    \I__4096\ : CEMux
    port map (
            O => \N__17947\,
            I => \N__17941\
        );

    \I__4095\ : Span4Mux_v
    port map (
            O => \N__17944\,
            I => \N__17938\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__17941\,
            I => \N__17935\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__17938\,
            I => \N__17932\
        );

    \I__4092\ : Span4Mux_h
    port map (
            O => \N__17935\,
            I => \N__17929\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__17932\,
            I => \this_vram.mem_WE_10\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__17929\,
            I => \this_vram.mem_WE_10\
        );

    \I__4089\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__17921\,
            I => \M_this_vram_read_data_3\
        );

    \I__4087\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__4085\ : Odrv4
    port map (
            O => \N__17912\,
            I => \this_vram.mem_out_bus4_1\
        );

    \I__4084\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__17906\,
            I => \N__17903\
        );

    \I__4082\ : Span12Mux_h
    port map (
            O => \N__17903\,
            I => \N__17900\
        );

    \I__4081\ : Span12Mux_v
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__4080\ : Odrv12
    port map (
            O => \N__17897\,
            I => \this_vram.mem_out_bus0_1\
        );

    \I__4079\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17891\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__17891\,
            I => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0\
        );

    \I__4077\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__17882\,
            I => \N__17879\
        );

    \I__4074\ : Sp12to4
    port map (
            O => \N__17879\,
            I => \N__17876\
        );

    \I__4073\ : Span12Mux_v
    port map (
            O => \N__17876\,
            I => \N__17873\
        );

    \I__4072\ : Odrv12
    port map (
            O => \N__17873\,
            I => \this_vram.mem_out_bus7_3\
        );

    \I__4071\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17867\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__4069\ : Span4Mux_v
    port map (
            O => \N__17864\,
            I => \N__17861\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__17861\,
            I => \this_vram.mem_out_bus3_3\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__17858\,
            I => \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_\
        );

    \I__4066\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__17852\,
            I => \this_vram.mem_N_102\
        );

    \I__4064\ : InMux
    port map (
            O => \N__17849\,
            I => \N__17845\
        );

    \I__4063\ : InMux
    port map (
            O => \N__17848\,
            I => \N__17842\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__17845\,
            I => \N__17838\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__17842\,
            I => \N__17834\
        );

    \I__4060\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17831\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__17838\,
            I => \N__17827\
        );

    \I__4058\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17824\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__17834\,
            I => \N__17819\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__17831\,
            I => \N__17819\
        );

    \I__4055\ : InMux
    port map (
            O => \N__17830\,
            I => \N__17816\
        );

    \I__4054\ : Span4Mux_h
    port map (
            O => \N__17827\,
            I => \N__17811\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__17824\,
            I => \N__17811\
        );

    \I__4052\ : Span4Mux_h
    port map (
            O => \N__17819\,
            I => \N__17806\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17806\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__17811\,
            I => \N__17803\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__17806\,
            I => \N__17800\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__17803\,
            I => \N__17795\
        );

    \I__4047\ : Span4Mux_v
    port map (
            O => \N__17800\,
            I => \N__17792\
        );

    \I__4046\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17789\
        );

    \I__4045\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17786\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__17795\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__17792\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__17789\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__17786\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__4040\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17774\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__17774\,
            I => \M_this_vram_read_data_2\
        );

    \I__4038\ : CEMux
    port map (
            O => \N__17771\,
            I => \N__17768\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__17768\,
            I => \N__17764\
        );

    \I__4036\ : CEMux
    port map (
            O => \N__17767\,
            I => \N__17761\
        );

    \I__4035\ : Span4Mux_v
    port map (
            O => \N__17764\,
            I => \N__17756\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__17761\,
            I => \N__17756\
        );

    \I__4033\ : Span4Mux_v
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__4032\ : Span4Mux_v
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__4031\ : Span4Mux_v
    port map (
            O => \N__17750\,
            I => \N__17747\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__17747\,
            I => \this_vram.mem_WE_12\
        );

    \I__4029\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17734\
        );

    \I__4027\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17731\
        );

    \I__4026\ : IoInMux
    port map (
            O => \N__17739\,
            I => \N__17728\
        );

    \I__4025\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17724\
        );

    \I__4024\ : CascadeMux
    port map (
            O => \N__17737\,
            I => \N__17721\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__17734\,
            I => \N__17716\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__17731\,
            I => \N__17716\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17713\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__17727\,
            I => \N__17706\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__17724\,
            I => \N__17703\
        );

    \I__4018\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17700\
        );

    \I__4017\ : Sp12to4
    port map (
            O => \N__17716\,
            I => \N__17697\
        );

    \I__4016\ : Span4Mux_s2_v
    port map (
            O => \N__17713\,
            I => \N__17694\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__17712\,
            I => \N__17691\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__17711\,
            I => \N__17688\
        );

    \I__4013\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17682\
        );

    \I__4012\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17679\
        );

    \I__4011\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17676\
        );

    \I__4010\ : Span4Mux_v
    port map (
            O => \N__17703\,
            I => \N__17673\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__17700\,
            I => \N__17670\
        );

    \I__4008\ : Span12Mux_v
    port map (
            O => \N__17697\,
            I => \N__17665\
        );

    \I__4007\ : Sp12to4
    port map (
            O => \N__17694\,
            I => \N__17665\
        );

    \I__4006\ : InMux
    port map (
            O => \N__17691\,
            I => \N__17658\
        );

    \I__4005\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17658\
        );

    \I__4004\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17658\
        );

    \I__4003\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17653\
        );

    \I__4002\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17653\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__17682\,
            I => \N__17646\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__17679\,
            I => \N__17646\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__17676\,
            I => \N__17646\
        );

    \I__3998\ : Span4Mux_h
    port map (
            O => \N__17673\,
            I => \N__17641\
        );

    \I__3997\ : Span4Mux_v
    port map (
            O => \N__17670\,
            I => \N__17641\
        );

    \I__3996\ : Span12Mux_h
    port map (
            O => \N__17665\,
            I => \N__17638\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__17658\,
            I => \M_this_reset_cond_out_0\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__17653\,
            I => \M_this_reset_cond_out_0\
        );

    \I__3993\ : Odrv12
    port map (
            O => \N__17646\,
            I => \M_this_reset_cond_out_0\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__17641\,
            I => \M_this_reset_cond_out_0\
        );

    \I__3991\ : Odrv12
    port map (
            O => \N__17638\,
            I => \M_this_reset_cond_out_0\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__17627\,
            I => \N__17620\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__17626\,
            I => \N__17616\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17625\,
            I => \N__17609\
        );

    \I__3987\ : InMux
    port map (
            O => \N__17624\,
            I => \N__17599\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17599\
        );

    \I__3985\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17592\
        );

    \I__3984\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17592\
        );

    \I__3983\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17592\
        );

    \I__3982\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17589\
        );

    \I__3981\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17584\
        );

    \I__3980\ : InMux
    port map (
            O => \N__17613\,
            I => \N__17584\
        );

    \I__3979\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17581\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__17609\,
            I => \N__17578\
        );

    \I__3977\ : InMux
    port map (
            O => \N__17608\,
            I => \N__17575\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17607\,
            I => \N__17570\
        );

    \I__3975\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17570\
        );

    \I__3974\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17562\
        );

    \I__3973\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17562\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__17599\,
            I => \N__17557\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__17592\,
            I => \N__17557\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__17589\,
            I => \N__17546\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__17584\,
            I => \N__17546\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__17581\,
            I => \N__17546\
        );

    \I__3967\ : Span4Mux_v
    port map (
            O => \N__17578\,
            I => \N__17546\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__17575\,
            I => \N__17546\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__17570\,
            I => \N__17543\
        );

    \I__3964\ : InMux
    port map (
            O => \N__17569\,
            I => \N__17540\
        );

    \I__3963\ : InMux
    port map (
            O => \N__17568\,
            I => \N__17537\
        );

    \I__3962\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17534\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__17562\,
            I => \N__17531\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__17557\,
            I => \N__17528\
        );

    \I__3959\ : Span4Mux_h
    port map (
            O => \N__17546\,
            I => \N__17525\
        );

    \I__3958\ : Span4Mux_v
    port map (
            O => \N__17543\,
            I => \N__17520\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17520\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17537\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__17534\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__3954\ : Odrv12
    port map (
            O => \N__17531\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__17528\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__3952\ : Odrv4
    port map (
            O => \N__17525\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__17520\,
            I => \M_this_start_data_delay_out_0\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__17507\,
            I => \M_state_q_ns_1_0__i12_mux_cascade_\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__17504\,
            I => \N__17496\
        );

    \I__3948\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17493\
        );

    \I__3947\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17490\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__17501\,
            I => \N__17487\
        );

    \I__3945\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17472\
        );

    \I__3944\ : InMux
    port map (
            O => \N__17499\,
            I => \N__17472\
        );

    \I__3943\ : InMux
    port map (
            O => \N__17496\,
            I => \N__17469\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__17493\,
            I => \N__17464\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__17490\,
            I => \N__17464\
        );

    \I__3940\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17457\
        );

    \I__3939\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17457\
        );

    \I__3938\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17457\
        );

    \I__3937\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17454\
        );

    \I__3936\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17446\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17446\
        );

    \I__3934\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17443\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17480\,
            I => \N__17434\
        );

    \I__3932\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17434\
        );

    \I__3931\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17434\
        );

    \I__3930\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17434\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17431\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17426\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__17464\,
            I => \N__17426\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__17457\,
            I => \N__17421\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17421\
        );

    \I__3924\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17418\
        );

    \I__3923\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17415\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17451\,
            I => \N__17412\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__17446\,
            I => \N__17407\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__17443\,
            I => \N__17407\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__17434\,
            I => \N__17404\
        );

    \I__3918\ : Span4Mux_h
    port map (
            O => \N__17431\,
            I => \N__17401\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__17426\,
            I => \N__17396\
        );

    \I__3916\ : Span4Mux_h
    port map (
            O => \N__17421\,
            I => \N__17396\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__17418\,
            I => \N__17393\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__17415\,
            I => \M_state_qZ0Z_1\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__17412\,
            I => \M_state_qZ0Z_1\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__17407\,
            I => \M_state_qZ0Z_1\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__17404\,
            I => \M_state_qZ0Z_1\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__17401\,
            I => \M_state_qZ0Z_1\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__17396\,
            I => \M_state_qZ0Z_1\
        );

    \I__3908\ : Odrv12
    port map (
            O => \N__17393\,
            I => \M_state_qZ0Z_1\
        );

    \I__3907\ : ClkMux
    port map (
            O => \N__17378\,
            I => \N__17147\
        );

    \I__3906\ : ClkMux
    port map (
            O => \N__17377\,
            I => \N__17147\
        );

    \I__3905\ : ClkMux
    port map (
            O => \N__17376\,
            I => \N__17147\
        );

    \I__3904\ : ClkMux
    port map (
            O => \N__17375\,
            I => \N__17147\
        );

    \I__3903\ : ClkMux
    port map (
            O => \N__17374\,
            I => \N__17147\
        );

    \I__3902\ : ClkMux
    port map (
            O => \N__17373\,
            I => \N__17147\
        );

    \I__3901\ : ClkMux
    port map (
            O => \N__17372\,
            I => \N__17147\
        );

    \I__3900\ : ClkMux
    port map (
            O => \N__17371\,
            I => \N__17147\
        );

    \I__3899\ : ClkMux
    port map (
            O => \N__17370\,
            I => \N__17147\
        );

    \I__3898\ : ClkMux
    port map (
            O => \N__17369\,
            I => \N__17147\
        );

    \I__3897\ : ClkMux
    port map (
            O => \N__17368\,
            I => \N__17147\
        );

    \I__3896\ : ClkMux
    port map (
            O => \N__17367\,
            I => \N__17147\
        );

    \I__3895\ : ClkMux
    port map (
            O => \N__17366\,
            I => \N__17147\
        );

    \I__3894\ : ClkMux
    port map (
            O => \N__17365\,
            I => \N__17147\
        );

    \I__3893\ : ClkMux
    port map (
            O => \N__17364\,
            I => \N__17147\
        );

    \I__3892\ : ClkMux
    port map (
            O => \N__17363\,
            I => \N__17147\
        );

    \I__3891\ : ClkMux
    port map (
            O => \N__17362\,
            I => \N__17147\
        );

    \I__3890\ : ClkMux
    port map (
            O => \N__17361\,
            I => \N__17147\
        );

    \I__3889\ : ClkMux
    port map (
            O => \N__17360\,
            I => \N__17147\
        );

    \I__3888\ : ClkMux
    port map (
            O => \N__17359\,
            I => \N__17147\
        );

    \I__3887\ : ClkMux
    port map (
            O => \N__17358\,
            I => \N__17147\
        );

    \I__3886\ : ClkMux
    port map (
            O => \N__17357\,
            I => \N__17147\
        );

    \I__3885\ : ClkMux
    port map (
            O => \N__17356\,
            I => \N__17147\
        );

    \I__3884\ : ClkMux
    port map (
            O => \N__17355\,
            I => \N__17147\
        );

    \I__3883\ : ClkMux
    port map (
            O => \N__17354\,
            I => \N__17147\
        );

    \I__3882\ : ClkMux
    port map (
            O => \N__17353\,
            I => \N__17147\
        );

    \I__3881\ : ClkMux
    port map (
            O => \N__17352\,
            I => \N__17147\
        );

    \I__3880\ : ClkMux
    port map (
            O => \N__17351\,
            I => \N__17147\
        );

    \I__3879\ : ClkMux
    port map (
            O => \N__17350\,
            I => \N__17147\
        );

    \I__3878\ : ClkMux
    port map (
            O => \N__17349\,
            I => \N__17147\
        );

    \I__3877\ : ClkMux
    port map (
            O => \N__17348\,
            I => \N__17147\
        );

    \I__3876\ : ClkMux
    port map (
            O => \N__17347\,
            I => \N__17147\
        );

    \I__3875\ : ClkMux
    port map (
            O => \N__17346\,
            I => \N__17147\
        );

    \I__3874\ : ClkMux
    port map (
            O => \N__17345\,
            I => \N__17147\
        );

    \I__3873\ : ClkMux
    port map (
            O => \N__17344\,
            I => \N__17147\
        );

    \I__3872\ : ClkMux
    port map (
            O => \N__17343\,
            I => \N__17147\
        );

    \I__3871\ : ClkMux
    port map (
            O => \N__17342\,
            I => \N__17147\
        );

    \I__3870\ : ClkMux
    port map (
            O => \N__17341\,
            I => \N__17147\
        );

    \I__3869\ : ClkMux
    port map (
            O => \N__17340\,
            I => \N__17147\
        );

    \I__3868\ : ClkMux
    port map (
            O => \N__17339\,
            I => \N__17147\
        );

    \I__3867\ : ClkMux
    port map (
            O => \N__17338\,
            I => \N__17147\
        );

    \I__3866\ : ClkMux
    port map (
            O => \N__17337\,
            I => \N__17147\
        );

    \I__3865\ : ClkMux
    port map (
            O => \N__17336\,
            I => \N__17147\
        );

    \I__3864\ : ClkMux
    port map (
            O => \N__17335\,
            I => \N__17147\
        );

    \I__3863\ : ClkMux
    port map (
            O => \N__17334\,
            I => \N__17147\
        );

    \I__3862\ : ClkMux
    port map (
            O => \N__17333\,
            I => \N__17147\
        );

    \I__3861\ : ClkMux
    port map (
            O => \N__17332\,
            I => \N__17147\
        );

    \I__3860\ : ClkMux
    port map (
            O => \N__17331\,
            I => \N__17147\
        );

    \I__3859\ : ClkMux
    port map (
            O => \N__17330\,
            I => \N__17147\
        );

    \I__3858\ : ClkMux
    port map (
            O => \N__17329\,
            I => \N__17147\
        );

    \I__3857\ : ClkMux
    port map (
            O => \N__17328\,
            I => \N__17147\
        );

    \I__3856\ : ClkMux
    port map (
            O => \N__17327\,
            I => \N__17147\
        );

    \I__3855\ : ClkMux
    port map (
            O => \N__17326\,
            I => \N__17147\
        );

    \I__3854\ : ClkMux
    port map (
            O => \N__17325\,
            I => \N__17147\
        );

    \I__3853\ : ClkMux
    port map (
            O => \N__17324\,
            I => \N__17147\
        );

    \I__3852\ : ClkMux
    port map (
            O => \N__17323\,
            I => \N__17147\
        );

    \I__3851\ : ClkMux
    port map (
            O => \N__17322\,
            I => \N__17147\
        );

    \I__3850\ : ClkMux
    port map (
            O => \N__17321\,
            I => \N__17147\
        );

    \I__3849\ : ClkMux
    port map (
            O => \N__17320\,
            I => \N__17147\
        );

    \I__3848\ : ClkMux
    port map (
            O => \N__17319\,
            I => \N__17147\
        );

    \I__3847\ : ClkMux
    port map (
            O => \N__17318\,
            I => \N__17147\
        );

    \I__3846\ : ClkMux
    port map (
            O => \N__17317\,
            I => \N__17147\
        );

    \I__3845\ : ClkMux
    port map (
            O => \N__17316\,
            I => \N__17147\
        );

    \I__3844\ : ClkMux
    port map (
            O => \N__17315\,
            I => \N__17147\
        );

    \I__3843\ : ClkMux
    port map (
            O => \N__17314\,
            I => \N__17147\
        );

    \I__3842\ : ClkMux
    port map (
            O => \N__17313\,
            I => \N__17147\
        );

    \I__3841\ : ClkMux
    port map (
            O => \N__17312\,
            I => \N__17147\
        );

    \I__3840\ : ClkMux
    port map (
            O => \N__17311\,
            I => \N__17147\
        );

    \I__3839\ : ClkMux
    port map (
            O => \N__17310\,
            I => \N__17147\
        );

    \I__3838\ : ClkMux
    port map (
            O => \N__17309\,
            I => \N__17147\
        );

    \I__3837\ : ClkMux
    port map (
            O => \N__17308\,
            I => \N__17147\
        );

    \I__3836\ : ClkMux
    port map (
            O => \N__17307\,
            I => \N__17147\
        );

    \I__3835\ : ClkMux
    port map (
            O => \N__17306\,
            I => \N__17147\
        );

    \I__3834\ : ClkMux
    port map (
            O => \N__17305\,
            I => \N__17147\
        );

    \I__3833\ : ClkMux
    port map (
            O => \N__17304\,
            I => \N__17147\
        );

    \I__3832\ : ClkMux
    port map (
            O => \N__17303\,
            I => \N__17147\
        );

    \I__3831\ : ClkMux
    port map (
            O => \N__17302\,
            I => \N__17147\
        );

    \I__3830\ : GlobalMux
    port map (
            O => \N__17147\,
            I => \N__17144\
        );

    \I__3829\ : gio2CtrlBuf
    port map (
            O => \N__17144\,
            I => clk_c_g
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__17141\,
            I => \N__17137\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17131\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17128\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__17131\,
            I => \N__17125\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__17128\,
            I => \N__17122\
        );

    \I__3822\ : Span12Mux_h
    port map (
            O => \N__17125\,
            I => \N__17119\
        );

    \I__3821\ : Span12Mux_h
    port map (
            O => \N__17122\,
            I => \N__17116\
        );

    \I__3820\ : Odrv12
    port map (
            O => \N__17119\,
            I => port_data_c_0
        );

    \I__3819\ : Odrv12
    port map (
            O => \N__17116\,
            I => port_data_c_0
        );

    \I__3818\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__17108\,
            I => \N__17104\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17101\
        );

    \I__3815\ : Span4Mux_s2_v
    port map (
            O => \N__17104\,
            I => \N__17095\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__17101\,
            I => \N__17095\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17092\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__17095\,
            I => \N__17086\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__3810\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17083\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__17086\,
            I => \N__17077\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17082\,
            I => \N__17074\
        );

    \I__3806\ : Span4Mux_v
    port map (
            O => \N__17077\,
            I => \N__17067\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17074\,
            I => \N__17067\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17064\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17060\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__17067\,
            I => \N__17055\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__17064\,
            I => \N__17055\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17063\,
            I => \N__17052\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__17060\,
            I => \N__17049\
        );

    \I__3798\ : Span4Mux_v
    port map (
            O => \N__17055\,
            I => \N__17044\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17052\,
            I => \N__17044\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__17049\,
            I => \N__17039\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__17044\,
            I => \N__17039\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__17039\,
            I => \M_this_vram_write_data_0\
        );

    \I__3793\ : CEMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17033\,
            I => \N__17029\
        );

    \I__3791\ : CEMux
    port map (
            O => \N__17032\,
            I => \N__17026\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__17029\,
            I => \N__17023\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__17026\,
            I => \N__17020\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__17023\,
            I => \this_vram.mem_WE_8\
        );

    \I__3787\ : Odrv12
    port map (
            O => \N__17020\,
            I => \this_vram.mem_WE_8\
        );

    \I__3786\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17012\,
            I => \N__17008\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17011\,
            I => \N__17005\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__17008\,
            I => \N__17000\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17005\,
            I => \N__17000\
        );

    \I__3781\ : Sp12to4
    port map (
            O => \N__17000\,
            I => \N__16996\
        );

    \I__3780\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16993\
        );

    \I__3779\ : Span12Mux_v
    port map (
            O => \N__16996\,
            I => \N__16988\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__16993\,
            I => \N__16988\
        );

    \I__3777\ : Odrv12
    port map (
            O => \N__16988\,
            I => \this_vram.mem_N_91\
        );

    \I__3776\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16981\
        );

    \I__3775\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16978\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__16981\,
            I => \N__16972\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__16978\,
            I => \N__16972\
        );

    \I__3772\ : InMux
    port map (
            O => \N__16977\,
            I => \N__16969\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__16972\,
            I => \N__16966\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__16969\,
            I => \N__16963\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__16966\,
            I => \N__16958\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__16963\,
            I => \N__16958\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__16955\,
            I => \this_vram.mem_N_88\
        );

    \I__3765\ : InMux
    port map (
            O => \N__16952\,
            I => \N__16948\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__16951\,
            I => \N__16945\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__16948\,
            I => \N__16942\
        );

    \I__3762\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__3761\ : Span4Mux_h
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__16939\,
            I => \N__16933\
        );

    \I__3759\ : Span4Mux_h
    port map (
            O => \N__16936\,
            I => \N__16930\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__16933\,
            I => \N__16927\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__16930\,
            I => \N_16_0\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__16927\,
            I => \N_16_0\
        );

    \I__3755\ : InMux
    port map (
            O => \N__16922\,
            I => \N__16919\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__3753\ : Span12Mux_s9_v
    port map (
            O => \N__16916\,
            I => \N__16913\
        );

    \I__3752\ : Odrv12
    port map (
            O => \N__16913\,
            I => port_address_c_4
        );

    \I__3751\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__16907\,
            I => \N__16904\
        );

    \I__3749\ : Span12Mux_v
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__3748\ : Span12Mux_v
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__3747\ : Odrv12
    port map (
            O => \N__16898\,
            I => port_address_c_7
        );

    \I__3746\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16888\
        );

    \I__3745\ : InMux
    port map (
            O => \N__16894\,
            I => \N__16888\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__16893\,
            I => \N__16884\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__16888\,
            I => \N__16881\
        );

    \I__3742\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16878\
        );

    \I__3741\ : InMux
    port map (
            O => \N__16884\,
            I => \N__16875\
        );

    \I__3740\ : Span4Mux_v
    port map (
            O => \N__16881\,
            I => \N__16870\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__16878\,
            I => \N__16870\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__16875\,
            I => \N__16867\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__16870\,
            I => \N__16864\
        );

    \I__3736\ : Span12Mux_v
    port map (
            O => \N__16867\,
            I => \N__16859\
        );

    \I__3735\ : Sp12to4
    port map (
            O => \N__16864\,
            I => \N__16859\
        );

    \I__3734\ : Span12Mux_h
    port map (
            O => \N__16859\,
            I => \N__16856\
        );

    \I__3733\ : Odrv12
    port map (
            O => \N__16856\,
            I => port_enb_c
        );

    \I__3732\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16850\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__16850\,
            I => \N__16847\
        );

    \I__3730\ : Span12Mux_v
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__3729\ : Odrv12
    port map (
            O => \N__16844\,
            I => port_address_c_2
        );

    \I__3728\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__16838\,
            I => \M_state_q_ns_1_0__m7Z0Z_5\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__16835\,
            I => \N__16831\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__16834\,
            I => \N__16827\
        );

    \I__3724\ : InMux
    port map (
            O => \N__16831\,
            I => \N__16824\
        );

    \I__3723\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16821\
        );

    \I__3722\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16818\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__16824\,
            I => \N__16815\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__16821\,
            I => \N__16810\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__16818\,
            I => \N__16810\
        );

    \I__3718\ : Span4Mux_v
    port map (
            O => \N__16815\,
            I => \N__16807\
        );

    \I__3717\ : Span4Mux_v
    port map (
            O => \N__16810\,
            I => \N__16804\
        );

    \I__3716\ : Sp12to4
    port map (
            O => \N__16807\,
            I => \N__16799\
        );

    \I__3715\ : Sp12to4
    port map (
            O => \N__16804\,
            I => \N__16799\
        );

    \I__3714\ : Span12Mux_h
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__3713\ : Odrv12
    port map (
            O => \N__16796\,
            I => port_data_c_1
        );

    \I__3712\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__16790\,
            I => \N__16786\
        );

    \I__3710\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16783\
        );

    \I__3709\ : Span4Mux_h
    port map (
            O => \N__16786\,
            I => \N__16779\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__16783\,
            I => \N__16776\
        );

    \I__3707\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16773\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__16779\,
            I => \N__16767\
        );

    \I__3705\ : Span4Mux_h
    port map (
            O => \N__16776\,
            I => \N__16767\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__16773\,
            I => \N__16764\
        );

    \I__3703\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16761\
        );

    \I__3702\ : Span4Mux_v
    port map (
            O => \N__16767\,
            I => \N__16755\
        );

    \I__3701\ : Span4Mux_h
    port map (
            O => \N__16764\,
            I => \N__16755\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__16761\,
            I => \N__16752\
        );

    \I__3699\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16749\
        );

    \I__3698\ : Span4Mux_v
    port map (
            O => \N__16755\,
            I => \N__16742\
        );

    \I__3697\ : Span4Mux_h
    port map (
            O => \N__16752\,
            I => \N__16742\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__16749\,
            I => \N__16739\
        );

    \I__3695\ : InMux
    port map (
            O => \N__16748\,
            I => \N__16736\
        );

    \I__3694\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16733\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__16742\,
            I => \N__16727\
        );

    \I__3692\ : Span4Mux_h
    port map (
            O => \N__16739\,
            I => \N__16727\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__16736\,
            I => \N__16724\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__16733\,
            I => \N__16721\
        );

    \I__3689\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16718\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__16727\,
            I => \N__16713\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__16724\,
            I => \N__16713\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__16721\,
            I => \N__16708\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__16718\,
            I => \N__16708\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__16713\,
            I => \M_this_vram_write_data_1\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__16708\,
            I => \M_this_vram_write_data_1\
        );

    \I__3682\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16700\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__16700\,
            I => \N__16697\
        );

    \I__3680\ : Span4Mux_v
    port map (
            O => \N__16697\,
            I => \N__16694\
        );

    \I__3679\ : Span4Mux_v
    port map (
            O => \N__16694\,
            I => \N__16691\
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__16691\,
            I => \this_vram.mem_out_bus2_1\
        );

    \I__3677\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__16685\,
            I => \N__16682\
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__16682\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_17\
        );

    \I__3674\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16676\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__16676\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_18\
        );

    \I__3672\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__16670\,
            I => \M_this_start_address_delay_out_0\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__16667\,
            I => \M_state_q_ns_1_0__N_24_mux_cascade_\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__16664\,
            I => \M_state_q_ns_1_0__N_10_cascade_\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__3667\ : CascadeBuf
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3665\ : CascadeBuf
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3663\ : CascadeBuf
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__3661\ : CascadeBuf
    port map (
            O => \N__16640\,
            I => \N__16637\
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__3659\ : CascadeBuf
    port map (
            O => \N__16634\,
            I => \N__16631\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \N__16628\
        );

    \I__3657\ : CascadeBuf
    port map (
            O => \N__16628\,
            I => \N__16625\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__3655\ : CascadeBuf
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__3654\ : CascadeMux
    port map (
            O => \N__16619\,
            I => \N__16616\
        );

    \I__3653\ : CascadeBuf
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__3651\ : CascadeBuf
    port map (
            O => \N__16610\,
            I => \N__16607\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__3649\ : CascadeBuf
    port map (
            O => \N__16604\,
            I => \N__16601\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3647\ : CascadeBuf
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__3645\ : CascadeBuf
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__16589\,
            I => \N__16586\
        );

    \I__3643\ : CascadeBuf
    port map (
            O => \N__16586\,
            I => \N__16583\
        );

    \I__3642\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3641\ : CascadeBuf
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__16577\,
            I => \N__16574\
        );

    \I__3639\ : CascadeBuf
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__16571\,
            I => \N__16568\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16563\
        );

    \I__3636\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16560\
        );

    \I__3635\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16557\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__16563\,
            I => \N__16554\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__16560\,
            I => \N__16551\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__16557\,
            I => \N__16546\
        );

    \I__3631\ : Span12Mux_s7_v
    port map (
            O => \N__16554\,
            I => \N__16546\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__16551\,
            I => \M_current_address_qZ0Z_1\
        );

    \I__3629\ : Odrv12
    port map (
            O => \N__16546\,
            I => \M_current_address_qZ0Z_1\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__16532\,
            I => \this_start_data_delay.this_edge_detector.N_211\
        );

    \I__3624\ : CascadeMux
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__3623\ : CascadeBuf
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__3621\ : CascadeBuf
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3619\ : CascadeBuf
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__16511\,
            I => \N__16508\
        );

    \I__3617\ : CascadeBuf
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3615\ : CascadeBuf
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__16499\,
            I => \N__16496\
        );

    \I__3613\ : CascadeBuf
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__3611\ : CascadeBuf
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__3609\ : CascadeBuf
    port map (
            O => \N__16484\,
            I => \N__16481\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__16481\,
            I => \N__16478\
        );

    \I__3607\ : CascadeBuf
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__16475\,
            I => \N__16472\
        );

    \I__3605\ : CascadeBuf
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__3603\ : CascadeBuf
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__3601\ : CascadeBuf
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__16457\,
            I => \N__16454\
        );

    \I__3599\ : CascadeBuf
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3597\ : CascadeBuf
    port map (
            O => \N__16448\,
            I => \N__16445\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__16445\,
            I => \N__16442\
        );

    \I__3595\ : CascadeBuf
    port map (
            O => \N__16442\,
            I => \N__16439\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__16439\,
            I => \N__16436\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16433\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__16433\,
            I => \N__16429\
        );

    \I__3591\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16426\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__16429\,
            I => \N__16423\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__16426\,
            I => \N__16417\
        );

    \I__3588\ : Span4Mux_v
    port map (
            O => \N__16423\,
            I => \N__16417\
        );

    \I__3587\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16414\
        );

    \I__3586\ : Span4Mux_v
    port map (
            O => \N__16417\,
            I => \N__16411\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__16414\,
            I => \M_current_address_qZ0Z_4\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__16411\,
            I => \M_current_address_qZ0Z_4\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16402\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__16405\,
            I => \N__16399\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16402\,
            I => \N__16396\
        );

    \I__3580\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16393\
        );

    \I__3579\ : Span4Mux_v
    port map (
            O => \N__16396\,
            I => \N__16390\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__16393\,
            I => \N__16387\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__16390\,
            I => \N__16384\
        );

    \I__3576\ : Sp12to4
    port map (
            O => \N__16387\,
            I => \N__16381\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__16384\,
            I => \N__16378\
        );

    \I__3574\ : Span12Mux_v
    port map (
            O => \N__16381\,
            I => \N__16375\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__16378\,
            I => port_data_c_4
        );

    \I__3572\ : Odrv12
    port map (
            O => \N__16375\,
            I => port_data_c_4
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \N__16367\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16364\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__3568\ : Span4Mux_v
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__16358\,
            I => \this_start_data_delay.this_edge_detector.N_214\
        );

    \I__3566\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__16352\,
            I => \N__16348\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16351\,
            I => \N__16345\
        );

    \I__3563\ : Span4Mux_h
    port map (
            O => \N__16348\,
            I => \N__16327\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__16345\,
            I => \N__16327\
        );

    \I__3561\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16322\
        );

    \I__3560\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16322\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16342\,
            I => \N__16315\
        );

    \I__3558\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16315\
        );

    \I__3557\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16315\
        );

    \I__3556\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16312\
        );

    \I__3555\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16309\
        );

    \I__3554\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16302\
        );

    \I__3553\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16302\
        );

    \I__3552\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16302\
        );

    \I__3551\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16297\
        );

    \I__3550\ : InMux
    port map (
            O => \N__16333\,
            I => \N__16297\
        );

    \I__3549\ : InMux
    port map (
            O => \N__16332\,
            I => \N__16276\
        );

    \I__3548\ : Span4Mux_h
    port map (
            O => \N__16327\,
            I => \N__16265\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__16322\,
            I => \N__16265\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__16315\,
            I => \N__16265\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__16312\,
            I => \N__16265\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__16309\,
            I => \N__16265\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16302\,
            I => \N__16260\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__16297\,
            I => \N__16260\
        );

    \I__3541\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16257\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16246\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16246\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16246\
        );

    \I__3537\ : InMux
    port map (
            O => \N__16292\,
            I => \N__16246\
        );

    \I__3536\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16246\
        );

    \I__3535\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16243\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16236\
        );

    \I__3533\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16236\
        );

    \I__3532\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16236\
        );

    \I__3531\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16229\
        );

    \I__3530\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16229\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16229\
        );

    \I__3528\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16222\
        );

    \I__3527\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16222\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16222\
        );

    \I__3525\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16217\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16217\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__16276\,
            I => \N__16214\
        );

    \I__3522\ : Span4Mux_v
    port map (
            O => \N__16265\,
            I => \N__16207\
        );

    \I__3521\ : Span4Mux_v
    port map (
            O => \N__16260\,
            I => \N__16207\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__16257\,
            I => \N__16207\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__16246\,
            I => \M_state_qZ0Z_0\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__16243\,
            I => \M_state_qZ0Z_0\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__16236\,
            I => \M_state_qZ0Z_0\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__16229\,
            I => \M_state_qZ0Z_0\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16222\,
            I => \M_state_qZ0Z_0\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16217\,
            I => \M_state_qZ0Z_0\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__16214\,
            I => \M_state_qZ0Z_0\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__16207\,
            I => \M_state_qZ0Z_0\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16187\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__3509\ : Span12Mux_h
    port map (
            O => \N__16184\,
            I => \N__16181\
        );

    \I__3508\ : Odrv12
    port map (
            O => \N__16181\,
            I => port_address_c_1
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__16178\,
            I => \N__16175\
        );

    \I__3506\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16172\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__16172\,
            I => \M_state_q_ns_1_0__N_24_mux\
        );

    \I__3504\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__16166\,
            I => \N__16162\
        );

    \I__3502\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16159\
        );

    \I__3501\ : Span4Mux_v
    port map (
            O => \N__16162\,
            I => \N__16154\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__16159\,
            I => \N__16154\
        );

    \I__3499\ : Sp12to4
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__3498\ : Span12Mux_h
    port map (
            O => \N__16151\,
            I => \N__16148\
        );

    \I__3497\ : Odrv12
    port map (
            O => \N__16148\,
            I => port_address_c_0
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__16145\,
            I => \N__16142\
        );

    \I__3495\ : CascadeBuf
    port map (
            O => \N__16142\,
            I => \N__16139\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__16139\,
            I => \N__16136\
        );

    \I__3493\ : CascadeBuf
    port map (
            O => \N__16136\,
            I => \N__16133\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__16133\,
            I => \N__16130\
        );

    \I__3491\ : CascadeBuf
    port map (
            O => \N__16130\,
            I => \N__16127\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__3489\ : CascadeBuf
    port map (
            O => \N__16124\,
            I => \N__16121\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__16121\,
            I => \N__16118\
        );

    \I__3487\ : CascadeBuf
    port map (
            O => \N__16118\,
            I => \N__16115\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__16115\,
            I => \N__16112\
        );

    \I__3485\ : CascadeBuf
    port map (
            O => \N__16112\,
            I => \N__16109\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__16109\,
            I => \N__16106\
        );

    \I__3483\ : CascadeBuf
    port map (
            O => \N__16106\,
            I => \N__16103\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__16103\,
            I => \N__16100\
        );

    \I__3481\ : CascadeBuf
    port map (
            O => \N__16100\,
            I => \N__16097\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__16097\,
            I => \N__16094\
        );

    \I__3479\ : CascadeBuf
    port map (
            O => \N__16094\,
            I => \N__16091\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__16091\,
            I => \N__16088\
        );

    \I__3477\ : CascadeBuf
    port map (
            O => \N__16088\,
            I => \N__16085\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__3475\ : CascadeBuf
    port map (
            O => \N__16082\,
            I => \N__16079\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__16079\,
            I => \N__16076\
        );

    \I__3473\ : CascadeBuf
    port map (
            O => \N__16076\,
            I => \N__16073\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__16073\,
            I => \N__16070\
        );

    \I__3471\ : CascadeBuf
    port map (
            O => \N__16070\,
            I => \N__16067\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__16067\,
            I => \N__16064\
        );

    \I__3469\ : CascadeBuf
    port map (
            O => \N__16064\,
            I => \N__16061\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__3467\ : CascadeBuf
    port map (
            O => \N__16058\,
            I => \N__16055\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__16055\,
            I => \N__16052\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16049\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__16049\,
            I => \N__16046\
        );

    \I__3463\ : Span4Mux_v
    port map (
            O => \N__16046\,
            I => \N__16042\
        );

    \I__3462\ : InMux
    port map (
            O => \N__16045\,
            I => \N__16038\
        );

    \I__3461\ : Span4Mux_h
    port map (
            O => \N__16042\,
            I => \N__16035\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16041\,
            I => \N__16032\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16038\,
            I => \N__16027\
        );

    \I__3458\ : Span4Mux_v
    port map (
            O => \N__16035\,
            I => \N__16027\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__16032\,
            I => \M_current_address_qZ0Z_8\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__16027\,
            I => \M_current_address_qZ0Z_8\
        );

    \I__3455\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__16019\,
            I => \N__16016\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__16016\,
            I => \this_start_data_delay.this_edge_detector.N_218\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__3451\ : CascadeBuf
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__3449\ : CascadeBuf
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__3447\ : CascadeBuf
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__3445\ : CascadeBuf
    port map (
            O => \N__15992\,
            I => \N__15989\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__3443\ : CascadeBuf
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__3441\ : CascadeBuf
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__15977\,
            I => \N__15974\
        );

    \I__3439\ : CascadeBuf
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__3437\ : CascadeBuf
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__15965\,
            I => \N__15962\
        );

    \I__3435\ : CascadeBuf
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__15959\,
            I => \N__15956\
        );

    \I__3433\ : CascadeBuf
    port map (
            O => \N__15956\,
            I => \N__15953\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__15953\,
            I => \N__15950\
        );

    \I__3431\ : CascadeBuf
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__3429\ : CascadeBuf
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__15941\,
            I => \N__15938\
        );

    \I__3427\ : CascadeBuf
    port map (
            O => \N__15938\,
            I => \N__15935\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__15935\,
            I => \N__15932\
        );

    \I__3425\ : CascadeBuf
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__3424\ : CascadeMux
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__3423\ : CascadeBuf
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__3421\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15917\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__15917\,
            I => \N__15914\
        );

    \I__3419\ : Span4Mux_s3_v
    port map (
            O => \N__15914\,
            I => \N__15910\
        );

    \I__3418\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15906\
        );

    \I__3417\ : Span4Mux_h
    port map (
            O => \N__15910\,
            I => \N__15903\
        );

    \I__3416\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15900\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__15906\,
            I => \N__15895\
        );

    \I__3414\ : Span4Mux_v
    port map (
            O => \N__15903\,
            I => \N__15895\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__15900\,
            I => \M_current_address_qZ0Z_10\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__15895\,
            I => \M_current_address_qZ0Z_10\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__15890\,
            I => \N__15887\
        );

    \I__3410\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__15884\,
            I => \this_start_data_delay.this_edge_detector.N_220\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__15881\,
            I => \N__15878\
        );

    \I__3407\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15875\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__15875\,
            I => \N__15872\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__15872\,
            I => \this_start_data_delay.this_edge_detector.N_221\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__15869\,
            I => \N__15865\
        );

    \I__3403\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15862\
        );

    \I__3402\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15859\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__15862\,
            I => \N__15854\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__15859\,
            I => \N__15854\
        );

    \I__3399\ : Span12Mux_s9_v
    port map (
            O => \N__15854\,
            I => \N__15851\
        );

    \I__3398\ : Span12Mux_v
    port map (
            O => \N__15851\,
            I => \N__15848\
        );

    \I__3397\ : Span12Mux_h
    port map (
            O => \N__15848\,
            I => \N__15845\
        );

    \I__3396\ : Odrv12
    port map (
            O => \N__15845\,
            I => port_data_c_6
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__15842\,
            I => \N__15839\
        );

    \I__3394\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15836\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__15836\,
            I => \this_start_data_delay.this_edge_detector.N_223\
        );

    \I__3392\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15830\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__15830\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_15\
        );

    \I__3390\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15824\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__15824\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_16\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__15821\,
            I => \N__15818\
        );

    \I__3387\ : CascadeBuf
    port map (
            O => \N__15818\,
            I => \N__15815\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__3385\ : CascadeBuf
    port map (
            O => \N__15812\,
            I => \N__15809\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__15809\,
            I => \N__15806\
        );

    \I__3383\ : CascadeBuf
    port map (
            O => \N__15806\,
            I => \N__15803\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__15803\,
            I => \N__15800\
        );

    \I__3381\ : CascadeBuf
    port map (
            O => \N__15800\,
            I => \N__15797\
        );

    \I__3380\ : CascadeMux
    port map (
            O => \N__15797\,
            I => \N__15794\
        );

    \I__3379\ : CascadeBuf
    port map (
            O => \N__15794\,
            I => \N__15791\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__15791\,
            I => \N__15788\
        );

    \I__3377\ : CascadeBuf
    port map (
            O => \N__15788\,
            I => \N__15785\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__15785\,
            I => \N__15782\
        );

    \I__3375\ : CascadeBuf
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__3373\ : CascadeBuf
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__3371\ : CascadeBuf
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__3369\ : CascadeBuf
    port map (
            O => \N__15764\,
            I => \N__15761\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__3367\ : CascadeBuf
    port map (
            O => \N__15758\,
            I => \N__15755\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__3365\ : CascadeBuf
    port map (
            O => \N__15752\,
            I => \N__15749\
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__3363\ : CascadeBuf
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__15743\,
            I => \N__15740\
        );

    \I__3361\ : CascadeBuf
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__15737\,
            I => \N__15734\
        );

    \I__3359\ : CascadeBuf
    port map (
            O => \N__15734\,
            I => \N__15731\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__15731\,
            I => \N__15728\
        );

    \I__3357\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15725\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__15725\,
            I => \N__15722\
        );

    \I__3355\ : Span4Mux_s2_v
    port map (
            O => \N__15722\,
            I => \N__15718\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__15721\,
            I => \N__15715\
        );

    \I__3353\ : Span4Mux_h
    port map (
            O => \N__15718\,
            I => \N__15711\
        );

    \I__3352\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15708\
        );

    \I__3351\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15705\
        );

    \I__3350\ : Span4Mux_v
    port map (
            O => \N__15711\,
            I => \N__15702\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__15708\,
            I => \M_current_address_qZ0Z_7\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__15705\,
            I => \M_current_address_qZ0Z_7\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__15702\,
            I => \M_current_address_qZ0Z_7\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__3345\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__15689\,
            I => \this_start_data_delay.this_edge_detector.N_217\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__3342\ : CascadeBuf
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__3340\ : CascadeBuf
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__3338\ : CascadeBuf
    port map (
            O => \N__15671\,
            I => \N__15668\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__3336\ : CascadeBuf
    port map (
            O => \N__15665\,
            I => \N__15662\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__15662\,
            I => \N__15659\
        );

    \I__3334\ : CascadeBuf
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__3332\ : CascadeBuf
    port map (
            O => \N__15653\,
            I => \N__15650\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__15650\,
            I => \N__15647\
        );

    \I__3330\ : CascadeBuf
    port map (
            O => \N__15647\,
            I => \N__15644\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__15644\,
            I => \N__15641\
        );

    \I__3328\ : CascadeBuf
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__3326\ : CascadeBuf
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__3324\ : CascadeBuf
    port map (
            O => \N__15629\,
            I => \N__15626\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__15626\,
            I => \N__15623\
        );

    \I__3322\ : CascadeBuf
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__15620\,
            I => \N__15617\
        );

    \I__3320\ : CascadeBuf
    port map (
            O => \N__15617\,
            I => \N__15614\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__15614\,
            I => \N__15611\
        );

    \I__3318\ : CascadeBuf
    port map (
            O => \N__15611\,
            I => \N__15608\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__15608\,
            I => \N__15605\
        );

    \I__3316\ : CascadeBuf
    port map (
            O => \N__15605\,
            I => \N__15602\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__15602\,
            I => \N__15599\
        );

    \I__3314\ : CascadeBuf
    port map (
            O => \N__15599\,
            I => \N__15596\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__15596\,
            I => \N__15593\
        );

    \I__3312\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15590\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__15590\,
            I => \N__15587\
        );

    \I__3310\ : Span4Mux_s3_v
    port map (
            O => \N__15587\,
            I => \N__15584\
        );

    \I__3309\ : Span4Mux_h
    port map (
            O => \N__15584\,
            I => \N__15579\
        );

    \I__3308\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15576\
        );

    \I__3307\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15573\
        );

    \I__3306\ : Span4Mux_v
    port map (
            O => \N__15579\,
            I => \N__15570\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__15576\,
            I => \M_current_address_qZ0Z_0\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__15573\,
            I => \M_current_address_qZ0Z_0\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__15570\,
            I => \M_current_address_qZ0Z_0\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__3301\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15557\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__15557\,
            I => \this_start_data_delay.this_edge_detector.N_210\
        );

    \I__3299\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15551\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__15551\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_13\
        );

    \I__3297\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15545\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__15545\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_14\
        );

    \I__3295\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15539\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__15539\,
            I => \M_current_address_q_RNIHDTUZ0Z_0\
        );

    \I__3293\ : InMux
    port map (
            O => \N__15536\,
            I => \N__15533\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__15533\,
            I => \un1_M_current_address_q_cry_5_c_RNIC9GNZ0\
        );

    \I__3291\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15527\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__15527\,
            I => \un1_M_current_address_q_cry_6_c_RNIECHNZ0\
        );

    \I__3289\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15521\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15521\,
            I => \un1_M_current_address_q_cry_10_c_RNI4KKHZ0\
        );

    \I__3287\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__15515\,
            I => \un1_M_current_address_q_cry_2_c_RNI60DNZ0\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15500\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15497\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15494\
        );

    \I__3282\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15491\
        );

    \I__3281\ : InMux
    port map (
            O => \N__15508\,
            I => \N__15488\
        );

    \I__3280\ : InMux
    port map (
            O => \N__15507\,
            I => \N__15485\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15506\,
            I => \N__15480\
        );

    \I__3278\ : InMux
    port map (
            O => \N__15505\,
            I => \N__15480\
        );

    \I__3277\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15477\
        );

    \I__3276\ : InMux
    port map (
            O => \N__15503\,
            I => \N__15474\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__15500\,
            I => \N__15459\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__15497\,
            I => \N__15456\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__15494\,
            I => \N__15453\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__15491\,
            I => \N__15450\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__15488\,
            I => \N__15447\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__15485\,
            I => \N__15444\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__15480\,
            I => \N__15441\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__15477\,
            I => \N__15438\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15474\,
            I => \N__15435\
        );

    \I__3266\ : SRMux
    port map (
            O => \N__15473\,
            I => \N__15392\
        );

    \I__3265\ : SRMux
    port map (
            O => \N__15472\,
            I => \N__15392\
        );

    \I__3264\ : SRMux
    port map (
            O => \N__15471\,
            I => \N__15392\
        );

    \I__3263\ : SRMux
    port map (
            O => \N__15470\,
            I => \N__15392\
        );

    \I__3262\ : SRMux
    port map (
            O => \N__15469\,
            I => \N__15392\
        );

    \I__3261\ : SRMux
    port map (
            O => \N__15468\,
            I => \N__15392\
        );

    \I__3260\ : SRMux
    port map (
            O => \N__15467\,
            I => \N__15392\
        );

    \I__3259\ : SRMux
    port map (
            O => \N__15466\,
            I => \N__15392\
        );

    \I__3258\ : SRMux
    port map (
            O => \N__15465\,
            I => \N__15392\
        );

    \I__3257\ : SRMux
    port map (
            O => \N__15464\,
            I => \N__15392\
        );

    \I__3256\ : SRMux
    port map (
            O => \N__15463\,
            I => \N__15392\
        );

    \I__3255\ : SRMux
    port map (
            O => \N__15462\,
            I => \N__15392\
        );

    \I__3254\ : Glb2LocalMux
    port map (
            O => \N__15459\,
            I => \N__15392\
        );

    \I__3253\ : Glb2LocalMux
    port map (
            O => \N__15456\,
            I => \N__15392\
        );

    \I__3252\ : Glb2LocalMux
    port map (
            O => \N__15453\,
            I => \N__15392\
        );

    \I__3251\ : Glb2LocalMux
    port map (
            O => \N__15450\,
            I => \N__15392\
        );

    \I__3250\ : Glb2LocalMux
    port map (
            O => \N__15447\,
            I => \N__15392\
        );

    \I__3249\ : Glb2LocalMux
    port map (
            O => \N__15444\,
            I => \N__15392\
        );

    \I__3248\ : Glb2LocalMux
    port map (
            O => \N__15441\,
            I => \N__15392\
        );

    \I__3247\ : Glb2LocalMux
    port map (
            O => \N__15438\,
            I => \N__15392\
        );

    \I__3246\ : Glb2LocalMux
    port map (
            O => \N__15435\,
            I => \N__15392\
        );

    \I__3245\ : GlobalMux
    port map (
            O => \N__15392\,
            I => \N__15389\
        );

    \I__3244\ : gio2CtrlBuf
    port map (
            O => \N__15389\,
            I => \N_339_g\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__15386\,
            I => \N__15383\
        );

    \I__3242\ : CascadeBuf
    port map (
            O => \N__15383\,
            I => \N__15380\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__3240\ : CascadeBuf
    port map (
            O => \N__15377\,
            I => \N__15374\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \N__15371\
        );

    \I__3238\ : CascadeBuf
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__3236\ : CascadeBuf
    port map (
            O => \N__15365\,
            I => \N__15362\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__3234\ : CascadeBuf
    port map (
            O => \N__15359\,
            I => \N__15356\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__3232\ : CascadeBuf
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__15350\,
            I => \N__15347\
        );

    \I__3230\ : CascadeBuf
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__15344\,
            I => \N__15341\
        );

    \I__3228\ : CascadeBuf
    port map (
            O => \N__15341\,
            I => \N__15338\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \N__15335\
        );

    \I__3226\ : CascadeBuf
    port map (
            O => \N__15335\,
            I => \N__15332\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__15332\,
            I => \N__15329\
        );

    \I__3224\ : CascadeBuf
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__15326\,
            I => \N__15323\
        );

    \I__3222\ : CascadeBuf
    port map (
            O => \N__15323\,
            I => \N__15320\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__3220\ : CascadeBuf
    port map (
            O => \N__15317\,
            I => \N__15314\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__15314\,
            I => \N__15311\
        );

    \I__3218\ : CascadeBuf
    port map (
            O => \N__15311\,
            I => \N__15308\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__15308\,
            I => \N__15305\
        );

    \I__3216\ : CascadeBuf
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__15302\,
            I => \N__15299\
        );

    \I__3214\ : CascadeBuf
    port map (
            O => \N__15299\,
            I => \N__15296\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__15296\,
            I => \N__15293\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15290\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15290\,
            I => \N__15285\
        );

    \I__3210\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15282\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15279\
        );

    \I__3208\ : Span12Mux_h
    port map (
            O => \N__15285\,
            I => \N__15276\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__15282\,
            I => \M_current_address_qZ0Z_6\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__15279\,
            I => \M_current_address_qZ0Z_6\
        );

    \I__3205\ : Odrv12
    port map (
            O => \N__15276\,
            I => \M_current_address_qZ0Z_6\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15266\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__15266\,
            I => \this_start_data_delay.this_edge_detector.N_216\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__3201\ : CascadeBuf
    port map (
            O => \N__15260\,
            I => \N__15257\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \N__15254\
        );

    \I__3199\ : CascadeBuf
    port map (
            O => \N__15254\,
            I => \N__15251\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__15251\,
            I => \N__15248\
        );

    \I__3197\ : CascadeBuf
    port map (
            O => \N__15248\,
            I => \N__15245\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__3195\ : CascadeBuf
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__3193\ : CascadeBuf
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__3191\ : CascadeBuf
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__15227\,
            I => \N__15224\
        );

    \I__3189\ : CascadeBuf
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__15221\,
            I => \N__15218\
        );

    \I__3187\ : CascadeBuf
    port map (
            O => \N__15218\,
            I => \N__15215\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__15215\,
            I => \N__15212\
        );

    \I__3185\ : CascadeBuf
    port map (
            O => \N__15212\,
            I => \N__15209\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \N__15206\
        );

    \I__3183\ : CascadeBuf
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__15203\,
            I => \N__15200\
        );

    \I__3181\ : CascadeBuf
    port map (
            O => \N__15200\,
            I => \N__15197\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__15197\,
            I => \N__15194\
        );

    \I__3179\ : CascadeBuf
    port map (
            O => \N__15194\,
            I => \N__15191\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__15191\,
            I => \N__15188\
        );

    \I__3177\ : CascadeBuf
    port map (
            O => \N__15188\,
            I => \N__15185\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__15185\,
            I => \N__15182\
        );

    \I__3175\ : CascadeBuf
    port map (
            O => \N__15182\,
            I => \N__15179\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__15179\,
            I => \N__15176\
        );

    \I__3173\ : CascadeBuf
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__15173\,
            I => \N__15170\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15164\
        );

    \I__3169\ : Span4Mux_s2_v
    port map (
            O => \N__15164\,
            I => \N__15161\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__15161\,
            I => \N__15156\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15160\,
            I => \N__15153\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15150\
        );

    \I__3165\ : Span4Mux_v
    port map (
            O => \N__15156\,
            I => \N__15147\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15153\,
            I => \M_current_address_qZ0Z_3\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__15150\,
            I => \M_current_address_qZ0Z_3\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__15147\,
            I => \M_current_address_qZ0Z_3\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__15140\,
            I => \N__15137\
        );

    \I__3160\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15134\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__15134\,
            I => \this_start_data_delay.this_edge_detector.N_213\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15131\,
            I => \N__15128\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__15128\,
            I => \N__15125\
        );

    \I__3156\ : Odrv12
    port map (
            O => \N__15125\,
            I => \un1_M_current_address_q_cry_11_c_RNI6NLHZ0\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15122\,
            I => \un1_M_current_address_q_cry_11\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15119\,
            I => \un1_M_current_address_q_cry_12\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__15116\,
            I => \N__15112\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15115\,
            I => \N__15109\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15106\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15109\,
            I => \N_177_0\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__15106\,
            I => \N_177_0\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15098\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15098\,
            I => \un1_M_current_address_q_cry_9_c_RNIRDIMZ0\
        );

    \I__3146\ : InMux
    port map (
            O => \N__15095\,
            I => \N__15092\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15092\,
            I => \N__15089\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__15089\,
            I => \un1_M_current_address_q_cry_0_c_RNI2QANZ0\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15083\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__15083\,
            I => \un1_M_current_address_q_cry_12_c_RNI8QMHZ0\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__15077\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_12\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15071\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_10\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__15065\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_11\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15062\,
            I => \un1_M_current_address_q_cry_2\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15056\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15056\,
            I => \un1_M_current_address_q_cry_3_c_RNI83ENZ0\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15053\,
            I => \un1_M_current_address_q_cry_3\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__15050\,
            I => \N__15047\
        );

    \I__3130\ : CascadeBuf
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__15044\,
            I => \N__15041\
        );

    \I__3128\ : CascadeBuf
    port map (
            O => \N__15041\,
            I => \N__15038\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__15038\,
            I => \N__15035\
        );

    \I__3126\ : CascadeBuf
    port map (
            O => \N__15035\,
            I => \N__15032\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__3124\ : CascadeBuf
    port map (
            O => \N__15029\,
            I => \N__15026\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__15026\,
            I => \N__15023\
        );

    \I__3122\ : CascadeBuf
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__15020\,
            I => \N__15017\
        );

    \I__3120\ : CascadeBuf
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__15014\,
            I => \N__15011\
        );

    \I__3118\ : CascadeBuf
    port map (
            O => \N__15011\,
            I => \N__15008\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__15008\,
            I => \N__15005\
        );

    \I__3116\ : CascadeBuf
    port map (
            O => \N__15005\,
            I => \N__15002\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__3114\ : CascadeBuf
    port map (
            O => \N__14999\,
            I => \N__14996\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__3112\ : CascadeBuf
    port map (
            O => \N__14993\,
            I => \N__14990\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__14990\,
            I => \N__14987\
        );

    \I__3110\ : CascadeBuf
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__14984\,
            I => \N__14981\
        );

    \I__3108\ : CascadeBuf
    port map (
            O => \N__14981\,
            I => \N__14978\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__3106\ : CascadeBuf
    port map (
            O => \N__14975\,
            I => \N__14972\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__3104\ : CascadeBuf
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__14966\,
            I => \N__14963\
        );

    \I__3102\ : CascadeBuf
    port map (
            O => \N__14963\,
            I => \N__14960\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__14960\,
            I => \N__14957\
        );

    \I__3100\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14954\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__14954\,
            I => \N__14951\
        );

    \I__3098\ : Span4Mux_s3_v
    port map (
            O => \N__14951\,
            I => \N__14946\
        );

    \I__3097\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14943\
        );

    \I__3096\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14940\
        );

    \I__3095\ : Sp12to4
    port map (
            O => \N__14946\,
            I => \N__14937\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__14943\,
            I => \N__14934\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__14940\,
            I => \N__14929\
        );

    \I__3092\ : Span12Mux_h
    port map (
            O => \N__14937\,
            I => \N__14929\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__14934\,
            I => \M_current_address_qZ0Z_5\
        );

    \I__3090\ : Odrv12
    port map (
            O => \N__14929\,
            I => \M_current_address_qZ0Z_5\
        );

    \I__3089\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__14921\,
            I => \un1_M_current_address_q_cry_4_c_RNIA6FNZ0\
        );

    \I__3087\ : InMux
    port map (
            O => \N__14918\,
            I => \un1_M_current_address_q_cry_4\
        );

    \I__3086\ : InMux
    port map (
            O => \N__14915\,
            I => \un1_M_current_address_q_cry_5\
        );

    \I__3085\ : InMux
    port map (
            O => \N__14912\,
            I => \un1_M_current_address_q_cry_6\
        );

    \I__3084\ : InMux
    port map (
            O => \N__14909\,
            I => \N__14906\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__14906\,
            I => \un1_M_current_address_q_cry_7_c_RNIGFINZ0\
        );

    \I__3082\ : InMux
    port map (
            O => \N__14903\,
            I => \bfn_19_24_0_\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \N__14897\
        );

    \I__3080\ : CascadeBuf
    port map (
            O => \N__14897\,
            I => \N__14894\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__3078\ : CascadeBuf
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__3076\ : CascadeBuf
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__3074\ : CascadeBuf
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__3072\ : CascadeBuf
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__14870\,
            I => \N__14867\
        );

    \I__3070\ : CascadeBuf
    port map (
            O => \N__14867\,
            I => \N__14864\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__3068\ : CascadeBuf
    port map (
            O => \N__14861\,
            I => \N__14858\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__14858\,
            I => \N__14855\
        );

    \I__3066\ : CascadeBuf
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__14852\,
            I => \N__14849\
        );

    \I__3064\ : CascadeBuf
    port map (
            O => \N__14849\,
            I => \N__14846\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__3062\ : CascadeBuf
    port map (
            O => \N__14843\,
            I => \N__14840\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__14840\,
            I => \N__14837\
        );

    \I__3060\ : CascadeBuf
    port map (
            O => \N__14837\,
            I => \N__14834\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__14834\,
            I => \N__14831\
        );

    \I__3058\ : CascadeBuf
    port map (
            O => \N__14831\,
            I => \N__14828\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__3056\ : CascadeBuf
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__3054\ : CascadeBuf
    port map (
            O => \N__14819\,
            I => \N__14816\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__3052\ : CascadeBuf
    port map (
            O => \N__14813\,
            I => \N__14810\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__3050\ : InMux
    port map (
            O => \N__14807\,
            I => \N__14804\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__14801\,
            I => \N__14796\
        );

    \I__3047\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14793\
        );

    \I__3046\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14790\
        );

    \I__3045\ : Span4Mux_h
    port map (
            O => \N__14796\,
            I => \N__14787\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__14793\,
            I => \N__14784\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__14790\,
            I => \N__14779\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__14787\,
            I => \N__14779\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__14784\,
            I => \M_current_address_qZ0Z_9\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__14779\,
            I => \M_current_address_qZ0Z_9\
        );

    \I__3039\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__14771\,
            I => \un1_M_current_address_q_cry_8_c_RNIIIJNZ0\
        );

    \I__3037\ : InMux
    port map (
            O => \N__14768\,
            I => \un1_M_current_address_q_cry_8\
        );

    \I__3036\ : InMux
    port map (
            O => \N__14765\,
            I => \un1_M_current_address_q_cry_9\
        );

    \I__3035\ : InMux
    port map (
            O => \N__14762\,
            I => \un1_M_current_address_q_cry_10\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14756\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__14756\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_8\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__14753\,
            I => \N__14749\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__14752\,
            I => \N__14746\
        );

    \I__3030\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14743\
        );

    \I__3029\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14740\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__14743\,
            I => \N__14735\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__14740\,
            I => \N__14735\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__3025\ : Sp12to4
    port map (
            O => \N__14732\,
            I => \N__14729\
        );

    \I__3024\ : Span12Mux_h
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__3023\ : Odrv12
    port map (
            O => \N__14726\,
            I => port_data_c_5
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__14723\,
            I => \N__14720\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__14717\,
            I => \this_start_data_delay.this_edge_detector.N_222\
        );

    \I__3019\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__14711\,
            I => \N__14708\
        );

    \I__3017\ : Span4Mux_h
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__14705\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_6\
        );

    \I__3015\ : InMux
    port map (
            O => \N__14702\,
            I => \N__14699\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__14699\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_7\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14693\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__14693\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_9\
        );

    \I__3011\ : InMux
    port map (
            O => \N__14690\,
            I => \un1_M_current_address_q_cry_0\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__3009\ : CascadeBuf
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__3007\ : CascadeBuf
    port map (
            O => \N__14678\,
            I => \N__14675\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__3005\ : CascadeBuf
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__3003\ : CascadeBuf
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__3001\ : CascadeBuf
    port map (
            O => \N__14660\,
            I => \N__14657\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__2999\ : CascadeBuf
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__2997\ : CascadeBuf
    port map (
            O => \N__14648\,
            I => \N__14645\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__2995\ : CascadeBuf
    port map (
            O => \N__14642\,
            I => \N__14639\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__14639\,
            I => \N__14636\
        );

    \I__2993\ : CascadeBuf
    port map (
            O => \N__14636\,
            I => \N__14633\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__14633\,
            I => \N__14630\
        );

    \I__2991\ : CascadeBuf
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__2989\ : CascadeBuf
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__2987\ : CascadeBuf
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__2985\ : CascadeBuf
    port map (
            O => \N__14612\,
            I => \N__14609\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__14609\,
            I => \N__14606\
        );

    \I__2983\ : CascadeBuf
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__2981\ : CascadeBuf
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14594\,
            I => \N__14590\
        );

    \I__2978\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14586\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__14590\,
            I => \N__14583\
        );

    \I__2976\ : InMux
    port map (
            O => \N__14589\,
            I => \N__14580\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__14586\,
            I => \N__14577\
        );

    \I__2974\ : Span12Mux_s9_v
    port map (
            O => \N__14583\,
            I => \N__14574\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__14580\,
            I => \M_current_address_qZ0Z_2\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__14577\,
            I => \M_current_address_qZ0Z_2\
        );

    \I__2971\ : Odrv12
    port map (
            O => \N__14574\,
            I => \M_current_address_qZ0Z_2\
        );

    \I__2970\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14564\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__14564\,
            I => \un1_M_current_address_q_cry_1_c_RNI4TBNZ0\
        );

    \I__2968\ : InMux
    port map (
            O => \N__14561\,
            I => \un1_M_current_address_q_cry_1\
        );

    \I__2967\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14555\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__14555\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_17\
        );

    \I__2965\ : InMux
    port map (
            O => \N__14552\,
            I => \N__14549\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__14549\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_18\
        );

    \I__2963\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14543\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__14543\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_7\
        );

    \I__2961\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14537\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__14537\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_8\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__14534\,
            I => \N__14531\
        );

    \I__2958\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14528\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__14525\,
            I => \this_start_data_delay.this_edge_detector.N_215\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__14522\,
            I => \N__14519\
        );

    \I__2954\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N__14513\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__14513\,
            I => \this_start_data_delay.this_edge_detector.N_212\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__14510\,
            I => \N__14507\
        );

    \I__2950\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14504\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__14504\,
            I => \this_start_data_delay.this_edge_detector.N_219\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__14501\,
            I => \N__14497\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__14500\,
            I => \N__14494\
        );

    \I__2946\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14491\
        );

    \I__2945\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14488\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14491\,
            I => \N__14485\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14482\
        );

    \I__2942\ : Span4Mux_h
    port map (
            O => \N__14485\,
            I => \N__14479\
        );

    \I__2941\ : Span4Mux_h
    port map (
            O => \N__14482\,
            I => \N__14476\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__14479\,
            I => \N__14473\
        );

    \I__2939\ : Span4Mux_h
    port map (
            O => \N__14476\,
            I => \N__14470\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__14473\,
            I => \this_vram.N_17_0\
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__14470\,
            I => \this_vram.N_17_0\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__14462\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_11\
        );

    \I__2934\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14456\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__14456\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_12\
        );

    \I__2932\ : IoInMux
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14447\
        );

    \I__2930\ : Span12Mux_s7_v
    port map (
            O => \N__14447\,
            I => \N__14444\
        );

    \I__2929\ : Span12Mux_h
    port map (
            O => \N__14444\,
            I => \N__14441\
        );

    \I__2928\ : Span12Mux_v
    port map (
            O => \N__14441\,
            I => \N__14438\
        );

    \I__2927\ : Odrv12
    port map (
            O => \N__14438\,
            I => debug_d
        );

    \I__2926\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14432\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__14432\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_13\
        );

    \I__2924\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14426\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14426\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_14\
        );

    \I__2922\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14420\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__14420\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_15\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__14414\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_16\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14408\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__14408\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_3\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14405\,
            I => \N__14402\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__14402\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_4\
        );

    \I__2914\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14396\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__14396\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_10\
        );

    \I__2912\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14390\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__14390\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_9\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14384\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__14384\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_6\
        );

    \I__2908\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14378\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14378\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_4\
        );

    \I__2906\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14372\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__14372\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_5\
        );

    \I__2904\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14365\
        );

    \I__2903\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14362\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__14365\,
            I => \N__14359\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__14362\,
            I => \N__14354\
        );

    \I__2900\ : Span4Mux_h
    port map (
            O => \N__14359\,
            I => \N__14345\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14342\
        );

    \I__2898\ : InMux
    port map (
            O => \N__14357\,
            I => \N__14339\
        );

    \I__2897\ : Span4Mux_h
    port map (
            O => \N__14354\,
            I => \N__14336\
        );

    \I__2896\ : InMux
    port map (
            O => \N__14353\,
            I => \N__14333\
        );

    \I__2895\ : InMux
    port map (
            O => \N__14352\,
            I => \N__14330\
        );

    \I__2894\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14327\
        );

    \I__2893\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14322\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14349\,
            I => \N__14322\
        );

    \I__2891\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14319\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__14345\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__14342\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__14339\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__14336\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__14333\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__14330\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__14327\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14322\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__14319\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__2881\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14296\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14293\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14296\,
            I => \N__14290\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14293\,
            I => \N__14281\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__14290\,
            I => \N__14278\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14289\,
            I => \N__14275\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14268\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14287\,
            I => \N__14268\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14286\,
            I => \N__14268\
        );

    \I__2872\ : InMux
    port map (
            O => \N__14285\,
            I => \N__14263\
        );

    \I__2871\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14263\
        );

    \I__2870\ : Odrv12
    port map (
            O => \N__14281\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__14278\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__14275\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__14268\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__14263\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__14252\,
            I => \N__14249\
        );

    \I__2864\ : CascadeBuf
    port map (
            O => \N__14249\,
            I => \N__14246\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__14246\,
            I => \N__14243\
        );

    \I__2862\ : CascadeBuf
    port map (
            O => \N__14243\,
            I => \N__14240\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__14240\,
            I => \N__14237\
        );

    \I__2860\ : CascadeBuf
    port map (
            O => \N__14237\,
            I => \N__14234\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__14234\,
            I => \N__14231\
        );

    \I__2858\ : CascadeBuf
    port map (
            O => \N__14231\,
            I => \N__14228\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__14228\,
            I => \N__14225\
        );

    \I__2856\ : CascadeBuf
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__14222\,
            I => \N__14219\
        );

    \I__2854\ : CascadeBuf
    port map (
            O => \N__14219\,
            I => \N__14216\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__14216\,
            I => \N__14213\
        );

    \I__2852\ : CascadeBuf
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__14210\,
            I => \N__14207\
        );

    \I__2850\ : CascadeBuf
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__14204\,
            I => \N__14201\
        );

    \I__2848\ : CascadeBuf
    port map (
            O => \N__14201\,
            I => \N__14198\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__14198\,
            I => \N__14195\
        );

    \I__2846\ : CascadeBuf
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__14192\,
            I => \N__14189\
        );

    \I__2844\ : CascadeBuf
    port map (
            O => \N__14189\,
            I => \N__14186\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__14186\,
            I => \N__14183\
        );

    \I__2842\ : CascadeBuf
    port map (
            O => \N__14183\,
            I => \N__14180\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__14180\,
            I => \N__14177\
        );

    \I__2840\ : CascadeBuf
    port map (
            O => \N__14177\,
            I => \N__14174\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__14174\,
            I => \N__14171\
        );

    \I__2838\ : CascadeBuf
    port map (
            O => \N__14171\,
            I => \N__14168\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__14168\,
            I => \N__14165\
        );

    \I__2836\ : CascadeBuf
    port map (
            O => \N__14165\,
            I => \N__14162\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__14162\,
            I => \N__14159\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14156\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14156\,
            I => \N__14153\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__14153\,
            I => \N__14150\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__14150\,
            I => \N__14147\
        );

    \I__2830\ : Span4Mux_v
    port map (
            O => \N__14147\,
            I => \N__14144\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__14144\,
            I => \M_this_vga_signals_address_10\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__14135\,
            I => \this_vram.M_this_vram_read_data_0\
        );

    \I__2825\ : InMux
    port map (
            O => \N__14132\,
            I => \N__14126\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14126\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__14126\,
            I => \N__14123\
        );

    \I__2822\ : Span4Mux_v
    port map (
            O => \N__14123\,
            I => \N__14119\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14122\,
            I => \N__14116\
        );

    \I__2820\ : Sp12to4
    port map (
            O => \N__14119\,
            I => \N__14111\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__14116\,
            I => \N__14111\
        );

    \I__2818\ : Span12Mux_h
    port map (
            O => \N__14111\,
            I => \N__14108\
        );

    \I__2817\ : Odrv12
    port map (
            O => \N__14108\,
            I => port_clk_c
        );

    \I__2816\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14101\
        );

    \I__2815\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14098\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14101\,
            I => \this_start_data_delay_this_edge_detector_M_last_q\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14098\,
            I => \this_start_data_delay_this_edge_detector_M_last_q\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14090\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__14090\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_0\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14084\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__14084\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_3\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14081\,
            I => \N__14078\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14078\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_1\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14075\,
            I => \N__14072\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14072\,
            I => \this_start_data_delay.this_delay.M_pipe_qZ0Z_2\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14069\,
            I => \N__14066\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__14066\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_5\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__14060\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_1\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14054\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14054\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_2\
        );

    \I__2798\ : InMux
    port map (
            O => \N__14051\,
            I => \N__14043\
        );

    \I__2797\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14043\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14039\
        );

    \I__2795\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14036\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__14043\,
            I => \N__14033\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14042\,
            I => \N__14030\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__14039\,
            I => \N__14025\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14036\,
            I => \N__14025\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__14033\,
            I => \N__14022\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14030\,
            I => \N__14017\
        );

    \I__2788\ : Span12Mux_v
    port map (
            O => \N__14025\,
            I => \N__14017\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__14022\,
            I => \this_vga_signals.un12_address_cry_2_c_RNIPIBB\
        );

    \I__2786\ : Odrv12
    port map (
            O => \N__14017\,
            I => \this_vga_signals.un12_address_cry_2_c_RNIPIBB\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__14009\,
            I => \N__14005\
        );

    \I__2783\ : InMux
    port map (
            O => \N__14008\,
            I => \N__14002\
        );

    \I__2782\ : Span12Mux_s10_h
    port map (
            O => \N__14005\,
            I => \N__13997\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14002\,
            I => \N__13997\
        );

    \I__2780\ : Span12Mux_h
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__2779\ : Odrv12
    port map (
            O => \N__13994\,
            I => \this_vga_signals.un12_address_cry_1_c_RNINFAB\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__13991\,
            I => \this_vga_signals.mult1_un96_sum_c5_0_1_0_1_cascade_\
        );

    \I__2777\ : InMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__13985\,
            I => \this_vga_signals.N_3_1_2\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__13979\,
            I => \this_vga_signals.g1_0_0_0_1\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__13976\,
            I => \this_vga_signals.mult1_un96_sum_c5_cascade_\
        );

    \I__2772\ : InMux
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__13967\,
            I => \this_vga_signals.g2_0\
        );

    \I__2769\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__13961\,
            I => \this_vga_signals.mult1_un96_sum_axbxc5_2\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__13958\,
            I => \this_vga_signals.g1_0_3_cascade_\
        );

    \I__2766\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__13952\,
            I => \this_vga_signals.mult1_un89_sum_c5_0_0_0_0\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__13949\,
            I => \N__13946\
        );

    \I__2763\ : CascadeBuf
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__2761\ : CascadeBuf
    port map (
            O => \N__13940\,
            I => \N__13937\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__2759\ : CascadeBuf
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__2757\ : CascadeBuf
    port map (
            O => \N__13928\,
            I => \N__13925\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__13925\,
            I => \N__13922\
        );

    \I__2755\ : CascadeBuf
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__2753\ : CascadeBuf
    port map (
            O => \N__13916\,
            I => \N__13913\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__13913\,
            I => \N__13910\
        );

    \I__2751\ : CascadeBuf
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__13907\,
            I => \N__13904\
        );

    \I__2749\ : CascadeBuf
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__2747\ : CascadeBuf
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2745\ : CascadeBuf
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__2743\ : CascadeBuf
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__2741\ : CascadeBuf
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__2739\ : CascadeBuf
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__2737\ : CascadeBuf
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__2735\ : CascadeBuf
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__2733\ : InMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__13853\,
            I => \N__13850\
        );

    \I__2731\ : Span12Mux_h
    port map (
            O => \N__13850\,
            I => \N__13847\
        );

    \I__2730\ : Span12Mux_v
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__2729\ : Odrv12
    port map (
            O => \N__13844\,
            I => \M_this_vga_signals_address_0\
        );

    \I__2728\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__13838\,
            I => \N__13835\
        );

    \I__2726\ : Span4Mux_h
    port map (
            O => \N__13835\,
            I => \N__13832\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__13832\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__2724\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13826\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__13826\,
            I => \this_vga_signals.if_N_3_2_i_1\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__13823\,
            I => \N__13810\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__13822\,
            I => \N__13807\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__13821\,
            I => \N__13803\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__13820\,
            I => \N__13799\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__13819\,
            I => \N__13795\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__13818\,
            I => \N__13792\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__13817\,
            I => \N__13789\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__13816\,
            I => \N__13786\
        );

    \I__2714\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13781\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__13814\,
            I => \N__13778\
        );

    \I__2712\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13766\
        );

    \I__2711\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13763\
        );

    \I__2710\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13757\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13806\,
            I => \N__13752\
        );

    \I__2708\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13752\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__13802\,
            I => \N__13749\
        );

    \I__2706\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13739\
        );

    \I__2705\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13739\
        );

    \I__2704\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13739\
        );

    \I__2703\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13739\
        );

    \I__2702\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13734\
        );

    \I__2701\ : InMux
    port map (
            O => \N__13786\,
            I => \N__13734\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__13785\,
            I => \N__13730\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__13784\,
            I => \N__13726\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__13781\,
            I => \N__13723\
        );

    \I__2697\ : InMux
    port map (
            O => \N__13778\,
            I => \N__13720\
        );

    \I__2696\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13717\
        );

    \I__2695\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13710\
        );

    \I__2694\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13710\
        );

    \I__2693\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13710\
        );

    \I__2692\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13706\
        );

    \I__2691\ : InMux
    port map (
            O => \N__13772\,
            I => \N__13703\
        );

    \I__2690\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13698\
        );

    \I__2689\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13698\
        );

    \I__2688\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13695\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__13766\,
            I => \N__13690\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__13763\,
            I => \N__13690\
        );

    \I__2685\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13687\
        );

    \I__2684\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13682\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13682\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__13757\,
            I => \N__13677\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__13752\,
            I => \N__13677\
        );

    \I__2680\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13674\
        );

    \I__2679\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13671\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__13739\,
            I => \N__13666\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__13734\,
            I => \N__13666\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13657\
        );

    \I__2675\ : InMux
    port map (
            O => \N__13730\,
            I => \N__13657\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13729\,
            I => \N__13657\
        );

    \I__2673\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13657\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__13723\,
            I => \N__13654\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__13720\,
            I => \N__13649\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__13717\,
            I => \N__13649\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__13710\,
            I => \N__13646\
        );

    \I__2668\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13643\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__13706\,
            I => \N__13640\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__13703\,
            I => \N__13633\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__13698\,
            I => \N__13633\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__13695\,
            I => \N__13633\
        );

    \I__2663\ : Span4Mux_v
    port map (
            O => \N__13690\,
            I => \N__13630\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__13687\,
            I => \N__13625\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__13682\,
            I => \N__13625\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__13677\,
            I => \N__13614\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__13674\,
            I => \N__13614\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__13671\,
            I => \N__13614\
        );

    \I__2657\ : Span4Mux_v
    port map (
            O => \N__13666\,
            I => \N__13614\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__13657\,
            I => \N__13614\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__13654\,
            I => \N__13611\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__13649\,
            I => \N__13604\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__13646\,
            I => \N__13604\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__13643\,
            I => \N__13604\
        );

    \I__2651\ : Span4Mux_h
    port map (
            O => \N__13640\,
            I => \N__13599\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__13633\,
            I => \N__13599\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__13630\,
            I => \N__13592\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__13625\,
            I => \N__13592\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__13614\,
            I => \N__13592\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__13611\,
            I => \this_vga_signals.un12_address_cry_4_c_RNITODB\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__13604\,
            I => \this_vga_signals.un12_address_cry_4_c_RNITODB\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__13599\,
            I => \this_vga_signals.un12_address_cry_4_c_RNITODB\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__13592\,
            I => \this_vga_signals.un12_address_cry_4_c_RNITODB\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13571\
        );

    \I__2640\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13566\
        );

    \I__2639\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13566\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__13577\,
            I => \N__13560\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__13576\,
            I => \N__13557\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13575\,
            I => \N__13549\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13574\,
            I => \N__13546\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__13571\,
            I => \N__13541\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__13566\,
            I => \N__13541\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13565\,
            I => \N__13532\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13532\
        );

    \I__2630\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13532\
        );

    \I__2629\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13532\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13529\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13524\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13524\
        );

    \I__2625\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13519\
        );

    \I__2624\ : InMux
    port map (
            O => \N__13553\,
            I => \N__13519\
        );

    \I__2623\ : InMux
    port map (
            O => \N__13552\,
            I => \N__13516\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13513\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__13546\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__13541\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__13532\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__13529\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__13524\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__13519\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__13516\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__13513\,
            I => \this_vga_signals.mult1_un75_sum_axbxc5\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13493\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__13493\,
            I => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_3\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \N__13483\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__13489\,
            I => \N__13479\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__13488\,
            I => \N__13475\
        );

    \I__2608\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13472\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13467\
        );

    \I__2606\ : InMux
    port map (
            O => \N__13483\,
            I => \N__13458\
        );

    \I__2605\ : InMux
    port map (
            O => \N__13482\,
            I => \N__13458\
        );

    \I__2604\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13455\
        );

    \I__2603\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13444\
        );

    \I__2602\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13441\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__13472\,
            I => \N__13438\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13471\,
            I => \N__13433\
        );

    \I__2599\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13433\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__13467\,
            I => \N__13430\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13425\
        );

    \I__2596\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13425\
        );

    \I__2595\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13422\
        );

    \I__2594\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13419\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__13458\,
            I => \N__13414\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__13455\,
            I => \N__13414\
        );

    \I__2591\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13409\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13453\,
            I => \N__13409\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__13452\,
            I => \N__13406\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__13451\,
            I => \N__13403\
        );

    \I__2587\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13396\
        );

    \I__2586\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13393\
        );

    \I__2585\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13390\
        );

    \I__2584\ : InMux
    port map (
            O => \N__13447\,
            I => \N__13387\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__13444\,
            I => \N__13378\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__13441\,
            I => \N__13378\
        );

    \I__2581\ : Span4Mux_v
    port map (
            O => \N__13438\,
            I => \N__13378\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__13433\,
            I => \N__13378\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__13430\,
            I => \N__13373\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__13425\,
            I => \N__13373\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__13422\,
            I => \N__13368\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13419\,
            I => \N__13368\
        );

    \I__2575\ : Span4Mux_v
    port map (
            O => \N__13414\,
            I => \N__13363\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__13409\,
            I => \N__13363\
        );

    \I__2573\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13360\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13403\,
            I => \N__13355\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13402\,
            I => \N__13355\
        );

    \I__2570\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13350\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13350\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13346\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__13396\,
            I => \N__13337\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__13393\,
            I => \N__13337\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13390\,
            I => \N__13337\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__13387\,
            I => \N__13337\
        );

    \I__2563\ : Span4Mux_h
    port map (
            O => \N__13378\,
            I => \N__13334\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__13373\,
            I => \N__13329\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__13368\,
            I => \N__13329\
        );

    \I__2560\ : Span4Mux_h
    port map (
            O => \N__13363\,
            I => \N__13324\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__13360\,
            I => \N__13324\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__13355\,
            I => \N__13319\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__13350\,
            I => \N__13319\
        );

    \I__2556\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13316\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__13346\,
            I => \this_vga_signals.un12_address_cry_5_c_RNIVREB\
        );

    \I__2554\ : Odrv12
    port map (
            O => \N__13337\,
            I => \this_vga_signals.un12_address_cry_5_c_RNIVREB\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__13334\,
            I => \this_vga_signals.un12_address_cry_5_c_RNIVREB\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__13329\,
            I => \this_vga_signals.un12_address_cry_5_c_RNIVREB\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__13324\,
            I => \this_vga_signals.un12_address_cry_5_c_RNIVREB\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__13319\,
            I => \this_vga_signals.un12_address_cry_5_c_RNIVREB\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__13316\,
            I => \this_vga_signals.un12_address_cry_5_c_RNIVREB\
        );

    \I__2548\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13295\
        );

    \I__2547\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13292\
        );

    \I__2546\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13289\
        );

    \I__2545\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13284\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__13295\,
            I => \N__13275\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__13292\,
            I => \N__13272\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__13289\,
            I => \N__13268\
        );

    \I__2541\ : InMux
    port map (
            O => \N__13288\,
            I => \N__13265\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13262\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__13284\,
            I => \N__13259\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13256\
        );

    \I__2537\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13253\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13250\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13245\
        );

    \I__2534\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13245\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13242\
        );

    \I__2532\ : Span4Mux_h
    port map (
            O => \N__13275\,
            I => \N__13237\
        );

    \I__2531\ : Span4Mux_h
    port map (
            O => \N__13272\,
            I => \N__13237\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13271\,
            I => \N__13234\
        );

    \I__2529\ : Odrv12
    port map (
            O => \N__13268\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13265\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13262\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__13259\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__13256\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__13253\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__13250\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__13245\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13242\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__13237\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13234\,
            I => this_vga_signals_un17_address_if_m2_2_0
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__13211\,
            I => \N__13207\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__13210\,
            I => \N__13204\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13207\,
            I => \N__13201\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13204\,
            I => \N__13198\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__13201\,
            I => \N__13193\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__13198\,
            I => \N__13193\
        );

    \I__2512\ : Odrv12
    port map (
            O => \N__13193\,
            I => \this_vga_signals.g0_38\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13190\,
            I => \N__13186\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13189\,
            I => \N__13183\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__13186\,
            I => \N__13180\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__13183\,
            I => \this_vga_signals.N_4_0_1\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__13180\,
            I => \this_vga_signals.N_4_0_1\
        );

    \I__2506\ : InMux
    port map (
            O => \N__13175\,
            I => \N__13172\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13172\,
            I => \this_vga_signals.if_N_3_2_i_2_0\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13166\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13166\,
            I => \this_start_address_delay.this_delay.M_pipe_qZ0Z_0\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13163\,
            I => \N__13160\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__13160\,
            I => \this_vga_signals.g1_0_0_0_0\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__13157\,
            I => \this_vga_signals.g0_0_3_cascade_\
        );

    \I__2499\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13151\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__13151\,
            I => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_4\
        );

    \I__2497\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__13145\,
            I => \this_vga_signals.g0_6\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13139\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__13139\,
            I => \this_vga_signals.g0_13\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13132\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13135\,
            I => \N__13129\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13132\,
            I => \this_vga_signals.if_N_3_2_i_0\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__13129\,
            I => \this_vga_signals.if_N_3_2_i_0\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__13121\,
            I => \N__13118\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__13118\,
            I => \this_vga_signals.g0_0_0_a2_1\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13112\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13112\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_0\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__13109\,
            I => \this_vga_signals.g1_2_cascade_\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__13106\,
            I => \this_vga_signals.r_N_2_0_0_2_cascade_\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13103\,
            I => \N__13100\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13100\,
            I => \this_vga_signals.N_3_1_1\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__13097\,
            I => \N__13094\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13091\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13091\,
            I => \N__13088\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__13088\,
            I => \this_vga_signals.g0_3_1\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13078\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13084\,
            I => \N__13073\
        );

    \I__2474\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13068\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13063\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13063\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13059\
        );

    \I__2470\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13054\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13054\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13051\
        );

    \I__2467\ : InMux
    port map (
            O => \N__13072\,
            I => \N__13046\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13071\,
            I => \N__13046\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13068\,
            I => \N__13036\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13063\,
            I => \N__13036\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13032\
        );

    \I__2462\ : Span4Mux_h
    port map (
            O => \N__13059\,
            I => \N__13027\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__13054\,
            I => \N__13027\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__13051\,
            I => \N__13022\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13046\,
            I => \N__13022\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13017\
        );

    \I__2457\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13017\
        );

    \I__2456\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13010\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13010\
        );

    \I__2454\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13010\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__13036\,
            I => \N__13007\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13035\,
            I => \N__13004\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__13032\,
            I => \this_vga_signals.mult1_un68_sum_c5\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__13027\,
            I => \this_vga_signals.mult1_un68_sum_c5\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__13022\,
            I => \this_vga_signals.mult1_un68_sum_c5\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__13017\,
            I => \this_vga_signals.mult1_un68_sum_c5\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__13010\,
            I => \this_vga_signals.mult1_un68_sum_c5\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__13007\,
            I => \this_vga_signals.mult1_un68_sum_c5\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__13004\,
            I => \this_vga_signals.mult1_un68_sum_c5\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__12989\,
            I => \N__12983\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__12988\,
            I => \N__12972\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__12987\,
            I => \N__12969\
        );

    \I__2441\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12964\
        );

    \I__2440\ : InMux
    port map (
            O => \N__12983\,
            I => \N__12964\
        );

    \I__2439\ : InMux
    port map (
            O => \N__12982\,
            I => \N__12961\
        );

    \I__2438\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12958\
        );

    \I__2437\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12954\
        );

    \I__2436\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12951\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__12978\,
            I => \N__12946\
        );

    \I__2434\ : InMux
    port map (
            O => \N__12977\,
            I => \N__12942\
        );

    \I__2433\ : InMux
    port map (
            O => \N__12976\,
            I => \N__12933\
        );

    \I__2432\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12933\
        );

    \I__2431\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12933\
        );

    \I__2430\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12933\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__12964\,
            I => \N__12930\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__12961\,
            I => \N__12925\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__12958\,
            I => \N__12925\
        );

    \I__2426\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12922\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__12954\,
            I => \N__12919\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__12951\,
            I => \N__12916\
        );

    \I__2423\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12913\
        );

    \I__2422\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12908\
        );

    \I__2421\ : InMux
    port map (
            O => \N__12946\,
            I => \N__12908\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__12945\,
            I => \N__12904\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__12942\,
            I => \N__12901\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__12933\,
            I => \N__12898\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__12930\,
            I => \N__12891\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__12925\,
            I => \N__12891\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__12922\,
            I => \N__12891\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__12919\,
            I => \N__12888\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__12916\,
            I => \N__12881\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__12913\,
            I => \N__12881\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__12908\,
            I => \N__12881\
        );

    \I__2410\ : InMux
    port map (
            O => \N__12907\,
            I => \N__12876\
        );

    \I__2409\ : InMux
    port map (
            O => \N__12904\,
            I => \N__12876\
        );

    \I__2408\ : Span4Mux_h
    port map (
            O => \N__12901\,
            I => \N__12873\
        );

    \I__2407\ : Span12Mux_v
    port map (
            O => \N__12898\,
            I => \N__12870\
        );

    \I__2406\ : Span4Mux_h
    port map (
            O => \N__12891\,
            I => \N__12867\
        );

    \I__2405\ : Span4Mux_h
    port map (
            O => \N__12888\,
            I => \N__12862\
        );

    \I__2404\ : Span4Mux_h
    port map (
            O => \N__12881\,
            I => \N__12862\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__12876\,
            I => \N__12859\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__12873\,
            I => \this_vga_signals.un12_address_cry_3_c_RNIRLCB\
        );

    \I__2401\ : Odrv12
    port map (
            O => \N__12870\,
            I => \this_vga_signals.un12_address_cry_3_c_RNIRLCB\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__12867\,
            I => \this_vga_signals.un12_address_cry_3_c_RNIRLCB\
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__12862\,
            I => \this_vga_signals.un12_address_cry_3_c_RNIRLCB\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__12859\,
            I => \this_vga_signals.un12_address_cry_3_c_RNIRLCB\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__12848\,
            I => \this_vga_signals.g0_5_3_cascade_\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__12845\,
            I => \this_vga_signals.g0_3_0_a2_1_cascade_\
        );

    \I__2395\ : InMux
    port map (
            O => \N__12842\,
            I => \N__12839\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__12839\,
            I => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_2\
        );

    \I__2393\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12829\
        );

    \I__2391\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12826\
        );

    \I__2390\ : Span4Mux_h
    port map (
            O => \N__12829\,
            I => \N__12823\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__12826\,
            I => \N__12820\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__12823\,
            I => \this_vga_signals.if_N_8_mux_2_0\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__12820\,
            I => \this_vga_signals.if_N_8_mux_2_0\
        );

    \I__2386\ : InMux
    port map (
            O => \N__12815\,
            I => \N__12809\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__12814\,
            I => \N__12791\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__12813\,
            I => \N__12787\
        );

    \I__2383\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12783\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__12809\,
            I => \N__12780\
        );

    \I__2381\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12775\
        );

    \I__2380\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12775\
        );

    \I__2379\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12772\
        );

    \I__2378\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12767\
        );

    \I__2377\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12767\
        );

    \I__2376\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12760\
        );

    \I__2375\ : InMux
    port map (
            O => \N__12802\,
            I => \N__12760\
        );

    \I__2374\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12760\
        );

    \I__2373\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12751\
        );

    \I__2372\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12751\
        );

    \I__2371\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12751\
        );

    \I__2370\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12751\
        );

    \I__2369\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12744\
        );

    \I__2368\ : InMux
    port map (
            O => \N__12795\,
            I => \N__12744\
        );

    \I__2367\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12744\
        );

    \I__2366\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12741\
        );

    \I__2365\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12734\
        );

    \I__2364\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12734\
        );

    \I__2363\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12734\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__12783\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__12780\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12775\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__12772\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__12767\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__12760\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__12751\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__12744\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__12741\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__12734\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5
        );

    \I__2352\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12707\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12704\
        );

    \I__2350\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12701\
        );

    \I__2349\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12698\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__12707\,
            I => \this_vga_signals.if_N_3_2_i\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__12704\,
            I => \this_vga_signals.if_N_3_2_i\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__12701\,
            I => \this_vga_signals.if_N_3_2_i\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__12698\,
            I => \this_vga_signals.if_N_3_2_i\
        );

    \I__2344\ : InMux
    port map (
            O => \N__12689\,
            I => \N__12686\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__12686\,
            I => \N__12683\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__12683\,
            I => \N__12680\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__12680\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__12677\,
            I => \N__12668\
        );

    \I__2339\ : InMux
    port map (
            O => \N__12676\,
            I => \N__12664\
        );

    \I__2338\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12656\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__12674\,
            I => \N__12653\
        );

    \I__2336\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12643\
        );

    \I__2335\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12643\
        );

    \I__2334\ : InMux
    port map (
            O => \N__12671\,
            I => \N__12643\
        );

    \I__2333\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12638\
        );

    \I__2332\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12638\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__12664\,
            I => \N__12634\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12629\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12662\,
            I => \N__12629\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__12661\,
            I => \N__12621\
        );

    \I__2327\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12615\
        );

    \I__2326\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12615\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__12656\,
            I => \N__12612\
        );

    \I__2324\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12607\
        );

    \I__2323\ : InMux
    port map (
            O => \N__12652\,
            I => \N__12607\
        );

    \I__2322\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12604\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__12650\,
            I => \N__12596\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__12643\,
            I => \N__12593\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__12638\,
            I => \N__12590\
        );

    \I__2318\ : InMux
    port map (
            O => \N__12637\,
            I => \N__12586\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__12634\,
            I => \N__12581\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__12629\,
            I => \N__12581\
        );

    \I__2315\ : InMux
    port map (
            O => \N__12628\,
            I => \N__12578\
        );

    \I__2314\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12569\
        );

    \I__2313\ : InMux
    port map (
            O => \N__12626\,
            I => \N__12569\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12569\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12624\,
            I => \N__12569\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12564\
        );

    \I__2309\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12564\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12615\,
            I => \N__12561\
        );

    \I__2307\ : Span4Mux_h
    port map (
            O => \N__12612\,
            I => \N__12554\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__12607\,
            I => \N__12554\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__12604\,
            I => \N__12554\
        );

    \I__2304\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12547\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12602\,
            I => \N__12547\
        );

    \I__2302\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12547\
        );

    \I__2301\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12540\
        );

    \I__2300\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12540\
        );

    \I__2299\ : InMux
    port map (
            O => \N__12596\,
            I => \N__12540\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__12593\,
            I => \N__12535\
        );

    \I__2297\ : Span4Mux_h
    port map (
            O => \N__12590\,
            I => \N__12535\
        );

    \I__2296\ : InMux
    port map (
            O => \N__12589\,
            I => \N__12532\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__12586\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__12581\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__12578\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__12569\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__12564\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__12561\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__12554\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12547\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__12540\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__12535\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__12532\,
            I => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2284\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__12506\,
            I => \N__12503\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__12503\,
            I => \this_vga_signals.g0_6_0\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__12500\,
            I => \this_vga_signals.g1_2_0_cascade_\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12494\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__12494\,
            I => \N__12491\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__12491\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__12488\,
            I => \this_vga_signals.g1_5_cascade_\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12478\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12484\,
            I => \N__12473\
        );

    \I__2274\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12473\
        );

    \I__2273\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12470\
        );

    \I__2272\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12467\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__12478\,
            I => \N__12462\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__12473\,
            I => \N__12459\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__12470\,
            I => \N__12456\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__12467\,
            I => \N__12453\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12448\
        );

    \I__2266\ : InMux
    port map (
            O => \N__12465\,
            I => \N__12448\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__12462\,
            I => \N__12437\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__12459\,
            I => \N__12437\
        );

    \I__2263\ : Span4Mux_h
    port map (
            O => \N__12456\,
            I => \N__12437\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__12453\,
            I => \N__12437\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12448\,
            I => \N__12437\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__12437\,
            I => \this_vga_signals.mult1_un75_sum_axb3\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12431\,
            I => \N__12428\
        );

    \I__2257\ : Odrv12
    port map (
            O => \N__12428\,
            I => \this_vga_signals.g0_0_1_1\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__12425\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_2_cascade_\
        );

    \I__2255\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12419\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__12419\,
            I => \this_vga_signals.g0_3\
        );

    \I__2253\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__12413\,
            I => \this_vga_signals.N_20_i_i_0\
        );

    \I__2251\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__12404\,
            I => \this_vga_signals.g0_0_a3_3\
        );

    \I__2248\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12397\
        );

    \I__2247\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12394\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12397\,
            I => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_0\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12394\,
            I => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_0\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__12389\,
            I => \this_vga_signals.N_11_cascade_\
        );

    \I__2243\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12383\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__12383\,
            I => \this_vga_signals.g0_0_a3_2\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__12380\,
            I => \this_vga_signals.g0_0_a3_5_cascade_\
        );

    \I__2240\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12374\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__12374\,
            I => \this_vga_signals.g0_i_x4_4_a3\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12368\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__12368\,
            I => \this_vga_signals.N_3_3_0\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12362\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__12362\,
            I => \N__12359\
        );

    \I__2234\ : Odrv12
    port map (
            O => \N__12359\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_1\
        );

    \I__2233\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12353\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__12353\,
            I => \this_vga_signals.g0_0_1_0\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__12350\,
            I => \this_vga_signals.g1_5_0_0_cascade_\
        );

    \I__2230\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12344\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__12344\,
            I => \this_vga_signals.r_N_2_0_0_0\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__12341\,
            I => \N__12338\
        );

    \I__2227\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12335\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__12335\,
            I => \N__12332\
        );

    \I__2225\ : Span4Mux_h
    port map (
            O => \N__12332\,
            I => \N__12329\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__12329\,
            I => \this_vga_signals.g0_1_0\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__12326\,
            I => \this_vga_signals.g0_1_2_cascade_\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12320\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__12320\,
            I => \N__12310\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12319\,
            I => \N__12303\
        );

    \I__2219\ : InMux
    port map (
            O => \N__12318\,
            I => \N__12303\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12295\
        );

    \I__2217\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12292\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12289\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12284\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12284\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__12310\,
            I => \N__12281\
        );

    \I__2212\ : InMux
    port map (
            O => \N__12309\,
            I => \N__12276\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12308\,
            I => \N__12276\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12273\
        );

    \I__2209\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12266\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12301\,
            I => \N__12266\
        );

    \I__2207\ : InMux
    port map (
            O => \N__12300\,
            I => \N__12266\
        );

    \I__2206\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12261\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12261\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12295\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12292\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__12289\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__12284\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__12281\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__12276\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__12273\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__12266\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__12261\,
            I => \this_vga_signals_un17_address_if_N_8_mux\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__12239\,
            I => \N__12236\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__12236\,
            I => \N__12233\
        );

    \I__2192\ : Span4Mux_v
    port map (
            O => \N__12233\,
            I => \N__12228\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12232\,
            I => \N__12223\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12223\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__12228\,
            I => \this_vga_signals.mult1_un54_sum_ac0_8\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__12223\,
            I => \this_vga_signals.mult1_un54_sum_ac0_8\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__2186\ : CascadeBuf
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__2184\ : CascadeBuf
    port map (
            O => \N__12209\,
            I => \N__12206\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__2182\ : CascadeBuf
    port map (
            O => \N__12203\,
            I => \N__12200\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__12200\,
            I => \N__12197\
        );

    \I__2180\ : CascadeBuf
    port map (
            O => \N__12197\,
            I => \N__12194\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__2178\ : CascadeBuf
    port map (
            O => \N__12191\,
            I => \N__12188\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \N__12185\
        );

    \I__2176\ : CascadeBuf
    port map (
            O => \N__12185\,
            I => \N__12182\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__12182\,
            I => \N__12179\
        );

    \I__2174\ : CascadeBuf
    port map (
            O => \N__12179\,
            I => \N__12176\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__12176\,
            I => \N__12173\
        );

    \I__2172\ : CascadeBuf
    port map (
            O => \N__12173\,
            I => \N__12170\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__12170\,
            I => \N__12167\
        );

    \I__2170\ : CascadeBuf
    port map (
            O => \N__12167\,
            I => \N__12164\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__12164\,
            I => \N__12161\
        );

    \I__2168\ : CascadeBuf
    port map (
            O => \N__12161\,
            I => \N__12158\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__12158\,
            I => \N__12155\
        );

    \I__2166\ : CascadeBuf
    port map (
            O => \N__12155\,
            I => \N__12152\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__12152\,
            I => \N__12149\
        );

    \I__2164\ : CascadeBuf
    port map (
            O => \N__12149\,
            I => \N__12146\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__12146\,
            I => \N__12143\
        );

    \I__2162\ : CascadeBuf
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__12140\,
            I => \N__12137\
        );

    \I__2160\ : CascadeBuf
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__12134\,
            I => \N__12131\
        );

    \I__2158\ : CascadeBuf
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12125\,
            I => \N__12122\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__12122\,
            I => \N__12119\
        );

    \I__2154\ : Sp12to4
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__2153\ : Span12Mux_s11_v
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__2152\ : Span12Mux_h
    port map (
            O => \N__12113\,
            I => \N__12110\
        );

    \I__2151\ : Odrv12
    port map (
            O => \N__12110\,
            I => \M_this_vga_signals_address_6\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12104\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__12104\,
            I => \this_vga_signals.N_4\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__12101\,
            I => \this_vram.M_this_vram_read_data_1_cascade_\
        );

    \I__2147\ : IoInMux
    port map (
            O => \N__12098\,
            I => \N__12095\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__2145\ : IoSpan4Mux
    port map (
            O => \N__12092\,
            I => \N__12089\
        );

    \I__2144\ : IoSpan4Mux
    port map (
            O => \N__12089\,
            I => \N__12085\
        );

    \I__2143\ : IoInMux
    port map (
            O => \N__12088\,
            I => \N__12082\
        );

    \I__2142\ : Sp12to4
    port map (
            O => \N__12085\,
            I => \N__12077\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__12082\,
            I => \N__12077\
        );

    \I__2140\ : Span12Mux_s6_h
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__2139\ : Odrv12
    port map (
            O => \N__12074\,
            I => rgb_c_2
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__12071\,
            I => \N__12068\
        );

    \I__2137\ : InMux
    port map (
            O => \N__12068\,
            I => \N__12065\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__12062\,
            I => \this_vga_signals.g0_4\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12056\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__12053\,
            I => \this_vga_signals.if_N_8_mux_2_2_1\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__12050\,
            I => \this_vga_signals.N_3_1_0_1_cascade_\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12044\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12044\,
            I => \this_vga_signals.g1_2_0_0\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12038\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12038\,
            I => \this_vga_signals.g0_0_0_0\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__12035\,
            I => \N__12026\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__12034\,
            I => \N__12018\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12014\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12032\,
            I => \N__12009\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12031\,
            I => \N__12004\
        );

    \I__2121\ : InMux
    port map (
            O => \N__12030\,
            I => \N__12004\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__12029\,
            I => \N__12001\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12026\,
            I => \N__11997\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__12025\,
            I => \N__11990\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12024\,
            I => \N__11986\
        );

    \I__2116\ : InMux
    port map (
            O => \N__12023\,
            I => \N__11983\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12022\,
            I => \N__11978\
        );

    \I__2114\ : InMux
    port map (
            O => \N__12021\,
            I => \N__11978\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12018\,
            I => \N__11973\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12017\,
            I => \N__11973\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12014\,
            I => \N__11970\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12013\,
            I => \N__11965\
        );

    \I__2109\ : InMux
    port map (
            O => \N__12012\,
            I => \N__11965\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__12009\,
            I => \N__11960\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__12004\,
            I => \N__11960\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12001\,
            I => \N__11955\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12000\,
            I => \N__11955\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__11997\,
            I => \N__11950\
        );

    \I__2103\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11943\
        );

    \I__2102\ : InMux
    port map (
            O => \N__11995\,
            I => \N__11943\
        );

    \I__2101\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11943\
        );

    \I__2100\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11940\
        );

    \I__2099\ : InMux
    port map (
            O => \N__11990\,
            I => \N__11935\
        );

    \I__2098\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11935\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__11986\,
            I => \N__11930\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__11983\,
            I => \N__11930\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__11978\,
            I => \N__11925\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__11973\,
            I => \N__11925\
        );

    \I__2093\ : Span4Mux_h
    port map (
            O => \N__11970\,
            I => \N__11916\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__11965\,
            I => \N__11916\
        );

    \I__2091\ : Span4Mux_v
    port map (
            O => \N__11960\,
            I => \N__11916\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__11955\,
            I => \N__11916\
        );

    \I__2089\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11913\
        );

    \I__2088\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11910\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__11950\,
            I => \N__11901\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__11943\,
            I => \N__11901\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__11940\,
            I => \N__11901\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__11935\,
            I => \N__11901\
        );

    \I__2083\ : Span4Mux_h
    port map (
            O => \N__11930\,
            I => \N__11896\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__11925\,
            I => \N__11896\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__11916\,
            I => \N__11893\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__11913\,
            I => \this_vga_signals.if_m1_0_0\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__11910\,
            I => \this_vga_signals.if_m1_0_0\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__11901\,
            I => \this_vga_signals.if_m1_0_0\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__11896\,
            I => \this_vga_signals.if_m1_0_0\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__11893\,
            I => \this_vga_signals.if_m1_0_0\
        );

    \I__2075\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11878\
        );

    \I__2074\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11875\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__11878\,
            I => \this_vga_signals.N_21\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__11875\,
            I => \this_vga_signals.N_21\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__11870\,
            I => \N__11866\
        );

    \I__2070\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11861\
        );

    \I__2069\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11856\
        );

    \I__2068\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11856\
        );

    \I__2067\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11853\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__11861\,
            I => \N__11848\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__11856\,
            I => \N__11841\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__11853\,
            I => \N__11828\
        );

    \I__2063\ : InMux
    port map (
            O => \N__11852\,
            I => \N__11823\
        );

    \I__2062\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11823\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__11848\,
            I => \N__11820\
        );

    \I__2060\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11817\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11810\
        );

    \I__2058\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11810\
        );

    \I__2057\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11810\
        );

    \I__2056\ : Span4Mux_h
    port map (
            O => \N__11841\,
            I => \N__11807\
        );

    \I__2055\ : InMux
    port map (
            O => \N__11840\,
            I => \N__11802\
        );

    \I__2054\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11802\
        );

    \I__2053\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11795\
        );

    \I__2052\ : InMux
    port map (
            O => \N__11837\,
            I => \N__11795\
        );

    \I__2051\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11795\
        );

    \I__2050\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11792\
        );

    \I__2049\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11783\
        );

    \I__2048\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11783\
        );

    \I__2047\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11783\
        );

    \I__2046\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11783\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__11828\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__11823\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__11820\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__11817\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__11810\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__11807\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__11802\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__11795\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__11792\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__11783\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__11762\,
            I => \N__11757\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__11761\,
            I => \N__11752\
        );

    \I__2033\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11749\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11744\
        );

    \I__2031\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11735\
        );

    \I__2030\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11735\
        );

    \I__2029\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11735\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__11749\,
            I => \N__11732\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__11748\,
            I => \N__11729\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__11747\,
            I => \N__11725\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__11744\,
            I => \N__11719\
        );

    \I__2024\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11714\
        );

    \I__2023\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11714\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__11735\,
            I => \N__11711\
        );

    \I__2021\ : Span4Mux_h
    port map (
            O => \N__11732\,
            I => \N__11708\
        );

    \I__2020\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11701\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11701\
        );

    \I__2018\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11701\
        );

    \I__2017\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11698\
        );

    \I__2016\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11693\
        );

    \I__2015\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11693\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__11719\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__11714\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__11711\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__11708\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__11701\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__11698\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__11693\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5\
        );

    \I__2007\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11673\
        );

    \I__2006\ : InMux
    port map (
            O => \N__11677\,
            I => \N__11670\
        );

    \I__2005\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11667\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__11673\,
            I => \this_vga_signals.N_12\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__11670\,
            I => \this_vga_signals.N_12\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__11667\,
            I => \this_vga_signals.N_12\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__11660\,
            I => \this_vga_signals.g0_0_0_a2_1_0_cascade_\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__11657\,
            I => \this_vga_signals.if_N_3_2_i_3_1_cascade_\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__1998\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__11648\,
            I => \this_vga_signals.N_31\
        );

    \I__1996\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__11642\,
            I => \this_vga_signals.N_20_i_i\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__11639\,
            I => \this_vga_signals.N_20_i_i_cascade_\
        );

    \I__1993\ : InMux
    port map (
            O => \N__11636\,
            I => \N__11633\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__11633\,
            I => \N__11630\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__11630\,
            I => \this_vga_signals.N_26_i_i\
        );

    \I__1990\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__11624\,
            I => \N__11619\
        );

    \I__1988\ : InMux
    port map (
            O => \N__11623\,
            I => \N__11616\
        );

    \I__1987\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11608\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__11619\,
            I => \N__11603\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__11616\,
            I => \N__11603\
        );

    \I__1984\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11600\
        );

    \I__1983\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11595\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11613\,
            I => \N__11595\
        );

    \I__1981\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11592\
        );

    \I__1980\ : InMux
    port map (
            O => \N__11611\,
            I => \N__11589\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__11608\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__11603\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__11600\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__11595\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__11592\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__11589\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1973\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11573\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__11573\,
            I => \N__11569\
        );

    \I__1971\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11566\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__11569\,
            I => \N__11557\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__11566\,
            I => \N__11557\
        );

    \I__1968\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11554\
        );

    \I__1967\ : InMux
    port map (
            O => \N__11564\,
            I => \N__11547\
        );

    \I__1966\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11547\
        );

    \I__1965\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11547\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__11557\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__11554\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__11547\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_1\
        );

    \I__1961\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11536\
        );

    \I__1960\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11533\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__11536\,
            I => \N__11530\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__11533\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__11530\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1956\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11521\
        );

    \I__1955\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11518\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__11521\,
            I => \N__11515\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__11518\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__11515\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__11510\,
            I => \N__11507\
        );

    \I__1950\ : CascadeBuf
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__1948\ : CascadeBuf
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__1946\ : CascadeBuf
    port map (
            O => \N__11495\,
            I => \N__11492\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__11492\,
            I => \N__11489\
        );

    \I__1944\ : CascadeBuf
    port map (
            O => \N__11489\,
            I => \N__11486\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__11486\,
            I => \N__11483\
        );

    \I__1942\ : CascadeBuf
    port map (
            O => \N__11483\,
            I => \N__11480\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__1940\ : CascadeBuf
    port map (
            O => \N__11477\,
            I => \N__11474\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__11474\,
            I => \N__11471\
        );

    \I__1938\ : CascadeBuf
    port map (
            O => \N__11471\,
            I => \N__11468\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__11468\,
            I => \N__11465\
        );

    \I__1936\ : CascadeBuf
    port map (
            O => \N__11465\,
            I => \N__11462\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__11462\,
            I => \N__11459\
        );

    \I__1934\ : CascadeBuf
    port map (
            O => \N__11459\,
            I => \N__11456\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__11456\,
            I => \N__11453\
        );

    \I__1932\ : CascadeBuf
    port map (
            O => \N__11453\,
            I => \N__11450\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__11450\,
            I => \N__11447\
        );

    \I__1930\ : CascadeBuf
    port map (
            O => \N__11447\,
            I => \N__11444\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__11444\,
            I => \N__11441\
        );

    \I__1928\ : CascadeBuf
    port map (
            O => \N__11441\,
            I => \N__11438\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__11438\,
            I => \N__11435\
        );

    \I__1926\ : CascadeBuf
    port map (
            O => \N__11435\,
            I => \N__11432\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__11432\,
            I => \N__11429\
        );

    \I__1924\ : CascadeBuf
    port map (
            O => \N__11429\,
            I => \N__11426\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__11426\,
            I => \N__11423\
        );

    \I__1922\ : CascadeBuf
    port map (
            O => \N__11423\,
            I => \N__11420\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__11420\,
            I => \N__11417\
        );

    \I__1920\ : InMux
    port map (
            O => \N__11417\,
            I => \N__11414\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__11414\,
            I => \N__11411\
        );

    \I__1918\ : Span12Mux_h
    port map (
            O => \N__11411\,
            I => \N__11408\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__11408\,
            I => \M_this_vga_signals_address_9\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11402\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11402\,
            I => \N__11398\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11401\,
            I => \N__11395\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__11398\,
            I => \N__11390\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__11395\,
            I => \N__11387\
        );

    \I__1911\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11382\
        );

    \I__1910\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11382\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__11390\,
            I => \this_vga_signals.mult1_un54_sum_ac0_7\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__11387\,
            I => \this_vga_signals.mult1_un54_sum_ac0_7\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11382\,
            I => \this_vga_signals.mult1_un54_sum_ac0_7\
        );

    \I__1906\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11372\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__11372\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_4\
        );

    \I__1904\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__11366\,
            I => \this_vga_signals.g0_i_x4_4_a3_1\
        );

    \I__1902\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__11357\,
            I => \this_vga_signals.if_m1_0\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11351\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__11351\,
            I => \this_vga_signals.if_N_3_3_i\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__11348\,
            I => \this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5_cascade_\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__11345\,
            I => \this_vga_signals.if_N_3_2_i_cascade_\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__1894\ : CascadeBuf
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__11336\,
            I => \N__11333\
        );

    \I__1892\ : CascadeBuf
    port map (
            O => \N__11333\,
            I => \N__11330\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__11330\,
            I => \N__11327\
        );

    \I__1890\ : CascadeBuf
    port map (
            O => \N__11327\,
            I => \N__11324\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__11324\,
            I => \N__11321\
        );

    \I__1888\ : CascadeBuf
    port map (
            O => \N__11321\,
            I => \N__11318\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__11318\,
            I => \N__11315\
        );

    \I__1886\ : CascadeBuf
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__11312\,
            I => \N__11309\
        );

    \I__1884\ : CascadeBuf
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__11306\,
            I => \N__11303\
        );

    \I__1882\ : CascadeBuf
    port map (
            O => \N__11303\,
            I => \N__11300\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__11300\,
            I => \N__11297\
        );

    \I__1880\ : CascadeBuf
    port map (
            O => \N__11297\,
            I => \N__11294\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__11294\,
            I => \N__11291\
        );

    \I__1878\ : CascadeBuf
    port map (
            O => \N__11291\,
            I => \N__11288\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__1876\ : CascadeBuf
    port map (
            O => \N__11285\,
            I => \N__11282\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \N__11279\
        );

    \I__1874\ : CascadeBuf
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__1872\ : CascadeBuf
    port map (
            O => \N__11273\,
            I => \N__11270\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__11270\,
            I => \N__11267\
        );

    \I__1870\ : CascadeBuf
    port map (
            O => \N__11267\,
            I => \N__11264\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__11264\,
            I => \N__11261\
        );

    \I__1868\ : CascadeBuf
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__11258\,
            I => \N__11255\
        );

    \I__1866\ : CascadeBuf
    port map (
            O => \N__11255\,
            I => \N__11252\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__1864\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11243\
        );

    \I__1862\ : Span12Mux_s9_h
    port map (
            O => \N__11243\,
            I => \N__11240\
        );

    \I__1861\ : Span12Mux_v
    port map (
            O => \N__11240\,
            I => \N__11237\
        );

    \I__1860\ : Odrv12
    port map (
            O => \N__11237\,
            I => \M_this_vga_signals_address_3\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__11234\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_3L3_cascade_\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11228\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__11228\,
            I => \N__11225\
        );

    \I__1856\ : Span4Mux_v
    port map (
            O => \N__11225\,
            I => \N__11222\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__11222\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_2L1\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__11219\,
            I => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5_cascade_\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11213\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__11213\,
            I => \this_vga_signals.N_21_0\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11204\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__11201\,
            I => \this_vga_signals.g0_6_0_0_2\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__11195\,
            I => \this_vga_signals.if_N_8_mux_2_2\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__11192\,
            I => \this_vga_signals.mult1_un82_sum_axb3_cascade_\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__11189\,
            I => \this_vga_signals.address_i2_mux_cascade_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__11186\,
            I => \N__11183\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__11183\,
            I => \this_vga_signals.address_N_11\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11180\,
            I => \N__11177\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__11177\,
            I => \this_vga_signals.address_i2_mux_0\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__11174\,
            I => \this_vga_signals.address_m21_ns_1_cascade_\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11168\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__11168\,
            I => \this_vga_signals.address_i2_mux_1\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__11165\,
            I => \this_vga_signals.address_N_22_cascade_\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11159\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11159\,
            I => \this_vga_signals.address_N_36\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1832\ : CascadeBuf
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__11150\,
            I => \N__11147\
        );

    \I__1830\ : CascadeBuf
    port map (
            O => \N__11147\,
            I => \N__11144\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__11144\,
            I => \N__11141\
        );

    \I__1828\ : CascadeBuf
    port map (
            O => \N__11141\,
            I => \N__11138\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__11138\,
            I => \N__11135\
        );

    \I__1826\ : CascadeBuf
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__1824\ : CascadeBuf
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__1822\ : CascadeBuf
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__1820\ : CascadeBuf
    port map (
            O => \N__11117\,
            I => \N__11114\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__11114\,
            I => \N__11111\
        );

    \I__1818\ : CascadeBuf
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__1816\ : CascadeBuf
    port map (
            O => \N__11105\,
            I => \N__11102\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__1814\ : CascadeBuf
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__11096\,
            I => \N__11093\
        );

    \I__1812\ : CascadeBuf
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1810\ : CascadeBuf
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1808\ : CascadeBuf
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__1806\ : CascadeBuf
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__1804\ : CascadeBuf
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__1800\ : Sp12to4
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__1799\ : Span12Mux_s9_v
    port map (
            O => \N__11054\,
            I => \N__11051\
        );

    \I__1798\ : Odrv12
    port map (
            O => \N__11051\,
            I => \M_this_vga_signals_address_7\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11043\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11047\,
            I => \N__11038\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11038\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__11043\,
            I => \N__11035\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__11038\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__11035\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11020\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11017\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11011\
        );

    \I__1788\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11011\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11026\,
            I => \N__11008\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11005\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__11024\,
            I => \N__10999\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11023\,
            I => \N__10994\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11020\,
            I => \N__10987\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11017\,
            I => \N__10987\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__11016\,
            I => \N__10983\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11011\,
            I => \N__10978\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__11008\,
            I => \N__10978\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11005\,
            I => \N__10975\
        );

    \I__1777\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10972\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10969\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10966\
        );

    \I__1774\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10959\
        );

    \I__1773\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10959\
        );

    \I__1772\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10959\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__10994\,
            I => \N__10956\
        );

    \I__1770\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10951\
        );

    \I__1769\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10951\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__10987\,
            I => \N__10948\
        );

    \I__1767\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10943\
        );

    \I__1766\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10943\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__10978\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__10975\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__10972\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__10969\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__10966\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__10959\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__10956\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__10951\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__10948\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__10943\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1755\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10918\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__10921\,
            I => \N__10914\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__10918\,
            I => \N__10910\
        );

    \I__1752\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10905\
        );

    \I__1751\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10905\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__10913\,
            I => \N__10900\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__10910\,
            I => \N__10895\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__10905\,
            I => \N__10895\
        );

    \I__1747\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10890\
        );

    \I__1746\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10890\
        );

    \I__1745\ : InMux
    port map (
            O => \N__10900\,
            I => \N__10887\
        );

    \I__1744\ : Span4Mux_h
    port map (
            O => \N__10895\,
            I => \N__10884\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__10890\,
            I => \N__10881\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10887\,
            I => \N__10878\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__10884\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__10881\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__10878\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__10871\,
            I => \N__10865\
        );

    \I__1737\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10857\
        );

    \I__1736\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10857\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10857\
        );

    \I__1734\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10853\
        );

    \I__1733\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10850\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__10857\,
            I => \N__10847\
        );

    \I__1731\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10844\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__10853\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_0\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__10850\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_0\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__10847\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_0\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__10844\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__10832\,
            I => \this_vga_signals.if_m16_0_o4\
        );

    \I__1724\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10824\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10818\
        );

    \I__1722\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10815\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__10824\,
            I => \N__10810\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10807\
        );

    \I__1719\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10804\
        );

    \I__1718\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10801\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__10818\,
            I => \N__10798\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__10815\,
            I => \N__10795\
        );

    \I__1715\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10792\
        );

    \I__1714\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10787\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__10810\,
            I => \N__10784\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__10807\,
            I => \N__10781\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__10804\,
            I => \N__10772\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__10801\,
            I => \N__10772\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__10798\,
            I => \N__10772\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__10795\,
            I => \N__10772\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10769\
        );

    \I__1706\ : InMux
    port map (
            O => \N__10791\,
            I => \N__10766\
        );

    \I__1705\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10763\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__10787\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__10784\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__10781\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__10772\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__10769\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__10766\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__10763\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__10748\,
            I => \N__10736\
        );

    \I__1696\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10726\
        );

    \I__1695\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10726\
        );

    \I__1694\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10723\
        );

    \I__1693\ : InMux
    port map (
            O => \N__10744\,
            I => \N__10720\
        );

    \I__1692\ : InMux
    port map (
            O => \N__10743\,
            I => \N__10715\
        );

    \I__1691\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10715\
        );

    \I__1690\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10712\
        );

    \I__1689\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10709\
        );

    \I__1688\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10704\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10704\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__10735\,
            I => \N__10701\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10697\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10694\
        );

    \I__1683\ : InMux
    port map (
            O => \N__10732\,
            I => \N__10689\
        );

    \I__1682\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10689\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__10726\,
            I => \N__10684\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__10723\,
            I => \N__10684\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__10720\,
            I => \N__10673\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__10715\,
            I => \N__10673\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__10712\,
            I => \N__10673\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10673\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10673\
        );

    \I__1674\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10670\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \N__10661\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__10697\,
            I => \N__10648\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__10694\,
            I => \N__10648\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__10689\,
            I => \N__10648\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__10684\,
            I => \N__10648\
        );

    \I__1668\ : Span4Mux_v
    port map (
            O => \N__10673\,
            I => \N__10648\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__10670\,
            I => \N__10648\
        );

    \I__1666\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10645\
        );

    \I__1665\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10638\
        );

    \I__1664\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10638\
        );

    \I__1663\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10638\
        );

    \I__1662\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10633\
        );

    \I__1661\ : InMux
    port map (
            O => \N__10664\,
            I => \N__10633\
        );

    \I__1660\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10630\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__10648\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__10645\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__10638\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__10633\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__10630\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1654\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__10616\,
            I => \N__10612\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10609\
        );

    \I__1651\ : Odrv4
    port map (
            O => \N__10612\,
            I => \this_vga_signals.address_N_40\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10609\,
            I => \this_vga_signals.address_N_40\
        );

    \I__1649\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__10598\,
            I => \this_vga_signals.if_m4_0_1_0_0\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__10595\,
            I => \N_11_0_cascade_\
        );

    \I__1645\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10586\
        );

    \I__1644\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10586\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__10586\,
            I => \this_vga_signals.N_5_i\
        );

    \I__1642\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10580\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__10580\,
            I => \this_vga_signals.G_12_0_1\
        );

    \I__1640\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__10574\,
            I => \this_vga_signals.N_25\
        );

    \I__1638\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10562\
        );

    \I__1637\ : InMux
    port map (
            O => \N__10570\,
            I => \N__10562\
        );

    \I__1636\ : InMux
    port map (
            O => \N__10569\,
            I => \N__10557\
        );

    \I__1635\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10557\
        );

    \I__1634\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10554\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__10562\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__10557\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__10554\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__1630\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10540\
        );

    \I__1629\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__10545\,
            I => \N__10535\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__10540\,
            I => \N__10532\
        );

    \I__1626\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10528\
        );

    \I__1625\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10523\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10523\
        );

    \I__1623\ : Span4Mux_h
    port map (
            O => \N__10532\,
            I => \N__10514\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10511\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__10528\,
            I => \N__10508\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__10523\,
            I => \N__10505\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10522\,
            I => \N__10502\
        );

    \I__1618\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10499\
        );

    \I__1617\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10494\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10494\
        );

    \I__1615\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10491\
        );

    \I__1614\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10488\
        );

    \I__1613\ : Odrv4
    port map (
            O => \N__10514\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__10511\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__10508\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__10505\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__10502\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__10499\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__10494\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10491\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10488\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__10466\,
            I => \this_vga_signals.N_275\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__10463\,
            I => \this_vga_signals.if_N_9_i_i_cascade_\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__10457\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__10454\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__1597\ : CascadeBuf
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1595\ : CascadeBuf
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__1593\ : CascadeBuf
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__1591\ : CascadeBuf
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1589\ : CascadeBuf
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__10421\,
            I => \N__10418\
        );

    \I__1587\ : CascadeBuf
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__10415\,
            I => \N__10412\
        );

    \I__1585\ : CascadeBuf
    port map (
            O => \N__10412\,
            I => \N__10409\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__1583\ : CascadeBuf
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__1581\ : CascadeBuf
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__1579\ : CascadeBuf
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__1577\ : CascadeBuf
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1575\ : CascadeBuf
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__1573\ : CascadeBuf
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \N__10370\
        );

    \I__1571\ : CascadeBuf
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__1569\ : CascadeBuf
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__1567\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__1565\ : Span12Mux_s5_v
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__1564\ : Span12Mux_h
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__10346\,
            I => \M_this_vga_signals_address_8\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__10343\,
            I => \this_vga_signals.address_m6_0_1_cascade_\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10336\
        );

    \I__1560\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10330\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__10336\,
            I => \N__10327\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10335\,
            I => \N__10320\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10320\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10320\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__10330\,
            I => \this_vga_signals.address_mZ0Z1\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__10327\,
            I => \this_vga_signals.address_mZ0Z1\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__10320\,
            I => \this_vga_signals.address_mZ0Z1\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \this_vga_signals.G_12_0_3_cascade_\
        );

    \I__1551\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__10307\,
            I => \N__10303\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10300\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__10303\,
            I => \this_vga_signals.if_m4_0_1\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__10300\,
            I => \this_vga_signals.if_m4_0_1\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__10295\,
            I => \this_vga_signals_un17_address_if_N_8_mux_cascade_\
        );

    \I__1545\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__10289\,
            I => \this_vga_signals.N_10_0\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \N_6_i_cascade_\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__10277\,
            I => \this_vga_signals.N_18_0\
        );

    \I__1539\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10271\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__10268\,
            I => \this_vga_signals.g0_6_1\
        );

    \I__1536\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__10262\,
            I => \this_vga_signals.G_12_0_x3_0\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1532\ : Span4Mux_h
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__10250\,
            I => \this_vga_signals.g0_6_0_0_1\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__10247\,
            I => \this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__10244\,
            I => \N__10236\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10231\
        );

    \I__1527\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10226\
        );

    \I__1526\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10226\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10219\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10216\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10213\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10208\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10208\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10231\,
            I => \N__10203\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__10226\,
            I => \N__10203\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10196\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10196\
        );

    \I__1516\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10196\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10222\,
            I => \N__10193\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__10219\,
            I => \this_vga_signals.mult1_un61_sum_axb3\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10216\,
            I => \this_vga_signals.mult1_un61_sum_axb3\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__10213\,
            I => \this_vga_signals.mult1_un61_sum_axb3\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__10208\,
            I => \this_vga_signals.mult1_un61_sum_axb3\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__10203\,
            I => \this_vga_signals.mult1_un61_sum_axb3\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10196\,
            I => \this_vga_signals.mult1_un61_sum_axb3\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__10193\,
            I => \this_vga_signals.mult1_un61_sum_axb3\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10178\,
            I => \this_vga_signals.if_m4_0_1_0_cascade_\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10169\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10169\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__10169\,
            I => \this_vga_signals.mult1_un54_sum_axbxc5\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__10166\,
            I => \N__10162\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10165\,
            I => \N__10151\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10151\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10151\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10144\
        );

    \I__1498\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10144\
        );

    \I__1497\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10137\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__10151\,
            I => \N__10134\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__10150\,
            I => \N__10131\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10125\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10144\,
            I => \N__10122\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10117\
        );

    \I__1491\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10117\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10112\
        );

    \I__1489\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10112\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__10137\,
            I => \N__10107\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__10134\,
            I => \N__10107\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10102\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10102\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10097\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10128\,
            I => \N__10097\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__10125\,
            I => \this_vga_signals.un12_address_cry_7_c_RNI32HB\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__10122\,
            I => \this_vga_signals.un12_address_cry_7_c_RNI32HB\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10117\,
            I => \this_vga_signals.un12_address_cry_7_c_RNI32HB\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__10112\,
            I => \this_vga_signals.un12_address_cry_7_c_RNI32HB\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__10107\,
            I => \this_vga_signals.un12_address_cry_7_c_RNI32HB\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__10102\,
            I => \this_vga_signals.un12_address_cry_7_c_RNI32HB\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10097\,
            I => \this_vga_signals.un12_address_cry_7_c_RNI32HB\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__10076\,
            I => \this_vga_signals.if_m2_3_0\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10070\,
            I => \this_vga_signals.mult1_un61_sum_axb3_1\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__10064\,
            I => \this_vga_signals.G_12_0_3_1\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__10061\,
            I => \this_vga_signals.N_9_cascade_\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10052\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10052\,
            I => \this_vga_signals.g1_1\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__10049\,
            I => \this_vga_signals.mult1_un61_sum_axb3_0_cascade_\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__10046\,
            I => \this_vga_signals.g0_4_0_1_cascade_\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10039\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10036\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10039\,
            I => \N__10033\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__10036\,
            I => \this_vga_signals.g1_1_0\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__10033\,
            I => \this_vga_signals.g1_1_0\
        );

    \I__1457\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10016\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10016\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10016\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10013\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10006\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10006\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10016\,
            I => \N__10003\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10013\,
            I => \N__9992\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10012\,
            I => \N__9987\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9987\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__10006\,
            I => \N__9982\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__10003\,
            I => \N__9982\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10002\,
            I => \N__9977\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9977\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9968\
        );

    \I__1442\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9968\
        );

    \I__1441\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9968\
        );

    \I__1440\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9968\
        );

    \I__1439\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9963\
        );

    \I__1438\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9963\
        );

    \I__1437\ : Odrv12
    port map (
            O => \N__9992\,
            I => \this_vga_signals.mult1_un54_sum_axb3_out\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__9987\,
            I => \this_vga_signals.mult1_un54_sum_axb3_out\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__9982\,
            I => \this_vga_signals.mult1_un54_sum_axb3_out\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__9977\,
            I => \this_vga_signals.mult1_un54_sum_axb3_out\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__9968\,
            I => \this_vga_signals.mult1_un54_sum_axb3_out\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__9963\,
            I => \this_vga_signals.mult1_un54_sum_axb3_out\
        );

    \I__1431\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__9947\,
            I => \N__9941\
        );

    \I__1429\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9938\
        );

    \I__1428\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9933\
        );

    \I__1427\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9933\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__9941\,
            I => \this_vga_signals.mult1_un54_sum_axb4\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__9938\,
            I => \this_vga_signals.mult1_un54_sum_axb4\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__9933\,
            I => \this_vga_signals.mult1_un54_sum_axb4\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__9926\,
            I => \N__9922\
        );

    \I__1422\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9915\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9912\
        );

    \I__1420\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9907\
        );

    \I__1419\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9907\
        );

    \I__1418\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9902\
        );

    \I__1417\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9902\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__9915\,
            I => \this_vga_signals.mult1_un47_sum_c5\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__9912\,
            I => \this_vga_signals.mult1_un47_sum_c5\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__9907\,
            I => \this_vga_signals.mult1_un47_sum_c5\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__9902\,
            I => \this_vga_signals.mult1_un47_sum_c5\
        );

    \I__1412\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9890\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__9890\,
            I => \this_vga_signals.mult1_un61_sum_axb4_x0\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__9887\,
            I => \this_vga_signals.mult1_un54_sum_ac0_7_cascade_\
        );

    \I__1409\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__9881\,
            I => \this_vga_signals.mult1_un61_sum_axb4_x1\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__9878\,
            I => \this_vga_signals.mult1_un61_sum_axb4_i_cascade_\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__9875\,
            I => \this_vga_signals.mult1_un61_sum_ac0_5_cascade_\
        );

    \I__1405\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__9869\,
            I => \this_vga_signals.mult1_un61_sum_axb4_i\
        );

    \I__1403\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9863\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__9863\,
            I => \N__9859\
        );

    \I__1401\ : InMux
    port map (
            O => \N__9862\,
            I => \N__9856\
        );

    \I__1400\ : Span4Mux_h
    port map (
            O => \N__9859\,
            I => \N__9853\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__9856\,
            I => \N__9850\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__9853\,
            I => \this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__9850\,
            I => \this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__9845\,
            I => \this_vga_signals.M_vcounter_q_RNI8OSG6BZ0Z_2_cascade_\
        );

    \I__1395\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9836\
        );

    \I__1394\ : InMux
    port map (
            O => \N__9841\,
            I => \N__9836\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9836\,
            I => \this_vga_signals.mult1_un61_sum_axb1_0\
        );

    \I__1392\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9826\
        );

    \I__1391\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9826\
        );

    \I__1390\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9817\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__9826\,
            I => \N__9814\
        );

    \I__1388\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9811\
        );

    \I__1387\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9806\
        );

    \I__1386\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9806\
        );

    \I__1385\ : InMux
    port map (
            O => \N__9822\,
            I => \N__9799\
        );

    \I__1384\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9799\
        );

    \I__1383\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9799\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__9817\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__9814\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__9811\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__9806\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__9799\,
            I => \this_vga_signals.mult1_un54_sum_c3\
        );

    \I__1377\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9785\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__9785\,
            I => \this_vga_signals.address_m35_1\
        );

    \I__1375\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9776\
        );

    \I__1374\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9773\
        );

    \I__1373\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9770\
        );

    \I__1372\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9767\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__9776\,
            I => \N__9760\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__9773\,
            I => \N__9757\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__9770\,
            I => \N__9752\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__9767\,
            I => \N__9752\
        );

    \I__1367\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9747\
        );

    \I__1366\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9747\
        );

    \I__1365\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9742\
        );

    \I__1364\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9742\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__9760\,
            I => \this_vga_signals.N_75_mux\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__9757\,
            I => \this_vga_signals.N_75_mux\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__9752\,
            I => \this_vga_signals.N_75_mux\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__9747\,
            I => \this_vga_signals.N_75_mux\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__9742\,
            I => \this_vga_signals.N_75_mux\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__1357\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9721\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9716\
        );

    \I__1355\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9716\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__9725\,
            I => \N__9713\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__9724\,
            I => \N__9710\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__9721\,
            I => \N__9706\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__9716\,
            I => \N__9703\
        );

    \I__1350\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9700\
        );

    \I__1349\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9697\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__9709\,
            I => \N__9694\
        );

    \I__1347\ : Span4Mux_v
    port map (
            O => \N__9706\,
            I => \N__9689\
        );

    \I__1346\ : Span4Mux_v
    port map (
            O => \N__9703\,
            I => \N__9689\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__9700\,
            I => \N__9686\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__9697\,
            I => \N__9683\
        );

    \I__1343\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9680\
        );

    \I__1342\ : Sp12to4
    port map (
            O => \N__9689\,
            I => \N__9677\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__9686\,
            I => \N__9674\
        );

    \I__1340\ : Sp12to4
    port map (
            O => \N__9683\,
            I => \N__9669\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__9680\,
            I => \N__9669\
        );

    \I__1338\ : Odrv12
    port map (
            O => \N__9677\,
            I => \this_vga_signals.N_84\
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__9674\,
            I => \this_vga_signals.N_84\
        );

    \I__1336\ : Odrv12
    port map (
            O => \N__9669\,
            I => \this_vga_signals.N_84\
        );

    \I__1335\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9659\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__9659\,
            I => \N__9656\
        );

    \I__1333\ : Span4Mux_h
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__9653\,
            I => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_2\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__1330\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9644\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__9644\,
            I => \this_vga_signals.address_m31_1\
        );

    \I__1328\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9638\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__9638\,
            I => \this_vga_signals.address_i2_mux_4\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__9635\,
            I => \N__9630\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9627\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9622\
        );

    \I__1323\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9622\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__9627\,
            I => \this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__9622\,
            I => \this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9614\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__9614\,
            I => \this_vga_signals.address_N_9_0\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__9611\,
            I => \this_vga_signals.address_N_33_cascade_\
        );

    \I__1317\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__9605\,
            I => \this_vga_signals.address_N_34\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9586\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9586\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9586\
        );

    \I__1312\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9586\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9586\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9583\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__9586\,
            I => \this_vga_signals.M_vstate_qZ0Z_1\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__9583\,
            I => \this_vga_signals.M_vstate_qZ0Z_1\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__9578\,
            I => \this_vga_signals.m35_e_1_cascade_\
        );

    \I__1306\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9572\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9568\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9565\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__9568\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_0\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__9565\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_0\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__9557\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1\
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__9554\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__9551\,
            I => \N__9547\
        );

    \I__1297\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9544\
        );

    \I__1296\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9541\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__9544\,
            I => \this_vga_signals.mult1_un68_sum_c2\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__9541\,
            I => \this_vga_signals.mult1_un68_sum_c2\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__9536\,
            I => \this_vga_signals.address_N_9_0_cascade_\
        );

    \I__1292\ : InMux
    port map (
            O => \N__9533\,
            I => \N__9530\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__9530\,
            I => \this_vga_signals.address_N_10_0\
        );

    \I__1290\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9523\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9520\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__9523\,
            I => \this_vga_signals.address_N_3\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__9520\,
            I => \this_vga_signals.address_N_3\
        );

    \I__1286\ : IoInMux
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__9512\,
            I => \N__9509\
        );

    \I__1284\ : IoSpan4Mux
    port map (
            O => \N__9509\,
            I => \N__9506\
        );

    \I__1283\ : IoSpan4Mux
    port map (
            O => \N__9506\,
            I => \N__9503\
        );

    \I__1282\ : Span4Mux_s3_v
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__9497\,
            I => \N__9494\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__9494\,
            I => vsync_c
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__9491\,
            I => \this_vga_signals.N_52_cascade_\
        );

    \I__1277\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9485\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__9485\,
            I => \this_vga_signals.N_76_mux\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__9482\,
            I => \this_vga_signals.N_76_mux_cascade_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9473\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9473\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__9473\,
            I => \this_vga_signals.N_72_mux\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__9470\,
            I => \this_vga_signals.N_55_cascade_\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__9467\,
            I => \this_vga_signals.M_vstate_q_RNO_1Z0Z_0_cascade_\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9464\,
            I => \N__9461\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__9461\,
            I => \this_vga_signals.M_vstate_q_RNO_2Z0Z_0\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__9455\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_3\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__9452\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\
        );

    \I__1264\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__9446\,
            I => \this_vga_signals.mult1_un54_sum_c4\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__9443\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_4_cascade_\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__9440\,
            I => \this_vga_signals.if_m4_0_1_cascade_\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__9437\,
            I => \this_vga_signals.G_12_0_x3_0_cascade_\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__9434\,
            I => \N__9430\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__9433\,
            I => \N__9425\
        );

    \I__1257\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9417\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9417\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9408\
        );

    \I__1254\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9408\
        );

    \I__1253\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9408\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9408\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9405\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__9417\,
            I => \this_vga_signals.un12_address_cry_10_c_RNINP5K\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__9408\,
            I => \this_vga_signals.un12_address_cry_10_c_RNINP5K\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__9405\,
            I => \this_vga_signals.un12_address_cry_10_c_RNINP5K\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__9398\,
            I => \this_vga_signals.un12_address_cry_9_c_RNIVF1R_cascade_\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__9395\,
            I => \N__9387\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__9394\,
            I => \N__9384\
        );

    \I__1244\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9378\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9378\
        );

    \I__1242\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9369\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9369\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9369\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9369\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9383\,
            I => \N__9366\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9378\,
            I => \this_vga_signals.un12_address_cry_9_c_RNIEJOE\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__9369\,
            I => \this_vga_signals.un12_address_cry_9_c_RNIEJOE\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9366\,
            I => \this_vga_signals.un12_address_cry_9_c_RNIEJOE\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__9359\,
            I => \this_vga_signals.mult1_un47_sum_c5_cascade_\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__9356\,
            I => \this_vga_signals.mult1_un61_sum_axb3_x1_cascade_\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__9353\,
            I => \this_vga_signals.mult1_un61_sum_axb3_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9347\,
            I => \this_vga_signals.if_m5_sn\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__9344\,
            I => \this_vga_signals.if_m5_rn_0_cascade_\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__9341\,
            I => \this_vga_signals.mult1_un68_sum_c5_cascade_\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__1226\ : CascadeBuf
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__1224\ : CascadeBuf
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__1222\ : CascadeBuf
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__1220\ : CascadeBuf
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__1218\ : CascadeBuf
    port map (
            O => \N__9311\,
            I => \N__9308\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__1216\ : CascadeBuf
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__9302\,
            I => \N__9299\
        );

    \I__1214\ : CascadeBuf
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__1212\ : CascadeBuf
    port map (
            O => \N__9293\,
            I => \N__9290\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__1210\ : CascadeBuf
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__1208\ : CascadeBuf
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__1206\ : CascadeBuf
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__1204\ : CascadeBuf
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__1202\ : CascadeBuf
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__1200\ : CascadeBuf
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__1198\ : CascadeBuf
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__1194\ : Span12Mux_h
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__1193\ : Span12Mux_v
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__1192\ : Odrv12
    port map (
            O => \N__9233\,
            I => \M_this_vga_signals_address_4\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__9230\,
            I => \this_vga_signals.mult1_un54_sum_ac0_8_cascade_\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__9224\,
            I => \this_vga_signals.g1_1_1\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9217\
        );

    \I__1187\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9211\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9206\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9201\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9201\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9214\,
            I => \N__9197\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__9211\,
            I => \N__9194\
        );

    \I__1181\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9189\
        );

    \I__1180\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9189\
        );

    \I__1179\ : Span4Mux_h
    port map (
            O => \N__9206\,
            I => \N__9184\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__9201\,
            I => \N__9184\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9181\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9197\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__9194\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__9189\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__9184\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__9181\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9166\
        );

    \I__1170\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9163\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9166\,
            I => \N__9158\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9163\,
            I => \N__9158\
        );

    \I__1167\ : Odrv12
    port map (
            O => \N__9158\,
            I => \this_vga_signals.M_hcounter_q_i_11\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9149\
        );

    \I__1165\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9149\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__9149\,
            I => \this_vga_signals.un12_address_cry_9_THRU_CO\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9136\
        );

    \I__1162\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9136\
        );

    \I__1161\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9127\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9127\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9127\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9127\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__9136\,
            I => \this_vga_signals.un12_address_cry_9_c_RNIVF1R\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__9127\,
            I => \this_vga_signals.un12_address_cry_9_c_RNIVF1R\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__9122\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_cascade_\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__9119\,
            I => \N__9114\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9108\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9108\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9103\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9103\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__9108\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__9103\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9092\
        );

    \I__1146\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9092\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9092\,
            I => \this_vga_signals.mult1_un61_sum_c2\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9083\,
            I => \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2\
        );

    \I__1141\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9077\,
            I => \this_vga_signals.address_i3_mux_i\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__9074\,
            I => \this_vga_signals.address_m27_ns_1_cascade_\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__9071\,
            I => \this_vga_signals.address_i2_mux_3_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__9065\,
            I => \this_vga_signals.address_i2_mux_2\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__1133\ : Span4Mux_h
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__9053\,
            I => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_1\
        );

    \I__1131\ : IoInMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__1129\ : Span4Mux_s3_h
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__9041\,
            I => \N__9037\
        );

    \I__1127\ : IoInMux
    port map (
            O => \N__9040\,
            I => \N__9034\
        );

    \I__1126\ : Span4Mux_v
    port map (
            O => \N__9037\,
            I => \N__9031\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__9034\,
            I => \N__9028\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__9031\,
            I => \N__9023\
        );

    \I__1123\ : Span4Mux_s3_h
    port map (
            O => \N__9028\,
            I => \N__9023\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__1121\ : Span4Mux_h
    port map (
            O => \N__9020\,
            I => \N__9017\
        );

    \I__1120\ : Odrv4
    port map (
            O => \N__9017\,
            I => rgb_c_0
        );

    \I__1119\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9009\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__9013\,
            I => \N__9004\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8997\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__9009\,
            I => \N__8993\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8988\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8988\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8985\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__9003\,
            I => \N__8982\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8979\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__9001\,
            I => \N__8976\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8973\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8970\
        );

    \I__1107\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8967\
        );

    \I__1106\ : Span4Mux_v
    port map (
            O => \N__8993\,
            I => \N__8962\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8962\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8959\
        );

    \I__1103\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8956\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__8979\,
            I => \N__8953\
        );

    \I__1101\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8950\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__8973\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__8970\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__8967\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1097\ : Odrv4
    port map (
            O => \N__8962\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__8959\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__8956\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1094\ : Odrv12
    port map (
            O => \N__8953\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__8950\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1092\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__8930\,
            I => \this_vga_signals.address_m1_1_1\
        );

    \I__1090\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8923\
        );

    \I__1089\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8920\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__8923\,
            I => \this_vga_signals.mult1_un54_sum_c2\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__8920\,
            I => \this_vga_signals.mult1_un54_sum_c2\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__8915\,
            I => \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2_cascade_\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1084\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__8906\,
            I => \this_vga_signals.mult1_un61_sum_c3_1\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__8903\,
            I => \this_vga_signals.mult1_un61_sum_c3_cascade_\
        );

    \I__1081\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8890\
        );

    \I__1080\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8885\
        );

    \I__1079\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8885\
        );

    \I__1078\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8874\
        );

    \I__1077\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8874\
        );

    \I__1076\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8874\
        );

    \I__1075\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8874\
        );

    \I__1074\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8874\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__8890\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__8885\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__8874\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1070\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8861\
        );

    \I__1069\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8861\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__8861\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_0\
        );

    \I__1067\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__8855\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_3_2\
        );

    \I__1065\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8848\
        );

    \I__1064\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8843\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__8848\,
            I => \N__8840\
        );

    \I__1062\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8837\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__8846\,
            I => \N__8833\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__8843\,
            I => \N__8825\
        );

    \I__1059\ : Span4Mux_v
    port map (
            O => \N__8840\,
            I => \N__8825\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8825\
        );

    \I__1057\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8822\
        );

    \I__1056\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8819\
        );

    \I__1055\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8816\
        );

    \I__1054\ : Span4Mux_h
    port map (
            O => \N__8825\,
            I => \N__8813\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8808\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__8819\,
            I => \N__8808\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__8816\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1050\ : Odrv4
    port map (
            O => \N__8813\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1049\ : Odrv12
    port map (
            O => \N__8808\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1048\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8797\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__8800\,
            I => \N__8794\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8791\
        );

    \I__1045\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8788\
        );

    \I__1044\ : Span4Mux_h
    port map (
            O => \N__8791\,
            I => \N__8785\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__8788\,
            I => \N__8782\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__8785\,
            I => \this_vga_signals.N_27\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__8782\,
            I => \this_vga_signals.N_27\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__8777\,
            I => \N__8770\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8765\
        );

    \I__1038\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8765\
        );

    \I__1037\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8762\
        );

    \I__1036\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8759\
        );

    \I__1035\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8756\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__8765\,
            I => \N__8752\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8749\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8759\,
            I => \N__8746\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__8756\,
            I => \N__8743\
        );

    \I__1030\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8740\
        );

    \I__1029\ : Span4Mux_h
    port map (
            O => \N__8752\,
            I => \N__8737\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__8749\,
            I => \N__8730\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__8746\,
            I => \N__8730\
        );

    \I__1026\ : Span4Mux_v
    port map (
            O => \N__8743\,
            I => \N__8730\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__8740\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__8737\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__8730\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__8717\,
            I => \this_vga_signals.hvisible_i_a2_2_0\
        );

    \I__1019\ : IoInMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__1017\ : Span4Mux_s2_h
    port map (
            O => \N__8708\,
            I => \N__8704\
        );

    \I__1016\ : IoInMux
    port map (
            O => \N__8707\,
            I => \N__8701\
        );

    \I__1015\ : Span4Mux_h
    port map (
            O => \N__8704\,
            I => \N__8698\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__8701\,
            I => \N__8695\
        );

    \I__1013\ : Span4Mux_h
    port map (
            O => \N__8698\,
            I => \N__8692\
        );

    \I__1012\ : Span12Mux_s10_h
    port map (
            O => \N__8695\,
            I => \N__8689\
        );

    \I__1011\ : Span4Mux_v
    port map (
            O => \N__8692\,
            I => \N__8686\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__8689\,
            I => rgb_c_4
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__8686\,
            I => rgb_c_4
        );

    \I__1008\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__8678\,
            I => \this_vga_signals.m30_3\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__8675\,
            I => \this_vga_signals.m30_4_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8667\
        );

    \I__1004\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8661\
        );

    \I__1003\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8658\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8655\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__8666\,
            I => \N__8652\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__8665\,
            I => \N__8649\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__8664\,
            I => \N__8643\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__8661\,
            I => \N__8639\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__8658\,
            I => \N__8636\
        );

    \I__996\ : Span4Mux_h
    port map (
            O => \N__8655\,
            I => \N__8633\
        );

    \I__995\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8630\
        );

    \I__994\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8625\
        );

    \I__993\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8625\
        );

    \I__992\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8622\
        );

    \I__991\ : InMux
    port map (
            O => \N__8646\,
            I => \N__8617\
        );

    \I__990\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8617\
        );

    \I__989\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8614\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__8639\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__8636\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__8633\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__8630\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__8625\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__8622\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8617\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__8614\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__980\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8593\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__8596\,
            I => \N__8584\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__8593\,
            I => \N__8580\
        );

    \I__977\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8577\
        );

    \I__976\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8574\
        );

    \I__975\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8571\
        );

    \I__974\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8568\
        );

    \I__973\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8565\
        );

    \I__972\ : InMux
    port map (
            O => \N__8587\,
            I => \N__8558\
        );

    \I__971\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8558\
        );

    \I__970\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8558\
        );

    \I__969\ : Span4Mux_v
    port map (
            O => \N__8580\,
            I => \N__8553\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__8577\,
            I => \N__8553\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__8574\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__8571\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__8568\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__8565\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__8558\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__8553\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__961\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8535\
        );

    \I__960\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8532\
        );

    \I__959\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8526\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8518\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__8532\,
            I => \N__8515\
        );

    \I__956\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8508\
        );

    \I__955\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8505\
        );

    \I__954\ : InMux
    port map (
            O => \N__8529\,
            I => \N__8502\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__8526\,
            I => \N__8499\
        );

    \I__952\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8494\
        );

    \I__951\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8494\
        );

    \I__950\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8489\
        );

    \I__949\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8489\
        );

    \I__948\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8486\
        );

    \I__947\ : Span4Mux_h
    port map (
            O => \N__8518\,
            I => \N__8483\
        );

    \I__946\ : Span4Mux_h
    port map (
            O => \N__8515\,
            I => \N__8480\
        );

    \I__945\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8477\
        );

    \I__944\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8470\
        );

    \I__943\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8470\
        );

    \I__942\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8470\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8465\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8465\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8502\,
            I => \N__8462\
        );

    \I__938\ : Span4Mux_h
    port map (
            O => \N__8499\,
            I => \N__8455\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__8494\,
            I => \N__8455\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8455\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__8486\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__8483\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__8480\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__8477\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8470\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__930\ : Odrv4
    port map (
            O => \N__8465\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__929\ : Odrv12
    port map (
            O => \N__8462\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__8455\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__8438\,
            I => \this_vga_signals.N_3_0_cascade_\
        );

    \I__926\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8430\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__8434\,
            I => \N__8421\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \N__8418\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__8430\,
            I => \N__8415\
        );

    \I__922\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8412\
        );

    \I__921\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8409\
        );

    \I__920\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8404\
        );

    \I__919\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8404\
        );

    \I__918\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8401\
        );

    \I__917\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8398\
        );

    \I__916\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8393\
        );

    \I__915\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8393\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__8415\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__8412\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__8409\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8404\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__8401\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__8398\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__8393\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__907\ : InMux
    port map (
            O => \N__8378\,
            I => \this_vga_signals.un12_address_cry_10\
        );

    \I__906\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8372\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__8372\,
            I => \N__8367\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__8371\,
            I => \N__8364\
        );

    \I__903\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8361\
        );

    \I__902\ : Span4Mux_v
    port map (
            O => \N__8367\,
            I => \N__8358\
        );

    \I__901\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8355\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8361\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__8358\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__8355\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__897\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8345\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__8345\,
            I => \N__8341\
        );

    \I__895\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8338\
        );

    \I__894\ : Span4Mux_h
    port map (
            O => \N__8341\,
            I => \N__8335\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__8338\,
            I => \this_vga_signals.N_49\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__8335\,
            I => \this_vga_signals.N_49\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__8330\,
            I => \N__8325\
        );

    \I__890\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8320\
        );

    \I__889\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8317\
        );

    \I__888\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8314\
        );

    \I__887\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8309\
        );

    \I__886\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8309\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__8320\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8317\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__8314\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__8309\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__881\ : IoInMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__879\ : Span4Mux_s3_v
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__878\ : Span4Mux_h
    port map (
            O => \N__8291\,
            I => \N__8287\
        );

    \I__877\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8284\
        );

    \I__876\ : Sp12to4
    port map (
            O => \N__8287\,
            I => \N__8281\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__8284\,
            I => \N__8278\
        );

    \I__874\ : Span12Mux_v
    port map (
            O => \N__8281\,
            I => \N__8274\
        );

    \I__873\ : Span12Mux_s10_h
    port map (
            O => \N__8278\,
            I => \N__8271\
        );

    \I__872\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8268\
        );

    \I__871\ : Odrv12
    port map (
            O => \N__8274\,
            I => \N_16\
        );

    \I__870\ : Odrv12
    port map (
            O => \N__8271\,
            I => \N_16\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__8268\,
            I => \N_16\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__8261\,
            I => \this_vga_signals.mult1_un61_sum_ac0_7_0_3_1_1_cascade_\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__8258\,
            I => \N__8253\
        );

    \I__866\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8250\
        );

    \I__865\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8247\
        );

    \I__864\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8244\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8241\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8247\,
            I => \N__8236\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__8244\,
            I => \N__8236\
        );

    \I__860\ : Span4Mux_h
    port map (
            O => \N__8241\,
            I => \N__8233\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__8236\,
            I => \N__8230\
        );

    \I__858\ : Odrv4
    port map (
            O => \N__8233\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__8230\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__856\ : InMux
    port map (
            O => \N__8225\,
            I => \this_vga_signals.un12_address_cry_1\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__854\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8214\
        );

    \I__853\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8211\
        );

    \I__852\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8208\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8214\,
            I => \N__8205\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8211\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__8208\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__8205\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__847\ : InMux
    port map (
            O => \N__8198\,
            I => \this_vga_signals.un12_address_cry_2\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__8195\,
            I => \N__8190\
        );

    \I__845\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8187\
        );

    \I__844\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8184\
        );

    \I__843\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8181\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8187\,
            I => \N__8178\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8184\,
            I => \N__8173\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__8181\,
            I => \N__8173\
        );

    \I__839\ : Span4Mux_h
    port map (
            O => \N__8178\,
            I => \N__8170\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__8170\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__8167\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__835\ : InMux
    port map (
            O => \N__8162\,
            I => \this_vga_signals.un12_address_cry_3\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__8159\,
            I => \N__8155\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__8158\,
            I => \N__8151\
        );

    \I__832\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8148\
        );

    \I__831\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8145\
        );

    \I__830\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8142\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8148\,
            I => \N__8139\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8134\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__8142\,
            I => \N__8134\
        );

    \I__826\ : Span4Mux_h
    port map (
            O => \N__8139\,
            I => \N__8131\
        );

    \I__825\ : Span4Mux_h
    port map (
            O => \N__8134\,
            I => \N__8128\
        );

    \I__824\ : Odrv4
    port map (
            O => \N__8131\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__8128\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__822\ : InMux
    port map (
            O => \N__8123\,
            I => \this_vga_signals.un12_address_cry_4\
        );

    \I__821\ : InMux
    port map (
            O => \N__8120\,
            I => \this_vga_signals.un12_address_cry_5\
        );

    \I__820\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8111\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__8116\,
            I => \N__8108\
        );

    \I__818\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8103\
        );

    \I__817\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8103\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8111\,
            I => \N__8100\
        );

    \I__815\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8097\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8103\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__8100\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__8097\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__811\ : InMux
    port map (
            O => \N__8090\,
            I => \this_vga_signals.un12_address_cry_6\
        );

    \I__810\ : InMux
    port map (
            O => \N__8087\,
            I => \bfn_11_18_0_\
        );

    \I__809\ : InMux
    port map (
            O => \N__8084\,
            I => \this_vga_signals.un12_address_cry_8\
        );

    \I__808\ : InMux
    port map (
            O => \N__8081\,
            I => \this_vga_signals.un12_address_cry_9\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__8078\,
            I => \this_vga_signals.address_m24_ns_1Z0Z_0_cascade_\
        );

    \I__806\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8068\
        );

    \I__804\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8060\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__8068\,
            I => \N__8057\
        );

    \I__802\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8054\
        );

    \I__801\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8049\
        );

    \I__800\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8049\
        );

    \I__799\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8044\
        );

    \I__798\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8044\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8060\,
            I => \N__8041\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__8057\,
            I => \this_vga_signals.mult1_un40_sum_c3\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8054\,
            I => \this_vga_signals.mult1_un40_sum_c3\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__8049\,
            I => \this_vga_signals.mult1_un40_sum_c3\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8044\,
            I => \this_vga_signals.mult1_un40_sum_c3\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__8041\,
            I => \this_vga_signals.mult1_un40_sum_c3\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__8030\,
            I => \this_vga_signals.mult1_un54_sum_c2_cascade_\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__789\ : InMux
    port map (
            O => \N__8024\,
            I => \N__8017\
        );

    \I__788\ : InMux
    port map (
            O => \N__8023\,
            I => \N__8017\
        );

    \I__787\ : InMux
    port map (
            O => \N__8022\,
            I => \N__8014\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__8017\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8014\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__8009\,
            I => \this_vga_signals.mult1_un54_sum_c3_cascade_\
        );

    \I__783\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__8003\,
            I => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_0\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__8000\,
            I => \N__7995\
        );

    \I__780\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7991\
        );

    \I__779\ : InMux
    port map (
            O => \N__7998\,
            I => \N__7988\
        );

    \I__778\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7985\
        );

    \I__777\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7982\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7975\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__7988\,
            I => \N__7975\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7975\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__7982\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__7975\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__771\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7966\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__7969\,
            I => \N__7962\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__7966\,
            I => \N__7959\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__7965\,
            I => \N__7956\
        );

    \I__767\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7953\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__7959\,
            I => \N__7950\
        );

    \I__765\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7947\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__7953\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__763\ : Odrv4
    port map (
            O => \N__7950\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__7947\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__761\ : InMux
    port map (
            O => \N__7940\,
            I => \this_vga_signals.un12_address_cry_0\
        );

    \I__760\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7931\
        );

    \I__759\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7924\
        );

    \I__758\ : InMux
    port map (
            O => \N__7935\,
            I => \N__7924\
        );

    \I__757\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7924\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__7931\,
            I => \N__7919\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__7924\,
            I => \N__7916\
        );

    \I__754\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7911\
        );

    \I__753\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7911\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__7919\,
            I => \this_vga_signals.N_70\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__7916\,
            I => \this_vga_signals.N_70\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__7911\,
            I => \this_vga_signals.N_70\
        );

    \I__749\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7900\
        );

    \I__748\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7897\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__7900\,
            I => \this_vga_signals.SUM_0\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__7897\,
            I => \this_vga_signals.SUM_0\
        );

    \I__745\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__7889\,
            I => \this_vga_signals.mult1_un40_sum_axbxc1\
        );

    \I__743\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__7883\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__7880\,
            I => \this_vga_signals.mult1_un40_sum_axbxc1_cascade_\
        );

    \I__740\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7873\
        );

    \I__739\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7870\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__7873\,
            I => \this_vga_signals.mult1_un47_sum_ac0_1\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__7870\,
            I => \this_vga_signals.mult1_un47_sum_ac0_1\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__7865\,
            I => \this_vga_signals.mult1_un47_sum_c3_cascade_\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__7862\,
            I => \N__7859\
        );

    \I__734\ : InMux
    port map (
            O => \N__7859\,
            I => \N__7853\
        );

    \I__733\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7853\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__7850\,
            I => \this_vga_signals.N_13_0\
        );

    \I__730\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7841\
        );

    \I__729\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7841\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__7841\,
            I => \this_vga_signals.if_i1_mux\
        );

    \I__727\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7835\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__7835\,
            I => \N__7832\
        );

    \I__725\ : Odrv4
    port map (
            O => \N__7832\,
            I => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_3\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__7829\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__7826\,
            I => \this_vga_signals.i9_mux_cascade_\
        );

    \I__722\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__7820\,
            I => \this_vga_signals.i9_mux\
        );

    \I__720\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7810\
        );

    \I__719\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7810\
        );

    \I__718\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7807\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__7810\,
            I => \this_vga_signals.address_1_c5_i\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__7807\,
            I => \this_vga_signals.address_1_c5_i\
        );

    \I__715\ : IoInMux
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__7799\,
            I => \N__7795\
        );

    \I__713\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7792\
        );

    \I__712\ : IoSpan4Mux
    port map (
            O => \N__7795\,
            I => \N__7789\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__7792\,
            I => \N__7786\
        );

    \I__710\ : Span4Mux_s1_h
    port map (
            O => \N__7789\,
            I => \N__7783\
        );

    \I__709\ : Span4Mux_v
    port map (
            O => \N__7786\,
            I => \N__7779\
        );

    \I__708\ : Span4Mux_h
    port map (
            O => \N__7783\,
            I => \N__7776\
        );

    \I__707\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7773\
        );

    \I__706\ : Span4Mux_h
    port map (
            O => \N__7779\,
            I => \N__7770\
        );

    \I__705\ : Span4Mux_h
    port map (
            O => \N__7776\,
            I => \N__7765\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__7773\,
            I => \N__7765\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__7770\,
            I => \N__7760\
        );

    \I__702\ : Span4Mux_v
    port map (
            O => \N__7765\,
            I => \N__7760\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__7760\,
            I => port_nmib_c
        );

    \I__700\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7752\
        );

    \I__699\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7747\
        );

    \I__698\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7747\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__7752\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__7747\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__695\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7736\
        );

    \I__694\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7736\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__7733\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCNZ0\
        );

    \I__691\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7726\
        );

    \I__690\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7723\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7720\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7717\
        );

    \I__687\ : Span4Mux_h
    port map (
            O => \N__7720\,
            I => \N__7714\
        );

    \I__686\ : Span4Mux_h
    port map (
            O => \N__7717\,
            I => \N__7711\
        );

    \I__685\ : Odrv4
    port map (
            O => \N__7714\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__7711\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0\
        );

    \I__683\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7700\
        );

    \I__682\ : InMux
    port map (
            O => \N__7705\,
            I => \N__7695\
        );

    \I__681\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7695\
        );

    \I__680\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7692\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__7700\,
            I => \N__7689\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7684\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__7692\,
            I => \N__7684\
        );

    \I__676\ : Span4Mux_v
    port map (
            O => \N__7689\,
            I => \N__7679\
        );

    \I__675\ : Span4Mux_v
    port map (
            O => \N__7684\,
            I => \N__7679\
        );

    \I__674\ : Sp12to4
    port map (
            O => \N__7679\,
            I => \N__7676\
        );

    \I__673\ : Span12Mux_h
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__672\ : Span12Mux_v
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__671\ : Odrv12
    port map (
            O => \N__7670\,
            I => rst_n_c
        );

    \I__670\ : InMux
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__668\ : Odrv4
    port map (
            O => \N__7661\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__667\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__7655\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__7652\,
            I => \this_vga_signals.address_1_c4_cascade_\
        );

    \I__664\ : InMux
    port map (
            O => \N__7649\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_9\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__7646\,
            I => \N__7642\
        );

    \I__662\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7636\
        );

    \I__661\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7633\
        );

    \I__660\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7630\
        );

    \I__659\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7627\
        );

    \I__658\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7624\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__7636\,
            I => \N__7619\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__7633\,
            I => \N__7619\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__7630\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__7627\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__7624\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__652\ : Odrv12
    port map (
            O => \N__7619\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__651\ : InMux
    port map (
            O => \N__7610\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_10\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__7607\,
            I => \this_vga_signals.g1_0_0_a2_0_cascade_\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__7604\,
            I => \this_vga_signals.g0_11_1_cascade_\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__647\ : InMux
    port map (
            O => \N__7598\,
            I => \N__7592\
        );

    \I__646\ : InMux
    port map (
            O => \N__7597\,
            I => \N__7592\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__7592\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__644\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__7586\,
            I => \N__7582\
        );

    \I__642\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7579\
        );

    \I__641\ : Span4Mux_v
    port map (
            O => \N__7582\,
            I => \N__7574\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7574\
        );

    \I__639\ : Odrv4
    port map (
            O => \N__7574\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KANZ0\
        );

    \I__638\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7562\
        );

    \I__637\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7562\
        );

    \I__636\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7562\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__7562\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__633\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__7553\,
            I => \this_vga_signals.N_2\
        );

    \I__631\ : InMux
    port map (
            O => \N__7550\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__630\ : InMux
    port map (
            O => \N__7547\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_0\
        );

    \I__629\ : InMux
    port map (
            O => \N__7544\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_1\
        );

    \I__628\ : InMux
    port map (
            O => \N__7541\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_2\
        );

    \I__627\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__7535\,
            I => \N__7531\
        );

    \I__625\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7528\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__7531\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__7528\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0\
        );

    \I__622\ : InMux
    port map (
            O => \N__7523\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_3\
        );

    \I__621\ : InMux
    port map (
            O => \N__7520\,
            I => \N__7517\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__7517\,
            I => \N__7513\
        );

    \I__619\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7510\
        );

    \I__618\ : Odrv4
    port map (
            O => \N__7513\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__7510\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0\
        );

    \I__616\ : InMux
    port map (
            O => \N__7505\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_4\
        );

    \I__615\ : InMux
    port map (
            O => \N__7502\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_5\
        );

    \I__614\ : InMux
    port map (
            O => \N__7499\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_6\
        );

    \I__613\ : InMux
    port map (
            O => \N__7496\,
            I => \bfn_9_24_0_\
        );

    \I__612\ : InMux
    port map (
            O => \N__7493\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_8\
        );

    \I__611\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__7487\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__7484\,
            I => \this_vga_signals.mult1_un40_sum_c3_cascade_\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__7481\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__7478\,
            I => \this_vga_signals.mult1_un47_sum_ac0_2_cascade_\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__7475\,
            I => \this_vga_signals.N_2_cascade_\
        );

    \I__605\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7468\
        );

    \I__604\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7465\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__7468\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__7465\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__7460\,
            I => \this_vga_signals.N_70_cascade_\
        );

    \I__600\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__7454\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_1_0\
        );

    \I__598\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7445\
        );

    \I__597\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7445\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__7445\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__595\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7439\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__7439\,
            I => \this_vga_signals.m44_0_0\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__7436\,
            I => \this_vga_signals.M_vcounter_q_RNIQE2J1Z0Z_9_cascade_\
        );

    \I__592\ : InMux
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__7430\,
            I => \this_vga_signals.M_vcounter_q_fast_RNI3BJLZ0Z_4\
        );

    \I__590\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__7424\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__588\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7417\
        );

    \I__587\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7414\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__7417\,
            I => \N__7411\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__7414\,
            I => \N__7408\
        );

    \I__584\ : Span4Mux_h
    port map (
            O => \N__7411\,
            I => \N__7405\
        );

    \I__583\ : Span4Mux_h
    port map (
            O => \N__7408\,
            I => \N__7402\
        );

    \I__582\ : Odrv4
    port map (
            O => \N__7405\,
            I => \this_vga_signals.N_32\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__7402\,
            I => \this_vga_signals.N_32\
        );

    \I__580\ : InMux
    port map (
            O => \N__7397\,
            I => \N__7392\
        );

    \I__579\ : InMux
    port map (
            O => \N__7396\,
            I => \N__7389\
        );

    \I__578\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7385\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__7392\,
            I => \N__7382\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__7389\,
            I => \N__7379\
        );

    \I__575\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7376\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__7385\,
            I => \N__7373\
        );

    \I__573\ : Span4Mux_v
    port map (
            O => \N__7382\,
            I => \N__7370\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__7379\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__7376\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__7373\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__7370\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__7361\,
            I => \N__7358\
        );

    \I__567\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7355\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__7355\,
            I => \this_vga_signals.N_26\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__7352\,
            I => \this_vga_signals.N_26_cascade_\
        );

    \I__564\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__7346\,
            I => \N__7342\
        );

    \I__562\ : InMux
    port map (
            O => \N__7345\,
            I => \N__7339\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__7342\,
            I => \N__7336\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__7339\,
            I => \N__7333\
        );

    \I__559\ : Sp12to4
    port map (
            O => \N__7336\,
            I => \N__7329\
        );

    \I__558\ : Span4Mux_h
    port map (
            O => \N__7333\,
            I => \N__7326\
        );

    \I__557\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7323\
        );

    \I__556\ : Odrv12
    port map (
            O => \N__7329\,
            I => \this_vga_signals.N_51\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__7326\,
            I => \this_vga_signals.N_51\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__7323\,
            I => \this_vga_signals.N_51\
        );

    \I__553\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7310\
        );

    \I__552\ : InMux
    port map (
            O => \N__7315\,
            I => \N__7310\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7307\
        );

    \I__550\ : Span4Mux_h
    port map (
            O => \N__7307\,
            I => \N__7304\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__7304\,
            I => \this_vga_signals.N_273\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__7301\,
            I => \this_vga_signals.N_18_cascade_\
        );

    \I__547\ : IoInMux
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7292\
        );

    \I__545\ : IoSpan4Mux
    port map (
            O => \N__7292\,
            I => \N__7289\
        );

    \I__544\ : Span4Mux_s2_v
    port map (
            O => \N__7289\,
            I => \N__7286\
        );

    \I__543\ : Span4Mux_v
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__541\ : Odrv4
    port map (
            O => \N__7280\,
            I => \this_vga_signals_N_274_i\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__7277\,
            I => \this_vga_signals.hvisible_i_a2_0_3_0_cascade_\
        );

    \I__539\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7266\
        );

    \I__538\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7266\
        );

    \I__537\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7263\
        );

    \I__536\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7258\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__7266\,
            I => \N__7253\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__7263\,
            I => \N__7253\
        );

    \I__533\ : InMux
    port map (
            O => \N__7262\,
            I => \N__7250\
        );

    \I__532\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7247\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__7258\,
            I => \N__7242\
        );

    \I__530\ : Span4Mux_h
    port map (
            O => \N__7253\,
            I => \N__7242\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__7250\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__7247\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__7242\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__7235\,
            I => \this_vga_signals.N_49_cascade_\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__7232\,
            I => \this_vga_signals.N_29_cascade_\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__7229\,
            I => \this_vga_signals.N_40_cascade_\
        );

    \I__523\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__521\ : Odrv4
    port map (
            O => \N__7220\,
            I => \this_vga_signals.N_20\
        );

    \I__520\ : IoInMux
    port map (
            O => \N__7217\,
            I => \N__7214\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__7214\,
            I => port_rw_c_i
        );

    \I__518\ : IoInMux
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__516\ : Odrv12
    port map (
            O => \N__7205\,
            I => port_nmib_c_i
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un12_address_cry_7\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_6_cry_7\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_19_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_23_0_\
        );

    \IN_MUX_bfv_19_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_current_address_q_cry_7\,
            carryinitout => \bfn_19_24_0_\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17739\,
            GLOBALBUFFEROUTPUT => \N_339_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \port_data_rw_obuf_RNO_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19705\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => port_rw_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIL6FA3_0_9_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7798\,
            lcout => port_nmib_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_6_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13486\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17351\,
            ce => 'H',
            sr => \N__15473\
        );

    \this_vga_signals.M_hstate_q_RNO_2_0_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001110111"
        )
    port map (
            in0 => \N__7273\,
            in1 => \N__8832\,
            in2 => \_gnd_net_\,
            in3 => \N__8755\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_1_0_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__8801\,
            in1 => \N__7395\,
            in2 => \N__7232\,
            in3 => \N__9221\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_0_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110001"
        )
    port map (
            in0 => \N__7274\,
            in1 => \N__7420\,
            in2 => \N__7229\,
            in3 => \N__7345\,
            lcout => \this_vga_signals.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_9_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10025\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17351\,
            ce => 'H',
            sr => \N__15473\
        );

    \this_vga_signals.M_hcounter_q_2_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14012\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17357\,
            ce => 'H',
            sr => \N__15471\
        );

    \this_vga_signals.M_hcounter_q_4_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12977\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17357\,
            ce => 'H',
            sr => \N__15471\
        );

    \this_vga_signals.M_hcounter_q_5_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13762\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17357\,
            ce => 'H',
            sr => \N__15471\
        );

    \this_vga_signals.M_hstate_q_0_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000010"
        )
    port map (
            in0 => \N__7315\,
            in1 => \N__7226\,
            in2 => \N__17737\,
            in3 => \N__7388\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_1_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__7421\,
            in1 => \N__7261\,
            in2 => \_gnd_net_\,
            in3 => \N__7349\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_1_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001110"
        )
    port map (
            in0 => \N__7316\,
            in1 => \N__7262\,
            in2 => \N__7301\,
            in3 => \N__17738\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17362\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__7396\,
            in1 => \N__7271\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals_N_274_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_13_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7782\,
            in1 => \N__8290\,
            in2 => \_gnd_net_\,
            in3 => \N__8075\,
            lcout => \this_vram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_3_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14042\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17336\,
            ce => 'H',
            sr => \N__15472\
        );

    \this_vga_signals.M_hcounter_q_0_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7999\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17336\,
            ce => 'H',
            sr => \N__15472\
        );

    \this_vga_signals.M_hcounter_q_RNI84D41_1_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8194\,
            in1 => \N__8257\,
            in2 => \N__8159\,
            in3 => \N__7970\,
            lcout => OPEN,
            ltout => \this_vga_signals.hvisible_i_a2_0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI9JJM1_0_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8217\,
            in2 => \N__7277\,
            in3 => \N__7994\,
            lcout => \this_vga_signals.N_49\,
            ltout => \this_vga_signals.N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7272\,
            in1 => \N__7332\,
            in2 => \N__7235\,
            in3 => \N__8324\,
            lcout => \this_vga_signals.M_hstate_d_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIHS8C_11_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8323\,
            lcout => \this_vga_signals.M_hcounter_q_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7706\,
            in2 => \_gnd_net_\,
            in3 => \N__7427\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17346\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIAU8U1_6_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__8776\,
            in1 => \N__9210\,
            in2 => \N__7361\,
            in3 => \N__8851\,
            lcout => \this_vga_signals.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNID7PV_0_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__7397\,
            in1 => \N__8375\,
            in2 => \_gnd_net_\,
            in3 => \N__8117\,
            lcout => \this_vga_signals.N_26\,
            ltout => \this_vga_signals.N_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIAU8U1_0_6_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__9209\,
            in1 => \N__8847\,
            in2 => \N__7352\,
            in3 => \N__8775\,
            lcout => \this_vga_signals.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8344\,
            in2 => \_gnd_net_\,
            in3 => \N__8328\,
            lcout => \this_vga_signals.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_5_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15508\,
            in2 => \_gnd_net_\,
            in3 => \N__7520\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_1_0_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110101"
        )
    port map (
            in0 => \N__7570\,
            in1 => \_gnd_net_\,
            in2 => \N__7601\,
            in3 => \N__7755\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_RNI3JK8_8_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7597\,
            in2 => \_gnd_net_\,
            in3 => \N__7569\,
            lcout => \this_vga_signals.N_2\,
            ltout => \this_vga_signals.N_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_RNI3BJL_4_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7451\,
            in1 => \N__7756\,
            in2 => \N__7475\,
            in3 => \N__7472\,
            lcout => \this_vga_signals.M_vcounter_q_fast_RNI3BJLZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_RNITCK8_4_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7471\,
            in2 => \_gnd_net_\,
            in3 => \N__7450\,
            lcout => \this_vga_signals.N_70\,
            ltout => \this_vga_signals.N_70_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_RNI61891_7_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7571\,
            in1 => \N__8592\,
            in2 => \N__7460\,
            in3 => \N__8529\,
            lcout => \this_vga_signals.address_1_c5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001000000"
        )
    port map (
            in0 => \N__8524\,
            in1 => \N__7457\,
            in2 => \N__8596\,
            in3 => \N__7923\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_RNIVBOE1_9_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001111111"
        )
    port map (
            in0 => \N__8523\,
            in1 => \N__8583\,
            in2 => \N__8664\,
            in3 => \N__7757\,
            lcout => \this_vga_signals.m44_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_4_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15507\,
            in2 => \_gnd_net_\,
            in3 => \N__7538\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7585\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17710\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQE2J1_9_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8642\,
            in1 => \N__8522\,
            in2 => \N__8433\,
            in3 => \N__7922\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_RNIQE2J1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_RNI27M05_4_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7442\,
            in1 => \N__7815\,
            in2 => \N__7436\,
            in3 => \N__7433\,
            lcout => \this_vga_signals.SUM_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_ac0_3_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000010"
        )
    port map (
            in0 => \N__8587\,
            in1 => \N__8646\,
            in2 => \N__8434\,
            in3 => \N__7490\,
            lcout => \this_vga_signals.mult1_un40_sum_c3\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000110"
        )
    port map (
            in0 => \N__10518\,
            in1 => \N__9002\,
            in2 => \N__7484\,
            in3 => \N__8525\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110011001"
        )
    port map (
            in0 => \N__8648\,
            in1 => \N__8424\,
            in2 => \_gnd_net_\,
            in3 => \N__8588\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__7935\,
            in1 => \_gnd_net_\,
            in2 => \N__7481\,
            in3 => \N__8512\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15506\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7516\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_2_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__8513\,
            in1 => \N__8065\,
            in2 => \_gnd_net_\,
            in3 => \N__7936\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__8066\,
            in1 => \N__7892\,
            in2 => \N__7478\,
            in3 => \N__7877\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_m3_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111000000110"
        )
    port map (
            in0 => \N__8511\,
            in1 => \N__7934\,
            in2 => \N__8665\,
            in3 => \N__7903\,
            lcout => \this_vga_signals.if_i1_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__15505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7534\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNO_0_0_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10813\,
            in2 => \N__7646\,
            in3 => \N__7645\,
            lcout => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNO_0_1_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10922\,
            in2 => \_gnd_net_\,
            in3 => \N__7547\,
            lcout => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNO_0_2_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11030\,
            in2 => \_gnd_net_\,
            in3 => \N__7544\,
            lcout => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNO_0_3_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10734\,
            in2 => \_gnd_net_\,
            in3 => \N__7541\,
            lcout => \this_vga_signals.M_vcounter_q_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7N_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10531\,
            in2 => \_gnd_net_\,
            in3 => \N__7523\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_3_c_RNIVA7NZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8N_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9000\,
            in2 => \_gnd_net_\,
            in3 => \N__7505\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_4_c_RNI1E8NZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15504\,
            in1 => \N__8521\,
            in2 => \_gnd_net_\,
            in3 => \N__7502\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_6\,
            clk => \N__17368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KAN_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8671\,
            in2 => \_gnd_net_\,
            in3 => \N__7499\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_6_c_RNI5KANZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBN_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8597\,
            in2 => \_gnd_net_\,
            in3 => \N__7496\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_7_c_RNI7NBNZ0\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCN_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8435\,
            in2 => \_gnd_net_\,
            in3 => \N__7493\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_RNI9QCNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7998\,
            in2 => \N__7969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_2_c_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8256\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_3_c_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8218\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_4_c_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8193\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_5_c_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8154\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_6_c_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8774\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_7_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7641\,
            in1 => \N__8115\,
            in2 => \_gnd_net_\,
            in3 => \N__7550\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__17324\,
            ce => 'H',
            sr => \N__15470\
        );

    \this_vga_signals.M_hcounter_q_RNIDR6I_8_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__8114\,
            in1 => \N__8370\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.N_27\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_9_c_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8836\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_10_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7640\,
            in1 => \N__9214\,
            in2 => \_gnd_net_\,
            in3 => \N__7649\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_10\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_9\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_10\,
            clk => \N__17329\,
            ce => 'H',
            sr => \N__15468\
        );

    \this_vga_signals.M_hcounter_q_11_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7639\,
            in1 => \N__8329\,
            in2 => \_gnd_net_\,
            in3 => \N__7610\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17329\,
            ce => 'H',
            sr => \N__15468\
        );

    \this_vga_signals.un17_address_g1_0_0_a2_0_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13761\,
            in2 => \_gnd_net_\,
            in3 => \N__12667\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g1_0_0_a2_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13465\,
            in1 => \N__18345\,
            in2 => \N__7607\,
            in3 => \N__13071\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_11_1_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12677\,
            in3 => \N__18346\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_11_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_11_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000110110111"
        )
    port map (
            in0 => \N__13072\,
            in1 => \N__13760\,
            in2 => \N__7604\,
            in3 => \N__13466\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_8_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17685\,
            in2 => \_gnd_net_\,
            in3 => \N__7730\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_7_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7589\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIPD2J1_5_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111111"
        )
    port map (
            in0 => \N__9012\,
            in1 => \N__10539\,
            in2 => \N__7559\,
            in3 => \N__8538\,
            lcout => \this_vga_signals.i9_mux\,
            ltout => \this_vga_signals.i9_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOO3P7_9_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8277\,
            in1 => \N__8426\,
            in2 => \N__7826\,
            in3 => \N__7816\,
            lcout => \this_vga_signals.rgb72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIL6FA3_9_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7823\,
            in1 => \N__8427\,
            in2 => \_gnd_net_\,
            in3 => \N__7817\,
            lcout => port_nmib_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_9_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011100000000"
        )
    port map (
            in0 => \N__9766\,
            in1 => \N__9727\,
            in2 => \N__17712\,
            in3 => \N__7742\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7705\,
            in2 => \_gnd_net_\,
            in3 => \N__7658\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011100000000"
        )
    port map (
            in0 => \N__9765\,
            in1 => \N__9726\,
            in2 => \N__17711\,
            in3 => \N__7741\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_8_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17687\,
            in2 => \_gnd_net_\,
            in3 => \N__7729\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__7704\,
            in1 => \N__7667\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17347\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIAGIO1_5_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__10517\,
            in1 => \N__8647\,
            in2 => \N__9001\,
            in3 => \N__8530\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_1_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNILURK2_9_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8425\,
            in2 => \N__7652\,
            in3 => \N__8589\,
            lcout => \this_vga_signals.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc3_1_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__7858\,
            in1 => \N__8063\,
            in2 => \_gnd_net_\,
            in3 => \N__7846\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un40_sum_axbxc1_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100010000111"
        )
    port map (
            in0 => \N__8531\,
            in1 => \N__7937\,
            in2 => \N__8666\,
            in3 => \N__7904\,
            lcout => \this_vga_signals.mult1_un40_sum_axbxc1\,
            ltout => \this_vga_signals.mult1_un40_sum_axbxc1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101010"
        )
    port map (
            in0 => \N__7886\,
            in1 => \N__8064\,
            in2 => \N__7880\,
            in3 => \N__7876\,
            lcout => \this_vga_signals.mult1_un47_sum_c3\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__9571\,
            in1 => \_gnd_net_\,
            in2 => \N__7865\,
            in3 => \N__11565\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI5CJTF_9_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8067\,
            in1 => \N__8022\,
            in2 => \N__7862\,
            in3 => \N__7847\,
            lcout => \this_vga_signals.address_m1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_1_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__8996\,
            in1 => \N__10522\,
            in2 => \N__10700\,
            in3 => \N__11615\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_3_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100000000"
        )
    port map (
            in0 => \N__15512\,
            in1 => \N__9781\,
            in2 => \N__9725\,
            in3 => \N__7838\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_0_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11614\,
            in1 => \N__8927\,
            in2 => \N__8027\,
            in3 => \N__11564\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_0\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_m24_ns_1_0_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8899\,
            in1 => \N__14348\,
            in2 => \N__7829\,
            in3 => \N__9825\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_m24_ns_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIS78CB9_2_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111011011101"
        )
    port map (
            in0 => \N__10665\,
            in1 => \N__9862\,
            in2 => \N__8078\,
            in3 => \N__11029\,
            lcout => \this_vga_signals.address_i2_mux_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__10519\,
            in1 => \N__8514\,
            in2 => \N__9003\,
            in3 => \N__8071\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c2_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010110010100"
        )
    port map (
            in0 => \N__10521\,
            in1 => \N__11611\,
            in2 => \N__9013\,
            in3 => \N__11562\,
            lcout => \this_vga_signals.mult1_un54_sum_c2\,
            ltout => \this_vga_signals.mult1_un54_sum_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_c3_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100110010000"
        )
    port map (
            in0 => \N__11563\,
            in1 => \N__11613\,
            in2 => \N__8030\,
            in3 => \N__8023\,
            lcout => \this_vga_signals.mult1_un54_sum_c3\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c2_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011101000"
        )
    port map (
            in0 => \N__10664\,
            in1 => \N__10520\,
            in2 => \N__8009\,
            in3 => \N__8898\,
            lcout => \this_vga_signals.mult1_un61_sum_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010011000100"
        )
    port map (
            in0 => \N__15511\,
            in1 => \N__8006\,
            in2 => \N__9731\,
            in3 => \N__9780\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITV8S_2_0_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10669\,
            in2 => \_gnd_net_\,
            in3 => \N__10791\,
            lcout => \this_vga_signals.M_vcounter_q_RNITV8S_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_0_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8000\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \this_vga_signals.un12_address_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7965\,
            in3 => \N__7940\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_0\,
            carryout => \this_vga_signals.un12_address_cry_1\,
            clk => \N__17318\,
            ce => 'H',
            sr => \N__15469\
        );

    \this_vga_signals.un12_address_un12_address_cry_1_c_RNINFAB_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8258\,
            in3 => \N__8225\,
            lcout => \this_vga_signals.un12_address_cry_1_c_RNINFAB\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_1\,
            carryout => \this_vga_signals.un12_address_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_2_c_RNIPIBB_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8222\,
            in3 => \N__8198\,
            lcout => \this_vga_signals.un12_address_cry_2_c_RNIPIBB\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_2\,
            carryout => \this_vga_signals.un12_address_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRLCB_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8195\,
            in3 => \N__8162\,
            lcout => \this_vga_signals.un12_address_cry_3_c_RNIRLCB\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_3\,
            carryout => \this_vga_signals.un12_address_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_4_c_RNITODB_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8158\,
            in3 => \N__8123\,
            lcout => \this_vga_signals.un12_address_cry_4_c_RNITODB\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_4\,
            carryout => \this_vga_signals.un12_address_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_5_c_RNIVREB_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8777\,
            in3 => \N__8120\,
            lcout => \this_vga_signals.un12_address_cry_5_c_RNIVREB\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_5\,
            carryout => \this_vga_signals.un12_address_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_6_c_RNI1VFB_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8116\,
            in3 => \N__8090\,
            lcout => \this_vga_signals.if_m1_0_0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_6\,
            carryout => \this_vga_signals.un12_address_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_7_c_RNI32HB_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8371\,
            in3 => \N__8087\,
            lcout => \this_vga_signals.un12_address_cry_7_c_RNI32HB\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \this_vga_signals.un12_address_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_8_c_RNI55IB_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18650\,
            in2 => \N__8846\,
            in3 => \N__8084\,
            lcout => \this_vga_signals.mult1_un54_sum_axb3_out\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_8\,
            carryout => \this_vga_signals.un12_address_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_cry_9_THRU_LUT4_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9200\,
            in2 => \N__18673\,
            in3 => \N__8081\,
            lcout => \this_vga_signals.un12_address_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un12_address_cry_9\,
            carryout => \this_vga_signals.un12_address_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_10_c_RNINP5K_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9170\,
            in2 => \_gnd_net_\,
            in3 => \N__8378\,
            lcout => \this_vga_signals.un12_address_cry_10_c_RNINP5K\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_8_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10149\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17325\,
            ce => 'H',
            sr => \N__15467\
        );

    \this_vga_signals.M_hcounter_q_RNI3IKE4_11_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__9146\,
            in1 => \N__8348\,
            in2 => \N__8330\,
            in3 => \N__8723\,
            lcout => \N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_1_0_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000111000011"
        )
    port map (
            in0 => \N__12030\,
            in1 => \N__11832\,
            in2 => \N__13452\,
            in3 => \N__10239\,
            lcout => \this_vga_signals.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_2L1_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101100110"
        )
    port map (
            in0 => \N__11833\,
            in1 => \N__12031\,
            in2 => \_gnd_net_\,
            in3 => \N__11760\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axbxc5_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11989\,
            in2 => \N__10244\,
            in3 => \N__11831\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_1_1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011011101"
        )
    port map (
            in0 => \N__10002\,
            in1 => \N__9392\,
            in2 => \_gnd_net_\,
            in3 => \N__9429\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_7_0_3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__10140\,
            in1 => \N__8858\,
            in2 => \N__8261\,
            in3 => \N__9145\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_7_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_7_c_RNI8RAPK_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000011010"
        )
    port map (
            in0 => \N__11834\,
            in1 => \N__9227\,
            in2 => \N__12025\,
            in3 => \N__10141\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_3_2_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000001010"
        )
    port map (
            in0 => \N__9393\,
            in1 => \_gnd_net_\,
            in2 => \N__9434\,
            in3 => \N__10001\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_7_0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIAIMG1_6_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9220\,
            in1 => \N__8852\,
            in2 => \N__8800\,
            in3 => \N__8773\,
            lcout => \this_vga_signals.hvisible_i_a2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_26_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__10243\,
            in1 => \N__12032\,
            in2 => \_gnd_net_\,
            in3 => \N__11847\,
            lcout => \this_vga_signals.g0_6_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7A9S_7_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8670\,
            in2 => \_gnd_net_\,
            in3 => \N__8540\,
            lcout => \this_vga_signals.m30_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI0FV6Q_11_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__16984\,
            in1 => \N__17799\,
            in2 => \N__14500\,
            in3 => \N__17011\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI39IO1_1_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10823\,
            in1 => \N__9014\,
            in2 => \N__10913\,
            in3 => \N__8428\,
            lcout => OPEN,
            ltout => \this_vga_signals.m30_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIEQ4H3_8_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8681\,
            in1 => \N__11026\,
            in2 => \N__8675\,
            in3 => \N__8591\,
            lcout => \this_vga_signals.N_75_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIS0EA1_8_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8672\,
            in1 => \N__8590\,
            in2 => \_gnd_net_\,
            in3 => \N__8539\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIHQRK2_9_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10829\,
            in1 => \N__9008\,
            in2 => \N__8438\,
            in3 => \N__8429\,
            lcout => \this_vga_signals.N_72_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_11_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__19946\,
            in1 => \N__8900\,
            in2 => \_gnd_net_\,
            in3 => \N__9831\,
            lcout => \this_vram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17348\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI0FV6Q_0_11_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__16985\,
            in1 => \N__17798\,
            in2 => \N__14501\,
            in3 => \N__17015\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__9007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11612\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9098\,
            in1 => \N__8897\,
            in2 => \N__9119\,
            in3 => \N__9824\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVOIR1_2_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8933\,
            in1 => \N__11622\,
            in2 => \N__11016\,
            in3 => \N__8926\,
            lcout => \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2\,
            ltout => \this_vga_signals.M_vcounter_q_RNIQVOIR1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI495CI5_2_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9822\,
            in1 => \N__9117\,
            in2 => \N__8915\,
            in3 => \N__8895\,
            lcout => \this_vga_signals.address_i3_mux_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_c3_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111001001101"
        )
    port map (
            in0 => \N__8894\,
            in1 => \N__9113\,
            in2 => \N__8912\,
            in3 => \N__9820\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_m1_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8867\,
            in1 => \N__8896\,
            in2 => \N__8903\,
            in3 => \N__9823\,
            lcout => \this_vga_signals.address_mZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__8893\,
            in1 => \N__9821\,
            in2 => \_gnd_net_\,
            in3 => \N__8866\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c2_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111010100"
        )
    port map (
            in0 => \N__10733\,
            in1 => \N__10986\,
            in2 => \N__9122\,
            in3 => \N__14353\,
            lcout => \this_vga_signals.mult1_un68_sum_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI9MJK5B_2_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011010011111"
        )
    port map (
            in0 => \N__9118\,
            in1 => \N__9097\,
            in2 => \N__9089\,
            in3 => \N__9080\,
            lcout => \this_vga_signals.address_N_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIDN3UA9_3_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111000101"
        )
    port map (
            in0 => \N__10667\,
            in1 => \N__14352\,
            in2 => \N__9635\,
            in3 => \N__14289\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_m27_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI2U4THK_2_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000101110001"
        )
    port map (
            in0 => \N__11002\,
            in1 => \N__9633\,
            in2 => \N__9074\,
            in3 => \N__9527\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_i2_mux_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNICBPF381_2_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__11048\,
            in1 => \N__10856\,
            in2 => \N__9071\,
            in3 => \N__9068\,
            lcout => \this_vga_signals.address_m35_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITV8S_1_0_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10790\,
            in2 => \_gnd_net_\,
            in3 => \N__10666\,
            lcout => \this_vga_signals.M_vcounter_q_RNITV8S_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITV8S_0_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__10668\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10821\,
            lcout => \this_vga_signals.address_m31_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_1_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001100000000"
        )
    port map (
            in0 => \N__9779\,
            in1 => \N__15510\,
            in2 => \N__9724\,
            in3 => \N__9062\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axb4_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101110110110"
        )
    port map (
            in0 => \N__9998\,
            in1 => \N__9424\,
            in2 => \N__9395\,
            in3 => \N__9142\,
            lcout => \this_vga_signals.mult1_un54_sum_axb4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g1_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001010000"
        )
    port map (
            in0 => \N__9143\,
            in1 => \_gnd_net_\,
            in2 => \N__9433\,
            in3 => \N__9390\,
            lcout => \this_vga_signals.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_30_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__13399\,
            in1 => \N__11954\,
            in2 => \_gnd_net_\,
            in3 => \N__10240\,
            lcout => \this_vga_signals.if_m4_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_8_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000001000"
        )
    port map (
            in0 => \N__9997\,
            in1 => \N__9423\,
            in2 => \N__9394\,
            in3 => \N__9141\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_8\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x0_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10128\,
            in1 => \N__9999\,
            in2 => \N__9230\,
            in3 => \N__9919\,
            lcout => \this_vga_signals.mult1_un61_sum_axb4_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g1_1_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001000100"
        )
    port map (
            in0 => \N__9391\,
            in1 => \N__9428\,
            in2 => \_gnd_net_\,
            in3 => \N__9144\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_x1_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10129\,
            in1 => \N__10000\,
            in2 => \_gnd_net_\,
            in3 => \N__9918\,
            lcout => \this_vga_signals.mult1_un61_sum_axb4_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc5_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110000111001"
        )
    port map (
            in0 => \N__9996\,
            in1 => \N__9945\,
            in2 => \N__10150\,
            in3 => \N__9925\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_9_c_RNIEJOE_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9216\,
            in1 => \N__18646\,
            in2 => \_gnd_net_\,
            in3 => \N__9155\,
            lcout => \this_vga_signals.un12_address_cry_9_c_RNIEJOE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g1_2_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__11401\,
            in1 => \N__10042\,
            in2 => \_gnd_net_\,
            in3 => \N__10024\,
            lcout => \this_vga_signals.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_9_c_RNIVF1R_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__9215\,
            in1 => \N__9169\,
            in2 => \_gnd_net_\,
            in3 => \N__9154\,
            lcout => \this_vga_signals.un12_address_cry_9_c_RNIVF1R\,
            ltout => \this_vga_signals.un12_address_cry_9_c_RNIVF1R_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un47_sum_ac0_7_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000101100"
        )
    port map (
            in0 => \N__9995\,
            in1 => \N__9422\,
            in2 => \N__9398\,
            in3 => \N__9383\,
            lcout => \this_vga_signals.mult1_un47_sum_c5\,
            ltout => \this_vga_signals.mult1_un47_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_x1_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110000001"
        )
    port map (
            in0 => \N__10023\,
            in1 => \N__10130\,
            in2 => \N__9359\,
            in3 => \N__12231\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axb3_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb3_ns_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001100110"
        )
    port map (
            in0 => \N__12232\,
            in1 => \N__10158\,
            in2 => \N__9356\,
            in3 => \N__9944\,
            lcout => \this_vga_signals.mult1_un61_sum_axb3\,
            ltout => \this_vga_signals.mult1_un61_sum_axb3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m5_sn_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13349\,
            in2 => \N__9353\,
            in3 => \N__11953\,
            lcout => \this_vga_signals.if_m5_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m5_rn_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111010"
        )
    port map (
            in0 => \N__13400\,
            in1 => \_gnd_net_\,
            in2 => \N__12034\,
            in3 => \N__10235\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m5_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m5_mb_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__11724\,
            in1 => \N__9350\,
            in2 => \N__9344\,
            in3 => \N__11835\,
            lcout => \this_vga_signals.mult1_un68_sum_c5\,
            ltout => \this_vga_signals.mult1_un68_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axb3_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13401\,
            in1 => \N__12589\,
            in2 => \N__9341\,
            in3 => \N__18310\,
            lcout => \this_vga_signals.mult1_un75_sum_axb3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_c4_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111011"
        )
    port map (
            in0 => \N__10142\,
            in1 => \N__10011\,
            in2 => \_gnd_net_\,
            in3 => \N__9920\,
            lcout => \this_vga_signals.mult1_un54_sum_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIAFTT93_9_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__12637\,
            in1 => \N__18311\,
            in2 => \N__19985\,
            in3 => \N__13062\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_axbxc3_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10143\,
            in1 => \N__10012\,
            in2 => \_gnd_net_\,
            in3 => \N__9921\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_7_0_4_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011011100"
        )
    port map (
            in0 => \N__9950\,
            in1 => \N__9458\,
            in2 => \N__9452\,
            in3 => \N__9449\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_7_0_4\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_7_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m1_0_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110000"
        )
    port map (
            in0 => \N__10234\,
            in1 => \_gnd_net_\,
            in2 => \N__9443\,
            in3 => \N__12017\,
            lcout => \this_vga_signals.if_m1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_i_o2_0_x2_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__13042\,
            in1 => \N__11851\,
            in2 => \N__11761\,
            in3 => \N__12675\,
            lcout => \this_vga_signals.N_26_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m4_0_1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__13402\,
            in1 => \N__11993\,
            in2 => \_gnd_net_\,
            in3 => \N__10241\,
            lcout => \this_vga_signals.if_m4_0_1\,
            ltout => \this_vga_signals.if_m4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_25_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011100000"
        )
    port map (
            in0 => \N__11755\,
            in1 => \N__11852\,
            in2 => \N__9440\,
            in3 => \N__11995\,
            lcout => \this_vga_signals.if_N_8_mux_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_6_c_RNIGPBEN_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000111100"
        )
    port map (
            in0 => \N__11994\,
            in1 => \N__11839\,
            in2 => \N__13451\,
            in3 => \N__10242\,
            lcout => \this_vga_signals.G_12_0_x3_0\,
            ltout => \this_vga_signals.G_12_0_x3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_3_c_RNI913733_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__13043\,
            in1 => \N__12907\,
            in2 => \N__9437\,
            in3 => \N__13300\,
            lcout => \this_vga_signals.G_12_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_38_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12651\,
            in2 => \N__18348\,
            in3 => \N__13041\,
            lcout => \this_vga_signals.g0_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_2_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__11996\,
            in1 => \N__11840\,
            in2 => \N__12945\,
            in3 => \N__11756\,
            lcout => \this_vga_signals.g0_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNITHP2_0_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10571\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9602\,
            lcout => vsync_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_0_1_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__9600\,
            in1 => \N__9764\,
            in2 => \_gnd_net_\,
            in3 => \N__9488\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_1_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001110"
        )
    port map (
            in0 => \N__10469\,
            in1 => \N__9601\,
            in2 => \N__9491\,
            in3 => \N__17709\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIEQ4H3_1_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9479\,
            in1 => \N__10904\,
            in2 => \_gnd_net_\,
            in3 => \N__11027\,
            lcout => \this_vga_signals.N_76_mux\,
            ltout => \this_vga_signals.N_76_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_2_0_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__9763\,
            in1 => \N__9598\,
            in2 => \N__9482\,
            in3 => \N__10743\,
            lcout => \this_vga_signals.M_vstate_q_RNO_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_3_0_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__9478\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10903\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_1_0_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111101111"
        )
    port map (
            in0 => \N__11028\,
            in1 => \N__9599\,
            in2 => \N__9470\,
            in3 => \N__10742\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vstate_q_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_0_0_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10570\,
            in2 => \N__9467\,
            in3 => \N__9464\,
            lcout => \this_vga_signals.N_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI149S_4_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10538\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10739\,
            lcout => OPEN,
            ltout => \this_vga_signals.m35_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNI4LE61_0_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9597\,
            in1 => \N__10567\,
            in2 => \N__9578\,
            in3 => \N__15503\,
            lcout => \this_vga_signals.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14285\,
            in1 => \N__9560\,
            in2 => \N__9551\,
            in3 => \N__14357\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIV7VFA9_0_2_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010001100001"
        )
    port map (
            in0 => \N__11023\,
            in1 => \N__14351\,
            in2 => \N__10748\,
            in3 => \N__14284\,
            lcout => \this_vga_signals.address_N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_0_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9575\,
            in1 => \N__11623\,
            in2 => \N__10545\,
            in3 => \N__11572\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9833\,
            in1 => \N__10732\,
            in2 => \_gnd_net_\,
            in3 => \N__9842\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc1\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_c3_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100110010000"
        )
    port map (
            in0 => \N__14288\,
            in1 => \N__14358\,
            in2 => \N__9554\,
            in3 => \N__9550\,
            lcout => \this_vga_signals.mult1_un68_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIV7VFA9_1_2_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000011000"
        )
    port map (
            in0 => \N__10992\,
            in1 => \N__14349\,
            in2 => \N__10735\,
            in3 => \N__14286\,
            lcout => \this_vga_signals.address_N_9_0\,
            ltout => \this_vga_signals.address_N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_0_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__10828\,
            in1 => \_gnd_net_\,
            in2 => \N__9536\,
            in3 => \N__9533\,
            lcout => \this_vga_signals.address_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI8OSG6B_2_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__10993\,
            in1 => \N__10731\,
            in2 => \_gnd_net_\,
            in3 => \N__9526\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_RNI8OSG6BZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI5UR0HK_2_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9866\,
            in2 => \N__9845\,
            in3 => \N__10339\,
            lcout => \this_vga_signals.address_i2_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10864\,
            in1 => \N__14350\,
            in2 => \_gnd_net_\,
            in3 => \N__14287\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9841\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9832\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI4G7F3B2_0_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__9641\,
            in1 => \N__9608\,
            in2 => \N__10871\,
            in3 => \N__9788\,
            lcout => \this_vga_signals.address_N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_2_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100000000"
        )
    port map (
            in0 => \N__15509\,
            in1 => \N__9782\,
            in2 => \N__9709\,
            in3 => \N__9662\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17353\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI9MCQB9_2_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000101111"
        )
    port map (
            in0 => \N__10619\,
            in1 => \N__10998\,
            in2 => \N__9650\,
            in3 => \N__10334\,
            lcout => \this_vga_signals.address_i2_mux_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIS78CB9_0_2_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100111000"
        )
    port map (
            in0 => \N__10335\,
            in1 => \N__9634\,
            in2 => \N__11024\,
            in3 => \N__10747\,
            lcout => \this_vga_signals.address_i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIV7VFA9_2_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101100110"
        )
    port map (
            in0 => \N__10746\,
            in1 => \N__10997\,
            in2 => \_gnd_net_\,
            in3 => \N__10333\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIBU2ELI_0_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__9617\,
            in1 => \_gnd_net_\,
            in2 => \N__9611\,
            in3 => \N__10822\,
            lcout => \this_vga_signals.address_N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_4_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111101100"
        )
    port map (
            in0 => \N__10028\,
            in1 => \N__11394\,
            in2 => \N__10058\,
            in3 => \N__10165\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axb3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_4_0_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100001000"
        )
    port map (
            in0 => \N__12023\,
            in1 => \N__10310\,
            in2 => \N__10049\,
            in3 => \N__11864\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_4_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13449\,
            in1 => \N__12628\,
            in2 => \N__10046\,
            in3 => \N__13083\,
            lcout => \this_vga_signals.g0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_2_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001011010"
        )
    port map (
            in0 => \N__11393\,
            in1 => \N__10027\,
            in2 => \N__10166\,
            in3 => \N__10043\,
            lcout => \this_vga_signals.mult1_un61_sum_axb3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un54_sum_ac0_7_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000100"
        )
    port map (
            in0 => \N__10026\,
            in1 => \N__9946\,
            in2 => \N__9926\,
            in3 => \N__10161\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_7\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_axb4_ns_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9893\,
            in2 => \N__9887\,
            in3 => \N__9884\,
            lcout => \this_vga_signals.mult1_un61_sum_axb4_i\,
            ltout => \this_vga_signals.mult1_un61_sum_axb4_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m2_3_0_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9878\,
            in3 => \N__10222\,
            lcout => \this_vga_signals.if_m2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un61_sum_ac0_5_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12000\,
            in2 => \_gnd_net_\,
            in3 => \N__10223\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_5\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000001011"
        )
    port map (
            in0 => \N__10159\,
            in1 => \N__10174\,
            in2 => \N__9875\,
            in3 => \N__9872\,
            lcout => this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0,
            ltout => \this_vga_signals_un17_address_if_generate_plus_mult1_un68_sum_axbxc5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_0_a2_1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10259\,
            in1 => \N__12832\,
            in2 => \N__10247\,
            in3 => \N__12806\,
            lcout => \this_vga_signals.g0_0_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_21_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010000"
        )
    port map (
            in0 => \N__10224\,
            in1 => \_gnd_net_\,
            in2 => \N__12029\,
            in3 => \N__11845\,
            lcout => \this_vga_signals.g0_6_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_41_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__12012\,
            in1 => \N__13471\,
            in2 => \_gnd_net_\,
            in3 => \N__10225\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m4_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_15_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101000"
        )
    port map (
            in0 => \N__11723\,
            in1 => \N__12013\,
            in2 => \N__10178\,
            in3 => \N__11846\,
            lcout => \this_vga_signals.if_N_8_mux_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m2_3_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111010010"
        )
    port map (
            in0 => \N__10175\,
            in1 => \N__10160\,
            in2 => \N__10082\,
            in3 => \N__11722\,
            lcout => \this_vga_signals.if_N_3_3_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_6_1_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__13470\,
            in1 => \N__10073\,
            in2 => \_gnd_net_\,
            in3 => \N__11844\,
            lcout => \this_vga_signals.g0_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_16_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__11728\,
            in1 => \N__11837\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.N_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_0_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000101100100"
        )
    port map (
            in0 => \N__12600\,
            in1 => \N__12315\,
            in2 => \N__13802\,
            in3 => \N__12805\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_3_c_RNIKCM73C_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__10292\,
            in1 => \N__10067\,
            in2 => \N__10061\,
            in3 => \N__13288\,
            lcout => OPEN,
            ltout => \this_vga_signals.G_12_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_3_c_RNIRBMU931_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__13554\,
            in1 => \N__10283\,
            in2 => \N__10313\,
            in3 => \N__10583\,
            lcout => \this_vga_signals.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m4_0_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101000"
        )
    port map (
            in0 => \N__12021\,
            in1 => \N__11836\,
            in2 => \N__11747\,
            in3 => \N__10306\,
            lcout => \this_vga_signals_un17_address_if_N_8_mux\,
            ltout => \this_vga_signals_un17_address_if_N_8_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_4_c_RNIU8UQ04_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010001001010"
        )
    port map (
            in0 => \N__12599\,
            in1 => \N__13748\,
            in2 => \N__10295\,
            in3 => \N__12804\,
            lcout => \this_vga_signals.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_i_x4_4_a3_1_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__12022\,
            in1 => \N__13553\,
            in2 => \N__11748\,
            in3 => \N__11838\,
            lcout => \this_vga_signals.g0_i_x4_4_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g1_2_0_a2_0_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12650\,
            in3 => \N__13035\,
            lcout => \this_vga_signals.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \G_12_0_x2_0_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12308\,
            in1 => \N__12794\,
            in2 => \_gnd_net_\,
            in3 => \N__13281\,
            lcout => OPEN,
            ltout => \N_6_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_4_c_RNID4564B_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__10592\,
            in1 => \N__13773\,
            in2 => \N__10286\,
            in3 => \N__13552\,
            lcout => \this_vga_signals.N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_6_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__10274\,
            in1 => \N__12795\,
            in2 => \N__12035\,
            in3 => \N__13045\,
            lcout => \this_vga_signals.g0_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_6_c_RNIHI8G23_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10265\,
            in1 => \N__12652\,
            in2 => \_gnd_net_\,
            in3 => \N__13044\,
            lcout => \this_vga_signals.N_5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \G_12_0_o7_1_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100101100000"
        )
    port map (
            in0 => \N__12796\,
            in1 => \N__12309\,
            in2 => \N__12674\,
            in3 => \N__13282\,
            lcout => OPEN,
            ltout => \N_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_3_c_RNIPAA128_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011101100"
        )
    port map (
            in0 => \N__12950\,
            in1 => \N__13772\,
            in2 => \N__10595\,
            in3 => \N__10591\,
            lcout => \this_vga_signals.G_12_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_0_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001101"
        )
    port map (
            in0 => \N__10547\,
            in1 => \N__10569\,
            in2 => \N__17727\,
            in3 => \N__10577\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNO_1_1_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10568\,
            in1 => \N__10744\,
            in2 => \_gnd_net_\,
            in3 => \N__10546\,
            lcout => \this_vga_signals.N_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_m16_0_x4_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10741\,
            in1 => \N__14368\,
            in2 => \_gnd_net_\,
            in3 => \N__14300\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_9_i_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101011100"
        )
    port map (
            in0 => \N__11025\,
            in1 => \N__10835\,
            in2 => \N__10463\,
            in3 => \N__10460\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIO5SOPF2_9_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__19986\,
            in1 => \N__11524\,
            in2 => \N__10454\,
            in3 => \N__11539\,
            lcout => \M_this_vga_signals_address_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITV8S_3_0_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10827\,
            in2 => \_gnd_net_\,
            in3 => \N__10740\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_m6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI9MCQB9_0_2_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111001100"
        )
    port map (
            in0 => \N__10615\,
            in1 => \N__11004\,
            in2 => \N__10343\,
            in3 => \N__10340\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI2QRE761_0_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__11046\,
            in1 => \N__10868\,
            in2 => \N__11189\,
            in3 => \N__11186\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_m21_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7GUI2B2_2_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__10870\,
            in1 => \N__11180\,
            in2 => \N__11174\,
            in3 => \N__11171\,
            lcout => OPEN,
            ltout => \this_vga_signals.address_N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIH8E9EM_1_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__10917\,
            in1 => \N__20008\,
            in2 => \N__11165\,
            in3 => \N__11162\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_address_if_m16_0_o4_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011010100"
        )
    port map (
            in0 => \N__11047\,
            in1 => \N__11003\,
            in2 => \N__10921\,
            in3 => \N__10869\,
            lcout => \this_vga_signals.if_m16_0_o4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNITV8S_0_0_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10745\,
            lcout => \this_vga_signals.address_N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_20_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__13082\,
            in1 => \_gnd_net_\,
            in2 => \N__12661\,
            in3 => \N__18355\,
            lcout => \this_vga_signals.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_14_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001000"
        )
    port map (
            in0 => \N__11743\,
            in1 => \N__12024\,
            in2 => \N__11870\,
            in3 => \N__10604\,
            lcout => \this_vga_signals.if_N_8_mux_2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_3L3_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12620\,
            in2 => \N__18361\,
            in3 => \N__13081\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_3L3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_N_4L5_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100111110011"
        )
    port map (
            in0 => \N__13709\,
            in1 => \N__13448\,
            in2 => \N__11234\,
            in3 => \N__12481\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5\,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4L5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11231\,
            in2 => \N__11219\,
            in3 => \N__13575\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc5_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_10_i_o2_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11865\,
            in2 => \_gnd_net_\,
            in3 => \N__11742\,
            lcout => \this_vga_signals.N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_16_0_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__13478\,
            in1 => \N__11881\,
            in2 => \N__13816\,
            in3 => \N__11678\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_3_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11216\,
            in1 => \N__13283\,
            in2 => \N__13488\,
            in3 => \N__13084\,
            lcout => \this_vga_signals.g0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_9_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12799\,
            in1 => \N__12314\,
            in2 => \_gnd_net_\,
            in3 => \N__12626\,
            lcout => \this_vga_signals.N_20_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_0_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12625\,
            in1 => \N__12798\,
            in2 => \N__11210\,
            in3 => \N__11198\,
            lcout => \this_vga_signals.g0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_22_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12797\,
            in1 => \N__12313\,
            in2 => \N__13823\,
            in3 => \N__12624\,
            lcout => \this_vga_signals.N_3_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_axb3_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12627\,
            in1 => \N__12800\,
            in2 => \N__13817\,
            in3 => \N__12316\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axb3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__12980\,
            in1 => \N__12401\,
            in2 => \N__11192\,
            in3 => \N__12713\,
            lcout => \this_vga_signals.mult1_un82_sum_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_i_x4_4_a3_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__11375\,
            in1 => \N__11369\,
            in2 => \N__11654\,
            in3 => \N__12041\,
            lcout => \this_vga_signals.g0_i_x4_4_a3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m5_2_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001100010"
        )
    port map (
            in0 => \N__11363\,
            in1 => \N__13463\,
            in2 => \N__13784\,
            in3 => \N__11354\,
            lcout => this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5,
            ltout => \this_vga_signals_un17_address_if_generate_plus_mult1_un75_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un75_sum_axbxc5_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12602\,
            in2 => \N__11348\,
            in3 => \N__12298\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m2_2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12299\,
            in1 => \N__13271\,
            in2 => \N__12814\,
            in3 => \N__12465\,
            lcout => \this_vga_signals.if_N_3_2_i\,
            ltout => \this_vga_signals.if_N_3_2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_generate_plus_mult1_un82_sum_ac0_7_0_1_0_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001100110"
        )
    port map (
            in0 => \N__12466\,
            in1 => \N__13733\,
            in2 => \N__11345\,
            in3 => \N__13574\,
            lcout => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_2_0_a3_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13464\,
            in1 => \N__18347\,
            in2 => \N__13785\,
            in3 => \N__11676\,
            lcout => \this_vga_signals.g1_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_if_m2_2_0_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13729\,
            in2 => \_gnd_net_\,
            in3 => \N__12601\,
            lcout => this_vga_signals_un17_address_if_m2_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIP8K884_9_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__12603\,
            in1 => \N__12317\,
            in2 => \N__20012\,
            in3 => \N__12812\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g1_0_0_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__13771\,
            in1 => \N__12660\,
            in2 => \N__12978\,
            in3 => \N__13189\,
            lcout => \this_vga_signals.g1_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_0_a2_2_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011010101001"
        )
    port map (
            in0 => \N__13453\,
            in1 => \N__11869\,
            in2 => \N__11762\,
            in3 => \N__12302\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_0_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_12_0_a3_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12790\,
            in1 => \N__11677\,
            in2 => \N__11660\,
            in3 => \N__13278\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_3_2_i_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_0_a2_3_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__13769\,
            in1 => \N__12949\,
            in2 => \N__11657\,
            in3 => \N__11645\,
            lcout => \this_vga_signals.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_14_0_a2_i_x2_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__12301\,
            in1 => \_gnd_net_\,
            in2 => \N__12813\,
            in3 => \N__12659\,
            lcout => \this_vga_signals.N_20_i_i\,
            ltout => \this_vga_signals.N_20_i_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_a3_3_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100101101"
        )
    port map (
            in0 => \N__13454\,
            in1 => \N__13770\,
            in2 => \N__11639\,
            in3 => \N__11636\,
            lcout => \this_vga_signals.g0_0_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_2_2_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12300\,
            in2 => \_gnd_net_\,
            in3 => \N__12786\,
            lcout => \this_vga_signals.N_4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_12_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__19995\,
            in1 => \N__11627\,
            in2 => \_gnd_net_\,
            in3 => \N__11576\,
            lcout => \this_vram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIL305C61_9_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__11540\,
            in1 => \N__19993\,
            in2 => \_gnd_net_\,
            in3 => \N__11525\,
            lcout => \M_this_vga_signals_address_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIR6TCF_9_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__19994\,
            in1 => \N__11405\,
            in2 => \_gnd_net_\,
            in3 => \N__12242\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_17_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011101110111"
        )
    port map (
            in0 => \N__13450\,
            in1 => \N__12107\,
            in2 => \N__13814\,
            in3 => \N__12485\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIETEJ4_11_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16977\,
            in1 => \N__17830\,
            in2 => \_gnd_net_\,
            in3 => \N__16999\,
            lcout => OPEN,
            ltout => \this_vram.M_this_vram_read_data_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI0FV6Q_1_11_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__14141\,
            in1 => \_gnd_net_\,
            in2 => \N__12101\,
            in3 => \N__16952\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_6_0_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19825\,
            in1 => \N__13298\,
            in2 => \N__12071\,
            in3 => \N__12815\,
            lcout => \this_vga_signals.g0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_5_0_a2_0_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12059\,
            in1 => \N__12663\,
            in2 => \N__13820\,
            in3 => \N__12808\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_3_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_5_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010110000101"
        )
    port map (
            in0 => \N__12976\,
            in1 => \N__14050\,
            in2 => \N__12050\,
            in3 => \N__12347\,
            lcout => \this_vga_signals.mult1_un89_sum_c5_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_0_0_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__13555\,
            in1 => \N__12047\,
            in2 => \N__13818\,
            in3 => \N__12710\,
            lcout => \this_vga_signals.g0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_a3_2_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12033\,
            in1 => \N__11882\,
            in2 => \N__12987\,
            in3 => \N__13556\,
            lcout => \this_vga_signals.g0_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_13_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12323\,
            in1 => \N__12662\,
            in2 => \N__13819\,
            in3 => \N__12807\,
            lcout => \this_vga_signals.g0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111101111"
        )
    port map (
            in0 => \N__12422\,
            in1 => \N__13798\,
            in2 => \N__12988\,
            in3 => \N__12416\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_a3_5_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101001100101"
        )
    port map (
            in0 => \N__12410\,
            in1 => \N__12400\,
            in2 => \N__12389\,
            in3 => \N__12386\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_a3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_a3_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000101101"
        )
    port map (
            in0 => \N__12975\,
            in1 => \N__14051\,
            in2 => \N__12380\,
            in3 => \N__12377\,
            lcout => \this_vga_signals.mult1_un96_sum_axbxc5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_29_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12957\,
            in1 => \N__12371\,
            in2 => \_gnd_net_\,
            in3 => \N__13135\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_5_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_27_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__12365\,
            in1 => \N__12356\,
            in2 => \N__12350\,
            in3 => \N__12842\,
            lcout => \this_vga_signals.r_N_2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_1_2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12318\,
            in1 => \N__12671\,
            in2 => \N__12341\,
            in3 => \N__13076\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_12_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13279\,
            in2 => \N__12326\,
            in3 => \N__12801\,
            lcout => \this_vga_signals.if_N_3_2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_3_0_a2_1_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12319\,
            in1 => \N__18356\,
            in2 => \N__13489\,
            in3 => \N__13077\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_3_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_3_0_a2_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12672\,
            in1 => \N__13280\,
            in2 => \N__12845\,
            in3 => \N__12802\,
            lcout => \this_vga_signals.if_N_3_2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_23_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011000000110"
        )
    port map (
            in0 => \N__13813\,
            in1 => \N__12482\,
            in2 => \N__13576\,
            in3 => \N__12711\,
            lcout => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_5_0_a2_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12673\,
            in1 => \N__12836\,
            in2 => \N__13822\,
            in3 => \N__12803\,
            lcout => \this_vga_signals.N_3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_37_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011000000110"
        )
    port map (
            in0 => \N__13774\,
            in1 => \N__12483\,
            in2 => \N__13577\,
            in3 => \N__12712\,
            lcout => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_5_c_RNI8HPEH2_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12689\,
            in1 => \N__13287\,
            in2 => \N__13490\,
            in3 => \N__12676\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_5_c_RNICKLJPG_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13564\,
            in1 => \N__12509\,
            in2 => \N__12500\,
            in3 => \N__12497\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_3_c_RNI5J0QQK_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111010010"
        )
    port map (
            in0 => \N__12979\,
            in1 => \N__13776\,
            in2 => \N__12488\,
            in3 => \N__13565\,
            lcout => \this_vga_signals.g1_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_36_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011100111111"
        )
    port map (
            in0 => \N__13775\,
            in1 => \N__13482\,
            in2 => \N__13211\,
            in3 => \N__12484\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc5_1_N_4_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_3_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12434\,
            in2 => \N__12425\,
            in3 => \N__13563\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_33_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111000"
        )
    port map (
            in0 => \N__13175\,
            in1 => \N__13163\,
            in2 => \N__13157\,
            in3 => \N__13154\,
            lcout => \this_vga_signals.N_3_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_5_0_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13777\,
            in2 => \_gnd_net_\,
            in3 => \N__13447\,
            lcout => \this_vga_signals.g0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_7_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100110011100"
        )
    port map (
            in0 => \N__13815\,
            in1 => \N__13148\,
            in2 => \N__12989\,
            in3 => \N__13583\,
            lcout => \this_vga_signals.g0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g1_4_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__12981\,
            in1 => \N__13142\,
            in2 => \_gnd_net_\,
            in3 => \N__13136\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_0_0_a2_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110010110"
        )
    port map (
            in0 => \N__13124\,
            in1 => \N__13115\,
            in2 => \N__13109\,
            in3 => \N__13496\,
            lcout => OPEN,
            ltout => \this_vga_signals.r_N_2_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_10_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100000110011"
        )
    port map (
            in0 => \N__14049\,
            in1 => \N__12986\,
            in2 => \N__13106\,
            in3 => \N__13103\,
            lcout => \this_vga_signals.mult1_un89_sum_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_5_3_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18357\,
            in1 => \N__13299\,
            in2 => \N__13097\,
            in3 => \N__13085\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_34_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110110110100"
        )
    port map (
            in0 => \N__13806\,
            in1 => \N__12982\,
            in2 => \N__12848\,
            in3 => \N__13579\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un96_sum_c5_0_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_32_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111101000"
        )
    port map (
            in0 => \N__14048\,
            in1 => \N__14008\,
            in2 => \N__13991\,
            in3 => \N__13988\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un96_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un12_address_un12_address_cry_3_c_RNI7M4QI33_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__13982\,
            in1 => \_gnd_net_\,
            in2 => \N__13976\,
            in3 => \N__13973\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIHKRBFB2_9_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__13964\,
            in1 => \N__19999\,
            in2 => \N__13958\,
            in3 => \N__13955\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_24_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__13841\,
            in1 => \N__13829\,
            in2 => \N__13821\,
            in3 => \N__13578\,
            lcout => \this_vga_signals.mult1_un82_sum_ac0_7_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un17_address_g0_35_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13487\,
            in1 => \N__13301\,
            in2 => \N__13210\,
            in3 => \N__13190\,
            lcout => \this_vga_signals.if_N_3_2_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_1_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13169\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_0_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14122\,
            in1 => \N__16887\,
            in2 => \_gnd_net_\,
            in3 => \N__14105\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_1_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14093\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_last_q_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16895\,
            lcout => \this_start_data_delay_this_edge_detector_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_0_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__14131\,
            in1 => \N__16894\,
            in2 => \_gnd_net_\,
            in3 => \N__14104\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_4_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14087\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_3_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14075\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_2_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14081\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_6_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14069\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_5_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14405\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_3_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14057\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_2_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14063\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_4_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14411\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_10_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14393\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_11_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14399\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17319\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_9_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14540\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_6_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14375\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_7_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14387\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_5_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14381\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOUPCH9_9_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__20019\,
            in1 => \N__14369\,
            in2 => \_gnd_net_\,
            in3 => \N__14299\,
            lcout => \M_this_vga_signals_address_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIETEJ4_0_11_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18716\,
            in1 => \N__17841\,
            in2 => \_gnd_net_\,
            in3 => \N__18079\,
            lcout => \this_vram.M_this_vram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIIHGJL_11_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__18080\,
            in1 => \N__17837\,
            in2 => \N__16951\,
            in3 => \N__18709\,
            lcout => \this_vram.N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_12_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14465\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_13_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14459\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_state_q_s2_0_a3_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__17503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16355\,
            lcout => debug_d,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_16_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14423\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_14_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14435\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_15_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14429\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_5_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__14949\,
            in1 => \N__17567\,
            in2 => \N__14753\,
            in3 => \N__16339\,
            lcout => \this_start_data_delay.this_edge_detector.N_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_17_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_19_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14552\,
            lcout => \M_this_start_data_delay_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_18_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14558\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_delay.M_pipe_q_8_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14546\,
            lcout => \this_start_data_delay.this_delay.M_pipe_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_2_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__16343\,
            in1 => \N__14567\,
            in2 => \N__14522\,
            in3 => \N__17500\,
            lcout => \M_current_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17338\,
            ce => 'H',
            sr => \N__15464\
        );

    \M_current_address_q_5_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__17499\,
            in1 => \N__14924\,
            in2 => \N__14534\,
            in3 => \N__16344\,
            lcout => \M_current_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17338\,
            ce => 'H',
            sr => \N__15464\
        );

    \M_current_address_q_9_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__14774\,
            in1 => \N__17486\,
            in2 => \N__14510\,
            in3 => \N__16342\,
            lcout => \M_current_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17342\,
            ce => 'H',
            sr => \N__15462\
        );

    \M_current_address_q_8_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110101001000"
        )
    port map (
            in0 => \N__16341\,
            in1 => \N__16022\,
            in2 => \N__17501\,
            in3 => \N__14909\,
            lcout => \M_current_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17342\,
            ce => 'H',
            sr => \N__15462\
        );

    \M_current_address_q_4_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__15059\,
            in1 => \N__17485\,
            in2 => \N__16370\,
            in3 => \N__16340\,
            lcout => \M_current_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17342\,
            ce => 'H',
            sr => \N__15462\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_2_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__14593\,
            in1 => \N__17604\,
            in2 => \N__19036\,
            in3 => \N__16333\,
            lcout => \this_start_data_delay.this_edge_detector.N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_9_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__14800\,
            in1 => \N__17605\,
            in2 => \N__19037\,
            in3 => \N__16334\,
            lcout => \this_start_data_delay.this_edge_detector.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_12_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__15131\,
            in1 => \N__17502\,
            in2 => \N__14723\,
            in3 => \N__16351\,
            lcout => \M_current_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17328\,
            ce => 'H',
            sr => \N__15466\
        );

    \this_start_address_delay.this_delay.M_pipe_q_9_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_8_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14702\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_12_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__19273\,
            in1 => \N__17568\,
            in2 => \N__14752\,
            in3 => \N__16338\,
            lcout => \this_start_data_delay.this_edge_detector.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_7_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14714\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_10_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14696\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNIHDTU_0_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15583\,
            in2 => \N__15116\,
            in3 => \N__15115\,
            lcout => \M_current_address_q_RNIHDTUZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_19_23_0_\,
            carryout => \un1_M_current_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_0_c_RNI2QAN_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16567\,
            in2 => \_gnd_net_\,
            in3 => \N__14690\,
            lcout => \un1_M_current_address_q_cry_0_c_RNI2QANZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_0\,
            carryout => \un1_M_current_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_1_c_RNI4TBN_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14589\,
            in2 => \_gnd_net_\,
            in3 => \N__14561\,
            lcout => \un1_M_current_address_q_cry_1_c_RNI4TBNZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_1\,
            carryout => \un1_M_current_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_2_c_RNI60DN_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15160\,
            in2 => \_gnd_net_\,
            in3 => \N__15062\,
            lcout => \un1_M_current_address_q_cry_2_c_RNI60DNZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_2\,
            carryout => \un1_M_current_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_3_c_RNI83EN_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16422\,
            in2 => \_gnd_net_\,
            in3 => \N__15053\,
            lcout => \un1_M_current_address_q_cry_3_c_RNI83ENZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_3\,
            carryout => \un1_M_current_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_4_c_RNIA6FN_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14950\,
            in2 => \_gnd_net_\,
            in3 => \N__14918\,
            lcout => \un1_M_current_address_q_cry_4_c_RNIA6FNZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_4\,
            carryout => \un1_M_current_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_5_c_RNIC9GN_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15289\,
            in2 => \_gnd_net_\,
            in3 => \N__14915\,
            lcout => \un1_M_current_address_q_cry_5_c_RNIC9GNZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_5\,
            carryout => \un1_M_current_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_6_c_RNIECHN_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15714\,
            in2 => \_gnd_net_\,
            in3 => \N__14912\,
            lcout => \un1_M_current_address_q_cry_6_c_RNIECHNZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_6\,
            carryout => \un1_M_current_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_7_c_RNIGFIN_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16041\,
            in2 => \_gnd_net_\,
            in3 => \N__14903\,
            lcout => \un1_M_current_address_q_cry_7_c_RNIGFINZ0\,
            ltout => OPEN,
            carryin => \bfn_19_24_0_\,
            carryout => \un1_M_current_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_8_c_RNIIIJN_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14799\,
            in2 => \_gnd_net_\,
            in3 => \N__14768\,
            lcout => \un1_M_current_address_q_cry_8_c_RNIIIJNZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_8\,
            carryout => \un1_M_current_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_9_c_RNIRDIM_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15909\,
            in2 => \_gnd_net_\,
            in3 => \N__14765\,
            lcout => \un1_M_current_address_q_cry_9_c_RNIRDIMZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_9\,
            carryout => \un1_M_current_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_10_c_RNI4KKH_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19185\,
            in2 => \_gnd_net_\,
            in3 => \N__14762\,
            lcout => \un1_M_current_address_q_cry_10_c_RNI4KKHZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_10\,
            carryout => \un1_M_current_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_11_c_RNI6NLH_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19286\,
            in2 => \_gnd_net_\,
            in3 => \N__15122\,
            lcout => \un1_M_current_address_q_cry_11_c_RNI6NLHZ0\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_11\,
            carryout => \un1_M_current_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_current_address_q_cry_12_c_RNI8QMH_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19082\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15119\,
            lcout => \un1_M_current_address_q_cry_12_c_RNI8QMHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.un1_M_state_q_1_i_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111001100"
        )
    port map (
            in0 => \N__17608\,
            in1 => \N__17484\,
            in2 => \_gnd_net_\,
            in3 => \N__16296\,
            lcout => \N_177_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_10_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__15101\,
            in1 => \N__17481\,
            in2 => \N__15890\,
            in3 => \N__16335\,
            lcout => \M_current_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17354\,
            ce => 'H',
            sr => \N__15463\
        );

    \M_current_address_q_1_LC_19_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__16337\,
            in1 => \N__15095\,
            in2 => \N__16541\,
            in3 => \N__17483\,
            lcout => \M_current_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17354\,
            ce => 'H',
            sr => \N__15463\
        );

    \M_current_address_q_13_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__16336\,
            in1 => \N__17482\,
            in2 => \N__15842\,
            in3 => \N__15086\,
            lcout => \M_current_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17354\,
            ce => 'H',
            sr => \N__15463\
        );

    \this_start_address_delay.this_delay.M_pipe_q_13_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15080\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_12_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15068\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_11_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15074\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_15_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15548\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_14_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15554\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_0_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__17477\,
            in1 => \N__15542\,
            in2 => \N__15563\,
            in3 => \N__16291\,
            lcout => \M_current_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17349\,
            ce => 'H',
            sr => \N__15465\
        );

    \M_current_address_q_6_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110101001000"
        )
    port map (
            in0 => \N__16294\,
            in1 => \N__15269\,
            in2 => \N__17504\,
            in3 => \N__15536\,
            lcout => \M_current_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17349\,
            ce => 'H',
            sr => \N__15465\
        );

    \M_current_address_q_7_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__16295\,
            in1 => \N__15530\,
            in2 => \N__15695\,
            in3 => \N__17480\,
            lcout => \M_current_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17349\,
            ce => 'H',
            sr => \N__15465\
        );

    \M_current_address_q_11_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__17478\,
            in1 => \N__15524\,
            in2 => \N__15881\,
            in3 => \N__16292\,
            lcout => \M_current_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17349\,
            ce => 'H',
            sr => \N__15465\
        );

    \M_current_address_q_3_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__16293\,
            in1 => \N__15518\,
            in2 => \N__15140\,
            in3 => \N__17479\,
            lcout => \M_current_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17349\,
            ce => 'H',
            sr => \N__15465\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_6_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__15288\,
            in1 => \N__17613\,
            in2 => \N__15869\,
            in3 => \N__16285\,
            lcout => \this_start_data_delay.this_edge_detector.N_216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_3_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__15159\,
            in1 => \N__17614\,
            in2 => \N__20372\,
            in3 => \N__16284\,
            lcout => \this_start_data_delay.this_edge_detector.N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_8_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__16286\,
            in1 => \N__16045\,
            in2 => \N__16835\,
            in3 => \N__17612\,
            lcout => \this_start_data_delay.this_edge_detector.N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_10_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__15913\,
            in1 => \N__17619\,
            in2 => \N__20368\,
            in3 => \N__16287\,
            lcout => \this_start_data_delay.this_edge_detector.N_220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_11_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16288\,
            in1 => \N__16406\,
            in2 => \N__17626\,
            in3 => \N__19203\,
            lcout => \this_start_data_delay.this_edge_detector.N_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_13_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16289\,
            in1 => \N__15868\,
            in2 => \N__17627\,
            in3 => \N__19081\,
            lcout => \this_start_data_delay.this_edge_detector.N_223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_17_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15827\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_this_vram_write_en_0_sqmuxa_0_a3_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17569\,
            in1 => \N__17453\,
            in2 => \_gnd_net_\,
            in3 => \N__16332\,
            lcout => \M_this_vram_write_en_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_16_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15833\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_7_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__16280\,
            in1 => \N__17624\,
            in2 => \N__15721\,
            in3 => \N__17140\,
            lcout => \this_start_data_delay.this_edge_detector.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_0_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__17623\,
            in1 => \N__15582\,
            in2 => \N__17141\,
            in3 => \N__16279\,
            lcout => \this_start_data_delay.this_edge_detector.N_210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_18_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16688\,
            lcout => \this_start_address_delay.this_delay.M_pipe_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.this_delay.M_pipe_q_19_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16679\,
            lcout => \M_this_start_address_delay_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_ns_1_0__m7_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19661\,
            in1 => \N__16841\,
            in2 => \_gnd_net_\,
            in3 => \N__16673\,
            lcout => \M_state_q_ns_1_0__N_24_mux\,
            ltout => \M_state_q_ns_1_0__N_24_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_ns_1_0__m9_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__16169\,
            in1 => \_gnd_net_\,
            in2 => \N__16667\,
            in3 => \N__17451\,
            lcout => OPEN,
            ltout => \M_state_q_ns_1_0__N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_0_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__17740\,
            in1 => \N__17615\,
            in2 => \N__16664\,
            in3 => \N__16290\,
            lcout => \M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17361\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_1_LC_21_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__16566\,
            in1 => \N__17606\,
            in2 => \N__16834\,
            in3 => \N__16281\,
            lcout => \this_start_data_delay.this_edge_detector.N_211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_current_address_q_3_0_4_LC_21_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__16282\,
            in1 => \N__16432\,
            in2 => \N__16405\,
            in3 => \N__17625\,
            lcout => \this_start_data_delay.this_edge_detector.N_214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_ns_1_0__m14_LC_21_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__16283\,
            in1 => \N__16190\,
            in2 => \N__16178\,
            in3 => \N__16165\,
            lcout => OPEN,
            ltout => \M_state_q_ns_1_0__i12_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_1_LC_21_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__17744\,
            in1 => \N__17607\,
            in2 => \N__17507\,
            in3 => \N__17452\,
            lcout => \M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_this_vram_write_data_0_LC_21_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17136\,
            in2 => \_gnd_net_\,
            in3 => \N__20285\,
            lcout => \M_this_vram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_wclke_3_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19318\,
            in1 => \N__19243\,
            in2 => \N__19155\,
            in3 => \N__20327\,
            lcout => \this_vram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI1GH72_12_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17993\,
            in1 => \N__19610\,
            in2 => \_gnd_net_\,
            in3 => \N__17894\,
            lcout => \this_vram.mem_N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5OL72_12_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19621\,
            in1 => \N__19412\,
            in2 => \_gnd_net_\,
            in3 => \N__18122\,
            lcout => \this_vram.mem_N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI4K10H_9_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17924\,
            in1 => \N__20006\,
            in2 => \_gnd_net_\,
            in3 => \N__17777\,
            lcout => \N_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_ns_1_0__m7_5_LC_22_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16922\,
            in1 => \N__16910\,
            in2 => \N__16893\,
            in3 => \N__16853\,
            lcout => \M_state_q_ns_1_0__m7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_this_vram_write_data_1_LC_22_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__16830\,
            in1 => \N__20284\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_0_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19470\,
            in1 => \N__16703\,
            in2 => \_gnd_net_\,
            in3 => \N__18008\,
            lcout => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_wclke_3_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19324\,
            in1 => \N__19239\,
            in2 => \N__19156\,
            in3 => \N__20329\,
            lcout => \this_vram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_wclke_3_LC_23_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20330\,
            in1 => \N__19149\,
            in2 => \N__19244\,
            in3 => \N__19325\,
            lcout => \this_vram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_11_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18806\,
            in1 => \N__17855\,
            in2 => \_gnd_net_\,
            in3 => \N__17848\,
            lcout => \M_this_vram_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_0_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17918\,
            in1 => \N__17909\,
            in2 => \_gnd_net_\,
            in3 => \N__19513\,
            lcout => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI25P11_0_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19514\,
            in1 => \N__17888\,
            in2 => \_gnd_net_\,
            in3 => \N__17870\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OL72_12_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18875\,
            in2 => \N__17858\,
            in3 => \N__19619\,
            lcout => \this_vram.mem_N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18914\,
            in1 => \N__19562\,
            in2 => \_gnd_net_\,
            in3 => \N__17849\,
            lcout => \M_this_vram_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_wclke_3_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__19308\,
            in1 => \N__19237\,
            in2 => \N__19142\,
            in3 => \N__20326\,
            lcout => \this_vram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19529\,
            in1 => \N__18845\,
            in2 => \_gnd_net_\,
            in3 => \N__19622\,
            lcout => \this_vram.mem_N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI9M0SU_9_LC_23_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20021\,
            in2 => \_gnd_net_\,
            in3 => \N__18362\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNIUSK11_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18176\,
            in1 => \N__18164\,
            in2 => \_gnd_net_\,
            in3 => \N__19473\,
            lcout => \this_vram.mem_mem_1_1_RNIUSKZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18149\,
            in1 => \N__19472\,
            in2 => \_gnd_net_\,
            in3 => \N__18134\,
            lcout => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18110\,
            in1 => \N__18095\,
            in2 => \_gnd_net_\,
            in3 => \N__19474\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_0_RNIU0NZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__18035\,
            in1 => \_gnd_net_\,
            in2 => \N__18083\,
            in3 => \N__19634\,
            lcout => \this_vram.mem_N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18059\,
            in1 => \N__18050\,
            in2 => \_gnd_net_\,
            in3 => \N__19471\,
            lcout => \this_vram.mem_mem_0_0_RNIQOIZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI25P11_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18029\,
            in1 => \N__19516\,
            in2 => \_gnd_net_\,
            in3 => \N__18023\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19633\,
            in1 => \_gnd_net_\,
            in2 => \N__18923\,
            in3 => \N__18920\,
            lcout => \this_vram.mem_N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18902\,
            in1 => \N__18890\,
            in2 => \_gnd_net_\,
            in3 => \N__19515\,
            lcout => \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18869\,
            in1 => \N__19519\,
            in2 => \_gnd_net_\,
            in3 => \N__18860\,
            lcout => \this_vram.mem_mem_3_0_RNI05PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18839\,
            in1 => \N__18824\,
            in2 => \_gnd_net_\,
            in3 => \N__19518\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_1_RNI01N11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5GH72_12_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19620\,
            in1 => \_gnd_net_\,
            in2 => \N__18809\,
            in3 => \N__18776\,
            lcout => \this_vram.mem_N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNISOI11_0_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18800\,
            in1 => \N__19517\,
            in2 => \_gnd_net_\,
            in3 => \N__18785\,
            lcout => \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNI01N11_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19522\,
            in1 => \N__18770\,
            in2 => \_gnd_net_\,
            in3 => \N__18755\,
            lcout => \this_vram.mem_mem_2_1_RNI01NZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNISOI11_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18740\,
            in1 => \N__19520\,
            in2 => \_gnd_net_\,
            in3 => \N__18725\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_0_1_RNISOIZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__19643\,
            in1 => \_gnd_net_\,
            in2 => \N__19637\,
            in3 => \N__19632\,
            lcout => \this_vram.mem_N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_RNISSK11_LC_24_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19556\,
            in1 => \N__19521\,
            in2 => \_gnd_net_\,
            in3 => \N__19541\,
            lcout => \this_vram.mem_mem_1_0_RNISSKZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19523\,
            in1 => \N__19439\,
            in2 => \_gnd_net_\,
            in3 => \N__19424\,
            lcout => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_wclke_3_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19307\,
            in1 => \N__19238\,
            in2 => \N__19157\,
            in3 => \N__20320\,
            lcout => \this_vram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_0_wclke_3_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19315\,
            in1 => \N__19204\,
            in2 => \N__19151\,
            in3 => \N__20317\,
            lcout => \this_vram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_6_0_wclke_3_LC_24_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19316\,
            in1 => \N__19221\,
            in2 => \N__19150\,
            in3 => \N__20318\,
            lcout => \this_vram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_7_0_wclke_3_LC_24_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19317\,
            in1 => \N__19222\,
            in2 => \N__19112\,
            in3 => \N__20319\,
            lcout => \this_vram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_this_vram_write_data_2_LC_24_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19035\,
            in2 => \_gnd_net_\,
            in3 => \N__20313\,
            lcout => \M_this_vram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.this_edge_detector.M_this_vram_write_data_3_LC_24_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20349\,
            in2 => \_gnd_net_\,
            in3 => \N__20328\,
            lcout => \M_this_vram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI3N285N2_9_LC_24_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__19864\,
            in1 => \N__20150\,
            in2 => \N__20020\,
            in3 => \N__20135\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIGKVAG41_9_LC_26_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20007\,
            in1 => \N__19865\,
            in2 => \_gnd_net_\,
            in3 => \N__19835\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_ns_1_0__m7_4_LC_32_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19715\,
            in1 => \N__19694\,
            in2 => \N__19682\,
            in3 => \N__19673\,
            lcout => \M_state_q_ns_1_0__m7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
