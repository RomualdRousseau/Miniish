-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 30 2022 22:04:54

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__42118\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41398\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40382\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \this_vga_signals.g1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2_mb_rn_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.g2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal \this_vga_signals.g2_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.g3_2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1_3_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_m2_1\ : std_logic;
signal \this_vga_signals.if_N_9_i\ : std_logic;
signal \this_vga_signals.if_m1_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb2_i_0\ : std_logic;
signal \this_vga_signals.g2_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1_3_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1_3_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_2\ : std_logic;
signal \this_vga_signals.g1_1_0\ : std_logic;
signal \this_vga_signals.g1_4_cascade_\ : std_logic;
signal rgb_c_4 : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.vaddress_m2_2\ : std_logic;
signal port_clk_c : std_logic;
signal \this_vga_signals.g2\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.N_935_0\ : std_logic;
signal port_data_rw_0_i : std_logic;
signal \this_vga_signals.g2_2_0\ : std_logic;
signal rgb_c_0 : std_logic;
signal rgb_c_1 : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.SUM_2_i_i_1_0_3_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_2_x1_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x1_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_i_1_1_3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_x0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x0\ : std_logic;
signal \this_vga_signals.SUM_2_i_i_1_0_3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_x1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_x1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_ns\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_ns_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2_mb_sn\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_3\ : std_logic;
signal \this_vga_signals.g1_0_0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_0_1_0\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_4_cascade_\ : std_logic;
signal \this_vga_signals.g2_1_0\ : std_logic;
signal \this_vga_signals.g0_4_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0\ : std_logic;
signal \this_vga_signals.g0_0_6\ : std_logic;
signal \this_vga_signals.g1_0_0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_4\ : std_logic;
signal \this_vga_signals.g3_0\ : std_logic;
signal \this_vga_signals.N_3_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.g2_0_0_0\ : std_logic;
signal \this_vga_signals.g3_x0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.g3_x1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb2_i\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_vga_signals.g3_0_a2_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2\ : std_logic;
signal \this_vga_signals.g0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.if_i4_mux_0\ : std_logic;
signal \this_vga_signals.vaddress_N_3_i_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g2_4_0\ : std_logic;
signal \this_vga_signals.g2_0_0\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_2_2_N_2L1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_2_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.N_1_4_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c2_2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c2_2\ : std_logic;
signal \this_vga_signals.N_4_3\ : std_logic;
signal \this_vga_signals.g1_1_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.g0_0_i_a5_1\ : std_logic;
signal \this_vga_signals.N_8\ : std_logic;
signal \this_vga_signals.N_6_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \this_vga_signals.g3_0_0\ : std_logic;
signal \this_vga_signals.g3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_0_2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i\ : std_logic;
signal \this_vga_signals.g0_15\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb2_0\ : std_logic;
signal rgb_c_3 : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_1_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i\ : std_logic;
signal \this_vga_signals.g3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_c_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_ac0_3_d\ : std_logic;
signal \this_vga_signals.M_vcounter_q_RNI0FQEQVZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_m6_0\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_4\ : std_logic;
signal \this_vga_signals.g0_0\ : std_logic;
signal \this_vga_signals.g0_0_0_0\ : std_logic;
signal \this_vga_signals.g3\ : std_logic;
signal \this_vga_signals.g0_0_0_a2_2_0\ : std_logic;
signal \this_vga_signals.g0_6_0_a2_3\ : std_logic;
signal \this_vga_signals.N_12_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3\ : std_logic;
signal \this_vga_signals.g0_1_1\ : std_logic;
signal rgb_c_2 : std_logic;
signal \this_vga_signals.vsync_1_0_a2_3\ : std_logic;
signal \this_vga_signals.vsync_1_0_a2_4\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_vga_signals.if_N_6_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0_0\ : std_logic;
signal \this_vga_signals.vvisibility_i_o2_1_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_m2_e_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.N_822_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_9_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_0_0\ : std_logic;
signal \this_vga_signals.r_N_4_mux_1_cascade_\ : std_logic;
signal \this_vga_signals.N_24_0_1\ : std_logic;
signal \this_vga_signals.un2_hsynclt6_0_cascade_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\ : std_logic;
signal \this_vga_signals.r_N_4_mux_0\ : std_logic;
signal \this_vga_signals.N_24_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_4_2_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.g0_0_i_a5_1_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.r_N_4_mux_cascade_\ : std_logic;
signal \this_vga_signals.N_24_0\ : std_logic;
signal \this_vga_signals.r_N_4_mux\ : std_logic;
signal \this_vga_signals.N_32_0\ : std_logic;
signal \this_vga_signals.N_24_0_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_0_0\ : std_logic;
signal \this_vga_signals.g0_23_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\ : std_logic;
signal \this_vga_signals.g0_1_0_0\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.g0_0_2_0\ : std_logic;
signal \this_vga_signals.un2_hsynclt7\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal rgb_c_5 : std_logic;
signal \this_vga_signals.if_N_8_i_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_9_0_0_cascade_\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \this_vga_signals.un4_hsynclto3_0_cascade_\ : std_logic;
signal this_vga_signals_un4_lvisibility_1 : std_logic;
signal \this_vga_signals_M_vcounter_q_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.N_935_0_g\ : std_logic;
signal \this_vga_signals.N_1212_g\ : std_logic;
signal \this_vga_signals.un4_hsynclto7_0\ : std_logic;
signal \this_vga_signals.un4_hsynclt9\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals_M_vcounter_q_7\ : std_logic;
signal \this_vga_signals.g0_0_2\ : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.g0_0_3_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9\ : std_logic;
signal \this_vga_signals.N_935_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \this_vga_signals.g0_0_0\ : std_logic;
signal \M_vcounter_q_esr_RNIQJSA2_0_9\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3\ : std_logic;
signal \this_vga_signals.d_N_11_cascade_\ : std_logic;
signal \this_vga_ramdac.m6\ : std_logic;
signal \this_vga_ramdac.N_2687_reto\ : std_logic;
signal \this_vga_ramdac.N_28_i_reto\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \this_vga_ramdac.N_2690_reto\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt4\ : std_logic;
signal \this_vga_ramdac.N_2691_reto\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \this_vga_ramdac.N_2689_reto\ : std_logic;
signal \this_vga_signals.N_822_0\ : std_logic;
signal \this_vga_signals.M_lcounter_q_3_i_o2_2_1_1\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \M_pcounter_q_ret_1_RNI4VLK7_cascade_\ : std_logic;
signal \this_vga_ramdac.N_2686_reto\ : std_logic;
signal \this_vga_ramdac.i2_mux\ : std_logic;
signal \M_pcounter_q_ret_1_RNI4VLK7\ : std_logic;
signal \this_vga_ramdac.N_2688_reto\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.g0_6_0_0\ : std_logic;
signal \M_hcounter_q_esr_RNIU8TO_9\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_0\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_vga_signals.N_2_8_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_2_am\ : std_logic;
signal \this_vga_signals.haddress_1Z0Z_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_0_3\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_2_bm\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.if_N_8_i_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.if_N_9_1\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_1_cascade_\ : std_logic;
signal \this_vga_signals.N_3_0\ : std_logic;
signal \this_vga_signals.SUM_3_i_0_0\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_1_0\ : std_logic;
signal \N_28_0\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt7_0\ : std_logic;
signal \this_vga_signals.M_lcounter_q_3_i_o2_0_1\ : std_logic;
signal \this_vga_signals.pixel_clk_i\ : std_logic;
signal \this_vga_signals.N_83_1_cascade_\ : std_logic;
signal \this_vga_signals.N_2_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_2_1\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_0Z0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.N_809_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \N_34_0\ : std_logic;
signal port_nmib_1_i : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal \M_this_map_ram_write_data_0\ : std_logic;
signal \M_this_map_ram_write_data_3\ : std_logic;
signal \M_this_map_ram_write_data_4\ : std_logic;
signal dma_0_i : std_logic;
signal \this_vga_signals.N_819_0\ : std_logic;
signal \this_vga_signals.N_827_0_cascade_\ : std_logic;
signal \this_vga_signals.N_826_0\ : std_logic;
signal \this_vga_signals.GZ0Z_406\ : std_logic;
signal \this_vga_signals.N_83_1\ : std_logic;
signal \this_pixel_clk_M_counter_q_0\ : std_logic;
signal \M_this_map_ram_write_data_1\ : std_logic;
signal \M_this_map_ram_write_data_2\ : std_logic;
signal \M_this_map_ram_write_data_7\ : std_logic;
signal \M_this_map_ram_write_data_5\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \N_825_0\ : std_logic;
signal \this_vga_signals_M_lcounter_q_0\ : std_logic;
signal \this_ppu.N_759_0\ : std_logic;
signal \this_vga_signals_M_lcounter_q_1\ : std_logic;
signal \this_vga_signals_M_vcounter_q_9\ : std_logic;
signal \this_ppu.N_5_4_cascade_\ : std_logic;
signal \this_ppu.oam_cache.mem_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\ : std_logic;
signal \M_this_map_ram_read_data_0\ : std_logic;
signal \M_this_ppu_spr_addr_6\ : std_logic;
signal \this_spr_ram.mem_out_bus4_2\ : std_logic;
signal \this_spr_ram.mem_out_bus0_2\ : std_logic;
signal \M_state_q_RNIQER3C_9\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \this_ppu.N_806\ : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \this_spr_ram.mem_out_bus4_0\ : std_logic;
signal \this_spr_ram.mem_out_bus0_0\ : std_logic;
signal \M_this_map_ram_read_data_2\ : std_logic;
signal \M_this_ppu_spr_addr_8\ : std_logic;
signal \M_this_map_ram_read_data_1\ : std_logic;
signal \M_this_ppu_spr_addr_7\ : std_logic;
signal \M_this_map_ram_read_data_3\ : std_logic;
signal \M_this_ppu_spr_addr_9\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \M_this_ppu_spr_addr_10\ : std_logic;
signal \this_ppu.oam_cache.mem_3\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_3\ : std_logic;
signal \this_ppu.oam_cache.mem_2\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_2\ : std_logic;
signal \M_this_map_ram_write_data_6\ : std_logic;
signal \this_spr_ram.mem_mem_0_1_RNIM6VFZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_2\ : std_logic;
signal \this_spr_ram.mem_out_bus3_2\ : std_logic;
signal \this_spr_ram.mem_mem_3_1_RNISI5GZ0_cascade_\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2\ : std_logic;
signal \M_this_spr_ram_read_data_2\ : std_logic;
signal \M_this_spr_ram_read_data_2_cascade_\ : std_logic;
signal \this_spr_ram.mem_out_bus6_2\ : std_logic;
signal \this_spr_ram.mem_out_bus2_2\ : std_logic;
signal \this_spr_ram.mem_mem_2_1_RNIQE3GZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_0\ : std_logic;
signal \this_spr_ram.mem_out_bus3_0\ : std_logic;
signal \this_spr_ram.mem_mem_3_0_RNIQI5GZ0_cascade_\ : std_logic;
signal \M_this_spr_ram_read_data_0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_1\ : std_logic;
signal \this_spr_ram.mem_out_bus3_1\ : std_logic;
signal \this_spr_ram.mem_out_bus6_0\ : std_logic;
signal \this_spr_ram.mem_out_bus2_0\ : std_logic;
signal \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\ : std_logic;
signal \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\ : std_logic;
signal \M_this_spr_ram_read_data_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c3_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c6_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c2\ : std_logic;
signal \this_ppu.M_state_qZ0Z_8\ : std_logic;
signal \this_spr_ram.mem_out_bus6_3\ : std_logic;
signal \this_spr_ram.mem_out_bus2_3\ : std_logic;
signal \this_spr_ram.mem_out_bus6_1\ : std_logic;
signal \this_spr_ram.mem_out_bus2_1\ : std_logic;
signal \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0_cascade_\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1\ : std_logic;
signal \this_spr_ram.mem_WE_6\ : std_logic;
signal \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\ : std_logic;
signal \M_this_spr_ram_read_data_3\ : std_logic;
signal \this_spr_ram.mem_out_bus4_1\ : std_logic;
signal \this_spr_ram.mem_out_bus0_1\ : std_logic;
signal \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_c6\ : std_logic;
signal \this_ppu.N_754_0\ : std_logic;
signal \this_ppu.M_last_q_RNIGL6V4\ : std_logic;
signal \this_spr_ram.mem_WE_8\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_11\ : std_logic;
signal \M_this_state_d_0_sqmuxa\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_11_cascade_\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_11\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_6_s1\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_7\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_2\ : std_logic;
signal \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_4_cascade_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_4\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_6\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_3\ : std_logic;
signal \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\ : std_logic;
signal \this_spr_ram.mem_out_bus4_3\ : std_logic;
signal \this_spr_ram.mem_out_bus0_3\ : std_logic;
signal \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_8\ : std_logic;
signal \this_spr_ram.mem_out_bus7_3\ : std_logic;
signal \this_spr_ram.mem_out_bus3_3\ : std_logic;
signal \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_5\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_3\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_4\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_spr_ram.mem_WE_10\ : std_logic;
signal \M_this_spr_ram_write_data_2\ : std_logic;
signal \this_ppu.oam_cache.mem_5\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_5\ : std_logic;
signal \M_this_spr_ram_write_data_1\ : std_logic;
signal \N_609\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_q_cry_1_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \M_this_data_count_q_cry_8_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_q_s_10\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_q_cry_10_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_q_cry_11_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_11\ : std_logic;
signal \this_ppu.N_91\ : std_logic;
signal \this_ppu.N_760_0_cascade_\ : std_logic;
signal \this_ppu.N_762_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_5\ : std_logic;
signal \this_ppu.M_last_q\ : std_logic;
signal \this_ppu.N_5_4\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_268_i_0_0_cascade_\ : std_logic;
signal \this_ppu.M_count_qZ0Z_5\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_1323_0_cascade_\ : std_logic;
signal \this_ppu.M_count_qZ0Z_1\ : std_logic;
signal \this_ppu.M_count_qZ0Z_7\ : std_logic;
signal \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_3\ : std_logic;
signal \M_this_oam_address_qZ0Z_6\ : std_logic;
signal \M_this_oam_address_qZ0Z_7\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_6\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_7\ : std_logic;
signal port_enb_c : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \N_309_0_cascade_\ : std_logic;
signal \M_this_data_count_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_q_cry_5_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_data_count_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_q_s_13\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_q_s_8\ : std_logic;
signal \N_660_i\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \N_257\ : std_logic;
signal \this_ppu.M_state_qZ0Z_7\ : std_logic;
signal \M_this_oam_address_qZ0Z_1\ : std_logic;
signal \M_this_oam_address_qZ0Z_0\ : std_logic;
signal \N_314_1\ : std_logic;
signal \this_ppu.N_268_i_0_0\ : std_logic;
signal \this_ppu.N_1323_0\ : std_logic;
signal \this_ppu.M_count_qZ0Z_0\ : std_logic;
signal \N_611\ : std_logic;
signal \M_this_ppu_oam_addr_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_13\ : std_logic;
signal \M_this_oam_ram_write_data_13\ : std_logic;
signal \M_this_oam_address_qZ0Z_2\ : std_logic;
signal \M_this_oam_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_oam_address_q_c2\ : std_logic;
signal \un1_M_this_oam_address_q_c4\ : std_logic;
signal \M_this_oam_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_oam_address_q_c4_cascade_\ : std_logic;
signal \M_this_oam_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_oam_address_q_c6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_18\ : std_logic;
signal \M_this_oam_ram_write_data_18\ : std_logic;
signal \M_this_data_tmp_qZ0Z_21\ : std_logic;
signal \M_this_oam_ram_write_data_21\ : std_logic;
signal \M_this_spr_address_qZ0Z_0\ : std_logic;
signal \bfn_19_13_0_\ : std_logic;
signal \M_this_spr_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_spr_address_q_cry_0\ : std_logic;
signal \M_this_spr_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_spr_address_q_cry_1\ : std_logic;
signal \M_this_spr_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_spr_address_q_cry_2\ : std_logic;
signal \M_this_spr_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_spr_address_q_cry_3\ : std_logic;
signal \M_this_spr_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_spr_address_q_cry_4\ : std_logic;
signal \M_this_spr_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_spr_address_q_cry_5\ : std_logic;
signal \M_this_spr_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_spr_address_q_cry_6\ : std_logic;
signal \un1_M_this_spr_address_q_cry_7\ : std_logic;
signal \M_this_spr_address_qZ0Z_8\ : std_logic;
signal \bfn_19_14_0_\ : std_logic;
signal \M_this_spr_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_spr_address_q_cry_8\ : std_logic;
signal \M_this_spr_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_spr_address_q_cry_9\ : std_logic;
signal \un1_M_this_spr_address_q_cry_10\ : std_logic;
signal \un1_M_this_spr_address_q_cry_11\ : std_logic;
signal \un1_M_this_spr_address_q_cry_12\ : std_logic;
signal \N_1310_0\ : std_logic;
signal \bfn_19_17_0_\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \M_this_scroll_qZ0Z_9\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_0\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \M_this_scroll_qZ0Z_10\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_1\ : std_logic;
signal \M_this_ppu_vram_addr_3\ : std_logic;
signal \M_this_scroll_qZ0Z_11\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_2\ : std_logic;
signal \M_this_ppu_vram_addr_4\ : std_logic;
signal \M_this_scroll_qZ0Z_12\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_3\ : std_logic;
signal \M_this_scroll_qZ0Z_13\ : std_logic;
signal \M_this_ppu_vram_addr_5\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_4\ : std_logic;
signal \M_this_scroll_qZ0Z_14\ : std_logic;
signal \M_this_ppu_vram_addr_6\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_5\ : std_logic;
signal \this_ppu.M_haddress_qZ0Z_7\ : std_logic;
signal \M_this_scroll_qZ0Z_15\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_6\ : std_logic;
signal \this_ppu.un1_M_hoffset_d_cry_7\ : std_logic;
signal \bfn_19_18_0_\ : std_logic;
signal \this_ppu.oam_cache.mem_1\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_1\ : std_logic;
signal \this_ppu.N_61_i_cascade_\ : std_logic;
signal \this_ppu.N_769_0\ : std_logic;
signal \this_ppu.M_state_q_srsts_i_i_o2_4_2\ : std_logic;
signal \this_ppu.M_state_qZ0Z_6\ : std_logic;
signal \this_ppu.un1_M_state_q_2_0_cascade_\ : std_logic;
signal \M_this_ppu_oam_addr_5\ : std_logic;
signal \this_ppu.M_oamcurr_qc_0_1\ : std_logic;
signal \this_ppu.un1_M_oamcurr_q_2_c5\ : std_logic;
signal \this_ppu.M_oamcurr_qZ0Z_6\ : std_logic;
signal \N_504_g\ : std_logic;
signal \this_ppu.N_17_0\ : std_logic;
signal \this_ppu.N_329_0_cascade_\ : std_logic;
signal \this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2\ : std_logic;
signal \this_ppu.N_21_0\ : std_logic;
signal \this_ppu.un1_M_oamcurr_q_2_c3\ : std_logic;
signal \this_ppu.N_23_0\ : std_logic;
signal \this_ppu.N_329_0\ : std_logic;
signal \M_this_ppu_oam_addr_0\ : std_logic;
signal \M_this_ppu_oam_addr_1\ : std_logic;
signal \this_ppu.un1_M_state_q_2_0\ : std_logic;
signal \this_ppu.N_19_0\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c2_cascade_\ : std_logic;
signal \M_this_data_tmp_qZ0Z_8\ : std_logic;
signal \M_this_oam_ram_write_data_8\ : std_logic;
signal \M_this_data_tmp_qZ0Z_9\ : std_logic;
signal \M_this_oam_ram_write_data_9\ : std_logic;
signal \N_1294_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_14\ : std_logic;
signal \M_this_oam_ram_write_data_14\ : std_logic;
signal \this_ppu.oam_cache.mem_6\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_6\ : std_logic;
signal \this_ppu.un20_i_a4_0_a3_0_a2_1Z0Z_3_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal \N_260\ : std_logic;
signal \this_ppu.N_406\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_12\ : std_logic;
signal dma_axb3 : std_logic;
signal \this_ppu_un20_i_a4_0_a3_0_a2_3_0_cascade_\ : std_logic;
signal dma_0 : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_10\ : std_logic;
signal \this_ppu.N_414_1_cascade_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \this_ppu.N_267\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_scroll_qZ0Z_8\ : std_logic;
signal \bfn_20_19_0_\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_1\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_2\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_3\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_4\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_5\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_6\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_7\ : std_logic;
signal \bfn_20_20_0_\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_8\ : std_logic;
signal \this_ppu.N_242_0\ : std_logic;
signal \this_ppu.oam_cache.mem_4\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_4\ : std_logic;
signal \this_ppu.M_hoffset_d_0_sqmuxa_7\ : std_logic;
signal \this_ppu.M_state_qZ0Z_9\ : std_logic;
signal \this_ppu.N_772_0\ : std_logic;
signal \this_ppu.N_760_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \this_ppu.N_799_cascade_\ : std_logic;
signal \this_ppu.N_779_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_4\ : std_logic;
signal \this_ppu.M_state_qZ0Z_2\ : std_logic;
signal \this_ppu.N_255\ : std_logic;
signal \this_ppu.N_756_0\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_c5\ : std_logic;
signal \this_ppu.M_last_q_RNIITCPC\ : std_logic;
signal \bfn_20_24_0_\ : std_logic;
signal \this_ppu.M_oamidx_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_oamidx_q_cry_0_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_oamidx_q_cry_0\ : std_logic;
signal \this_ppu.un1_M_oamidx_q_cry_1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_oamidx_q_cry_1\ : std_logic;
signal \this_ppu.un1_M_oamidx_q_cry_2\ : std_logic;
signal \this_ppu.M_oamidx_qZ1Z_2\ : std_logic;
signal \M_this_ppu_oam_addr_3\ : std_logic;
signal \this_ppu.M_oamidx_qZ0Z_3\ : std_logic;
signal \M_this_ppu_oam_addr_2\ : std_logic;
signal \this_ppu.M_state_q_srsts_0_a3_0_o2_0_6\ : std_logic;
signal \this_ppu.N_228_0_i_1_0\ : std_logic;
signal \this_ppu.M_oamidx_qZ0Z_0\ : std_logic;
signal \N_332_0\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_7_cascade_\ : std_logic;
signal \this_ppu.N_405\ : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_13_cascade_\ : std_logic;
signal \this_ppu.N_324_0\ : std_logic;
signal \this_ppu.N_424_cascade_\ : std_logic;
signal \this_ppu.N_449\ : std_logic;
signal \M_this_state_q_RNI1G0LZ0Z_1\ : std_logic;
signal \this_ppu.N_341_0\ : std_logic;
signal \this_ppu.N_934\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal this_ppu_un20_i_a4_0_a2_0_a2_0_2 : std_logic;
signal \N_311_0_cascade_\ : std_logic;
signal \M_this_state_q_RNI244K2Z0Z_10\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \M_this_state_q_RNIR71EZ0Z_10\ : std_logic;
signal \this_ppu.hspr_cry_0_c_inv_RNI1203\ : std_logic;
signal \bfn_21_17_0_\ : std_logic;
signal \M_this_ppu_spr_addr_1\ : std_logic;
signal \this_ppu.hspr_cry_0\ : std_logic;
signal \this_ppu.hspr_cry_1\ : std_logic;
signal \M_this_ppu_spr_addr_2\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_9\ : std_logic;
signal \bfn_21_18_0_\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_0\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_1\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_2\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_3\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_4\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_5\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_6\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_7\ : std_logic;
signal \this_ppu.M_hoffset_q_i_8\ : std_logic;
signal \bfn_21_19_0_\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_2_cry_8\ : std_logic;
signal \this_ppu.vspr12_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNOZ0\ : std_logic;
signal \bfn_21_20_0_\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_1\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_2\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_3\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_4\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_5\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_6\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_7\ : std_logic;
signal \bfn_21_21_0_\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_8\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_8_THRU_CO\ : std_logic;
signal \this_ppu.vspr_cry_0_c_inv_RNIFK43\ : std_logic;
signal \bfn_21_22_0_\ : std_logic;
signal \M_this_ppu_spr_addr_4\ : std_logic;
signal \this_ppu.vspr_cry_0\ : std_logic;
signal \this_ppu.vspr_cry_1\ : std_logic;
signal \M_this_ppu_spr_addr_5\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_17\ : std_logic;
signal \this_ppu.oam_cache.mem_17\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_17\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \bfn_21_23_0_\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_0\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_1\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_3\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_2\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_4\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_3\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_5\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_4\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_6\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_5\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_7\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_6\ : std_logic;
signal \this_ppu.un1_M_voffset_d_cry_7\ : std_logic;
signal \bfn_21_24_0_\ : std_logic;
signal \this_ppu.N_756_0_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_2\ : std_logic;
signal \M_this_oam_ram_write_data_2\ : std_logic;
signal \M_this_data_tmp_qZ0Z_16\ : std_logic;
signal \M_this_oam_ram_write_data_16\ : std_logic;
signal \M_this_data_tmp_qZ0Z_5\ : std_logic;
signal \M_this_oam_ram_write_data_5\ : std_logic;
signal \M_this_data_tmp_qZ0Z_15\ : std_logic;
signal \M_this_oam_ram_write_data_15\ : std_logic;
signal \M_this_data_tmp_qZ0Z_19\ : std_logic;
signal \M_this_oam_ram_write_data_19\ : std_logic;
signal \N_1286_0\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \this_ppu.N_511\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_0_i_1Z0Z_6_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal this_ppu_un20_i_a4_0_a3_0_a2_1_1 : std_logic;
signal port_rw_in : std_logic;
signal \this_ppu.N_321_0\ : std_logic;
signal \this_ppu.N_328_0\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0_cascade_\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_i_1_0Z0Z_0\ : std_logic;
signal \this_ppu.N_416\ : std_logic;
signal \this_ppu.M_hoffset_q_i_0\ : std_logic;
signal \bfn_22_18_0_\ : std_logic;
signal \this_ppu.M_hoffset_q_i_1\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_0\ : std_logic;
signal \this_ppu.M_hoffset_q_i_2\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_1\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_0\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_2\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_1\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_3\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_2\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_4\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_3\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_4\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_cry_7\ : std_logic;
signal \bfn_22_19_0_\ : std_logic;
signal \this_ppu.vspr16_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_ac0_13_i\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNOZ0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNOZ0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNOZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_6\ : std_logic;
signal \this_ppu.un1_oam_data_1_8\ : std_logic;
signal \this_ppu.un1_oam_data_1_7\ : std_logic;
signal \this_ppu.un1_oam_data_1_5\ : std_logic;
signal \bfn_22_21_0_\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_1\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_2\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNOZ0\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_3\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_3\ : std_logic;
signal \this_ppu.read_data_RNI3DGK1_14\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_5\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_6\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_7\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNOZ0\ : std_logic;
signal \this_ppu.M_hoffset_qZ0Z_8\ : std_logic;
signal \bfn_22_22_0_\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_8\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_CO\ : std_logic;
signal \this_ppu.oam_cache.mem_18\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_18\ : std_logic;
signal \M_this_scroll_qZ0Z_0\ : std_logic;
signal \M_this_scroll_qZ0Z_1\ : std_logic;
signal \M_this_scroll_qZ0Z_5\ : std_logic;
signal \M_this_scroll_qZ0Z_3\ : std_logic;
signal \M_this_scroll_qZ0Z_4\ : std_logic;
signal \M_this_scroll_qZ0Z_6\ : std_logic;
signal \M_this_scroll_qZ0Z_7\ : std_logic;
signal \this_ppu.M_voffset_q_i_0\ : std_logic;
signal \bfn_22_24_0_\ : std_logic;
signal \this_ppu.M_voffset_qZ0Z_1\ : std_logic;
signal \this_ppu.M_voffset_q_i_1\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_0\ : std_logic;
signal \this_ppu.M_voffset_qZ0Z_2\ : std_logic;
signal \this_ppu.M_voffset_q_i_2\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_1\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_5\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_2\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_6\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_3\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_7\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_8\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_8\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_5\ : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_9\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_7\ : std_logic;
signal \this_ppu.M_voffset_qZ0Z_8\ : std_logic;
signal \this_ppu.M_voffset_q_i_8\ : std_logic;
signal \bfn_22_25_0_\ : std_logic;
signal \this_ppu.un1_M_voffset_q_cry_8\ : std_logic;
signal \this_ppu.M_state_d14_1\ : std_logic;
signal \N_433\ : std_logic;
signal \N_438\ : std_logic;
signal \M_this_data_tmp_qZ0Z_12\ : std_logic;
signal \M_this_oam_ram_write_data_12\ : std_logic;
signal \M_this_scroll_qZ0Z_2\ : std_logic;
signal \N_1318_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_0\ : std_logic;
signal \M_this_oam_ram_write_data_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_1\ : std_logic;
signal \M_this_oam_ram_write_data_1\ : std_logic;
signal \N_434\ : std_logic;
signal \this_spr_ram.mem_out_bus5_3\ : std_logic;
signal \this_spr_ram.mem_out_bus1_3\ : std_logic;
signal \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_WE_0\ : std_logic;
signal \this_ppu.oam_cache.mem_7\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_7\ : std_logic;
signal \this_ppu.hspr\ : std_logic;
signal \M_this_ppu_spr_addr_0\ : std_logic;
signal \M_this_spr_ram_write_data_0\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_2\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_3\ : std_logic;
signal \this_ppu.N_510\ : std_logic;
signal port_address_in_1 : std_logic;
signal \this_ppu.N_916\ : std_logic;
signal \this_ppu.M_state_q_inv_1\ : std_logic;
signal \this_ppu.vspr\ : std_logic;
signal \M_this_ppu_spr_addr_3\ : std_logic;
signal \this_ppu.oam_cache.mem_15\ : std_logic;
signal \this_ppu.oam_cache.mem_14\ : std_logic;
signal \M_this_oam_ram_read_data_22\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_21\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_21\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_9\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_c7\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_10\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_c7_cascade_\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNOZ0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNOZ0\ : std_logic;
signal \this_ppu.oam_cache.mem_12\ : std_logic;
signal \this_ppu.M_hoffset_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNOZ0\ : std_logic;
signal \this_ppu.oam_cache.mem_9\ : std_logic;
signal \this_ppu.oam_cache.mem_8\ : std_logic;
signal \this_ppu.oam_cache.mem_13\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_c4\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_8\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_c4_cascade_\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_7\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNOZ0\ : std_logic;
signal \this_ppu.read_data_RNI80ET_11\ : std_logic;
signal \M_this_oam_ram_read_data_11\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_11\ : std_logic;
signal \this_ppu.oam_cache.mem_11\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_6\ : std_logic;
signal \this_ppu.M_hoffset_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_4\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNOZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_4_c5_0\ : std_logic;
signal \M_this_oam_ram_read_data_23\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_23\ : std_logic;
signal port_data_c_0 : std_logic;
signal port_data_c_1 : std_logic;
signal \this_ppu.oam_cache.mem_16\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_16\ : std_logic;
signal \M_this_data_tmp_qZ0Z_20\ : std_logic;
signal \M_this_oam_ram_write_data_20\ : std_logic;
signal \M_this_oam_ram_write_data_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_7\ : std_logic;
signal \M_this_oam_ram_write_data_3\ : std_logic;
signal \M_this_data_tmp_qZ0Z_3\ : std_logic;
signal \M_this_oam_ram_write_data_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_4\ : std_logic;
signal \N_1302_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_23\ : std_logic;
signal \M_this_oam_ram_write_data_23\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_17\ : std_logic;
signal \N_440\ : std_logic;
signal \N_437\ : std_logic;
signal \M_this_data_tmp_qZ0Z_22\ : std_logic;
signal \M_this_oam_ram_write_data_22\ : std_logic;
signal port_data_c_6 : std_logic;
signal \N_439\ : std_logic;
signal \this_spr_ram.mem_WE_2\ : std_logic;
signal \this_spr_ram.mem_WE_4\ : std_logic;
signal \this_spr_ram.mem_out_bus5_1\ : std_logic;
signal \this_spr_ram.mem_out_bus1_1\ : std_logic;
signal \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_WE_14\ : std_logic;
signal \N_260_0\ : std_logic;
signal \M_this_spr_address_qZ0Z_13\ : std_logic;
signal \M_this_spr_address_qZ0Z_12\ : std_logic;
signal \M_this_spr_address_qZ0Z_11\ : std_logic;
signal \this_spr_ram.mem_WE_12\ : std_logic;
signal \this_ppu.N_545\ : std_logic;
signal \M_this_spr_ram_write_data_3\ : std_logic;
signal port_address_in_4 : std_logic;
signal port_address_in_0 : std_logic;
signal \this_ppu.N_610\ : std_logic;
signal \M_this_state_d_0_sqmuxa_2\ : std_logic;
signal led_c_1 : std_logic;
signal \N_608\ : std_logic;
signal \M_this_substate_qZ0\ : std_logic;
signal \M_this_state_qZ0Z_13\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \this_ppu.oam_cache.mem_10\ : std_logic;
signal \this_ppu.un1_M_hoffset_q_5\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_18\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal port_data_c_7 : std_logic;
signal \M_this_ctrl_flags_qZ0Z_7\ : std_logic;
signal \N_312_0\ : std_logic;
signal \M_this_ext_address_qZ0Z_0\ : std_logic;
signal \bfn_24_21_0_\ : std_logic;
signal \M_this_ext_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_ext_address_q_cry_0_THRU_CO\ : std_logic;
signal \un1_M_this_ext_address_q_cry_0\ : std_logic;
signal \M_this_ext_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_ext_address_q_cry_1_THRU_CO\ : std_logic;
signal \un1_M_this_ext_address_q_cry_1\ : std_logic;
signal \M_this_ext_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_ext_address_q_cry_2_THRU_CO\ : std_logic;
signal \un1_M_this_ext_address_q_cry_2\ : std_logic;
signal \un1_M_this_ext_address_q_cry_3\ : std_logic;
signal \un1_M_this_ext_address_q_cry_4\ : std_logic;
signal \un1_M_this_ext_address_q_cry_5\ : std_logic;
signal \un1_M_this_ext_address_q_cry_6\ : std_logic;
signal \un1_M_this_ext_address_q_cry_7\ : std_logic;
signal \M_this_ext_address_qZ0Z_8\ : std_logic;
signal \un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0\ : std_logic;
signal \bfn_24_22_0_\ : std_logic;
signal \M_this_ext_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_8\ : std_logic;
signal \un1_M_this_ext_address_q_cry_9\ : std_logic;
signal \un1_M_this_ext_address_q_cry_10\ : std_logic;
signal \un1_M_this_ext_address_q_cry_11\ : std_logic;
signal \un1_M_this_ext_address_q_cry_12\ : std_logic;
signal \M_this_ext_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_13\ : std_logic;
signal \M_this_ext_address_qZ0Z_15\ : std_logic;
signal \un1_M_this_ext_address_q_cry_14\ : std_logic;
signal \un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0\ : std_logic;
signal \M_this_oam_ram_read_data_13\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_13\ : std_logic;
signal \M_this_oam_ram_read_data_15\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_15\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_3\ : std_logic;
signal \M_this_oam_ram_read_data_8\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_8\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_16\ : std_logic;
signal \M_this_oam_ram_read_data_10\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_10\ : std_logic;
signal \M_this_oam_ram_read_data_25\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_25\ : std_logic;
signal \M_this_oam_ram_read_data_26\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_26\ : std_logic;
signal \M_this_data_tmp_qZ0Z_10\ : std_logic;
signal \M_this_oam_ram_write_data_10\ : std_logic;
signal \M_this_data_tmp_qZ0Z_6\ : std_logic;
signal \M_this_oam_ram_write_data_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_11\ : std_logic;
signal \M_this_oam_ram_write_data_11\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_2\ : std_logic;
signal \this_ppu.un12lto7Z0Z_4\ : std_logic;
signal \M_this_oam_ram_read_data_4\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_4\ : std_logic;
signal \M_this_oam_ram_read_data_5\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_5\ : std_logic;
signal \M_this_oam_ram_read_data_6\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_6\ : std_logic;
signal \M_this_oam_ram_read_data_7\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_7\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_1\ : std_logic;
signal \M_this_oam_ram_read_data_2\ : std_logic;
signal \M_this_oam_ram_read_data_1\ : std_logic;
signal \M_this_oam_ram_read_data_3\ : std_logic;
signal \M_this_oam_ram_read_data_0\ : std_logic;
signal \this_ppu.un12lto7Z0Z_5\ : std_logic;
signal \M_this_oam_ram_read_data_27\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_27\ : std_logic;
signal \this_ppu.un1_oam_data_1_3\ : std_logic;
signal \M_this_oam_ram_read_data_29\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_29\ : std_logic;
signal \this_ppu.un1_oam_data_1_4\ : std_logic;
signal \M_this_oam_ram_read_data_31\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_31\ : std_logic;
signal \M_this_oam_ram_read_data_19\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_19\ : std_logic;
signal \M_this_oam_ram_read_data_20\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_20\ : std_logic;
signal \M_this_oam_ram_read_data_24\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_24\ : std_logic;
signal \M_this_oam_ram_read_data_18\ : std_logic;
signal \this_ppu.un1_oam_data_1_2\ : std_logic;
signal \M_this_data_tmp_qZ0Z_17\ : std_logic;
signal \M_this_oam_ram_write_data_17\ : std_logic;
signal \this_ppu.un1_oam_data_1_4_c2\ : std_logic;
signal \M_this_oam_ram_read_data_30\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_30\ : std_logic;
signal \M_this_oam_ram_read_data_9\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_9\ : std_logic;
signal \N_435\ : std_logic;
signal \M_this_oam_ram_read_data_17\ : std_logic;
signal \M_this_oam_ram_read_data_16\ : std_logic;
signal \this_ppu.un1_oam_data_1_1\ : std_logic;
signal \this_spr_ram.mem_out_bus5_2\ : std_logic;
signal \this_spr_ram.mem_out_bus1_2\ : std_logic;
signal \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\ : std_logic;
signal \this_spr_ram.mem_out_bus5_0\ : std_logic;
signal \this_spr_ram.mem_out_bus1_0\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\ : std_logic;
signal \un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0\ : std_logic;
signal port_data_c_2 : std_logic;
signal \M_this_ext_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_ext_address_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_ext_address_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_ext_address_q_cry_5_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_ext_address_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_ext_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0\ : std_logic;
signal \M_this_ext_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0\ : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_ext_address_qZ0Z_12\ : std_logic;
signal \N_309_0\ : std_logic;
signal \N_311_0\ : std_logic;
signal port_data_c_5 : std_logic;
signal \un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0\ : std_logic;
signal \M_this_ext_address_qZ0Z_13\ : std_logic;
signal clk_0_c_g : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;
signal \M_this_oam_ram_read_data_12\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_12\ : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_oam_ram_write_data_0_sqmuxa\ : std_logic;
signal \N_436\ : std_logic;
signal \M_this_oam_ram_read_data_28\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_28\ : std_logic;
signal \M_this_oam_ram_read_data_14\ : std_logic;
signal \this_ppu.M_state_qZ0Z_3\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_14\ : std_logic;
signal port_address_in_2 : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_6 : std_logic;
signal port_address_in_5 : std_logic;
signal \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1Z0Z_0\ : std_logic;
signal port_address_in_7 : std_logic;
signal \this_ppu.N_173\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_map_ram_read_data_3\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_2\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_1\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_0\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__33298\&\N__33349\&\N__33397\&\N__33448\&\N__33502\&\N__34306\&\N__32923\&\N__35206\&\N__33004\&\N__33073\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__19234\&\N__19267\&\N__19297\&\N__19324\&\N__19351\&\N__19381\&\N__19408\&\N__18685\&\N__18715\&\N__18742\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__19645\&'0'&'0'&'0'&\N__19768\&'0'&'0'&'0'&\N__19780\&'0'&'0'&'0'&\N__19657\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__33292\&\N__33342\&\N__33391\&\N__33442\&\N__33496\&\N__34297\&\N__32916\&\N__35200\&\N__32998\&\N__33067\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__19228\&\N__19261\&\N__19291\&\N__19318\&\N__19345\&\N__19375\&\N__19402\&\N__18679\&\N__18709\&\N__18736\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__19759\&'0'&'0'&'0'&\N__21706\&'0'&'0'&'0'&\N__19747\&'0'&'0'&'0'&\N__19636\&'0';
    \M_this_oam_ram_read_data_15\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_14\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_13\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_12\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_11\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_10\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_9\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_8\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_7\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_6\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_5\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_4\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_3\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_2\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_1\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_0\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__28480\&\N__25384\&\N__30196\&\N__30091\&\N__28687\&\N__28753\;
    \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24298\&\N__24334\&\N__25195\&\N__25150\&\N__25270\&\N__25312\;
    \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ <= \N__31939\&\N__28996\&\N__25327\&\N__33664\&\N__38065\&\N__38101\&\N__29074\&\N__28570\&\N__36085\&\N__38089\&\N__31960\&\N__36049\&\N__36067\&\N__32005\&\N__33592\&\N__33610\;
    \M_this_oam_ram_read_data_31\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_30\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_29\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_28\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_27\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_26\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_25\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_24\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_23\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_22\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_21\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_20\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_19\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_18\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_17\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_16\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__28474\&\N__25378\&\N__30190\&\N__30085\&\N__28681\&\N__28747\;
    \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24292\&\N__24328\&\N__25189\&\N__25144\&\N__25264\&\N__25306\;
    \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ <= \N__36349\&\N__36184\&\N__33688\&\N__36340\&\N__39163\&\N__39109\&\N__33580\&\N__33700\&\N__35965\&\N__36322\&\N__26974\&\N__35365\&\N__31924\&\N__26995\&\N__38365\&\N__31978\;
    \this_ppu.oam_cache.mem_15\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(15);
    \this_ppu.oam_cache.mem_14\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(14);
    \this_ppu.oam_cache.mem_13\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(13);
    \this_ppu.oam_cache.mem_12\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(12);
    \this_ppu.oam_cache.mem_11\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_ppu.oam_cache.mem_10\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(10);
    \this_ppu.oam_cache.mem_9\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(9);
    \this_ppu.oam_cache.mem_8\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(8);
    \this_ppu.oam_cache.mem_7\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(7);
    \this_ppu.oam_cache.mem_6\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(6);
    \this_ppu.oam_cache.mem_5\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(5);
    \this_ppu.oam_cache.mem_4\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(4);
    \this_ppu.oam_cache.mem_3\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_ppu.oam_cache.mem_2\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(2);
    \this_ppu.oam_cache.mem_1\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_ppu.oam_cache.mem_0\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28783\&\N__28828\&\N__28597\&\N__28861\;
    \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__30127\&\N__30229\&\N__30307\&\N__29896\;
    \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\ <= \N__37909\&\N__41356\&\N__37927\&\N__39529\&\N__34990\&\N__37858\&\N__39121\&\N__37882\&\N__38290\&\N__38311\&\N__38332\&\N__38026\&\N__37900\&\N__38056\&\N__38272\&\N__38281\;
    \this_ppu.oam_cache.mem_18\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(2);
    \this_ppu.oam_cache.mem_17\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_ppu.oam_cache.mem_16\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28777\&\N__28822\&\N__28591\&\N__28855\;
    \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__30121\&\N__30223\&\N__30301\&\N__29889\;
    \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\ <= \N__38575\&\N__39148\&\N__38161\&\N__41629\&\N__38194\&\N__38119\&\N__38137\&\N__38455\&\N__35635\&\N__34516\&\N__34444\&\N__38473\&\N__38521\&\N__36535\&\N__35953\&\N__37873\;
    \this_spr_ram.mem_out_bus0_1\ <= \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus0_0\ <= \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__20779\&\N__21008\&\N__21424\&\N__21175\&\N__20350\&\N__31165\&\N__31388\&\N__34727\&\N__30802\&\N__30995\&\N__33994\;
    \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__27235\&\N__27409\&\N__27642\&\N__27892\&\N__25618\&\N__25864\&\N__26040\&\N__26297\&\N__26467\&\N__26745\&\N__26945\;
    \this_spr_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22945\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33863\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus0_3\ <= \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus0_2\ <= \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__20838\&\N__21009\&\N__21423\&\N__21176\&\N__20351\&\N__31190\&\N__31417\&\N__34796\&\N__30750\&\N__30949\&\N__33993\;
    \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__27213\&\N__27377\&\N__27615\&\N__27887\&\N__25604\&\N__25793\&\N__26039\&\N__26278\&\N__26466\&\N__26731\&\N__26944\;
    \this_spr_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37111\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22733\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus1_1\ <= \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus1_0\ <= \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__20780\&\N__21010\&\N__21425\&\N__21201\&\N__20363\&\N__31219\&\N__31447\&\N__34797\&\N__30787\&\N__30983\&\N__33988\;
    \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__27186\&\N__27376\&\N__27614\&\N__27875\&\N__25584\&\N__25836\&\N__26000\&\N__26231\&\N__26465\&\N__26725\&\N__26911\;
    \this_spr_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22926\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33844\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus1_3\ <= \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus1_2\ <= \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__20815\&\N__21011\&\N__21426\&\N__21202\&\N__20274\&\N__31245\&\N__31473\&\N__34760\&\N__30815\&\N__31010\&\N__33989\;
    \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__27176\&\N__27307\&\N__27539\&\N__27855\&\N__25555\&\N__25840\&\N__25999\&\N__26239\&\N__26482\&\N__26726\&\N__26893\;
    \this_spr_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37099\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22707\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus2_1\ <= \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus2_0\ <= \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__20837\&\N__20992\&\N__21409\&\N__21128\&\N__20262\&\N__31231\&\N__31459\&\N__34785\&\N__30866\&\N__31022\&\N__34011\;
    \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__27221\&\N__27420\&\N__27650\&\N__27879\&\N__25638\&\N__25873\&\N__26050\&\N__26308\&\N__26521\&\N__26748\&\N__26954\;
    \this_spr_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22953\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33876\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus2_3\ <= \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus2_2\ <= \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__20836\&\N__21018\&\N__21410\&\N__21164\&\N__20234\&\N__31232\&\N__31460\&\N__34809\&\N__30880\&\N__31047\&\N__34072\;
    \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__27223\&\N__27393\&\N__27629\&\N__27847\&\N__25630\&\N__25869\&\N__26049\&\N__26300\&\N__26522\&\N__26740\&\N__26955\;
    \this_spr_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37154\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22729\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus3_1\ <= \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus3_0\ <= \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__20835\&\N__21019\&\N__21439\&\N__21171\&\N__20302\&\N__31257\&\N__31485\&\N__34810\&\N__30881\&\N__31069\&\N__34087\;
    \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__27222\&\N__27421\&\N__27651\&\N__27851\&\N__25619\&\N__25868\&\N__26051\&\N__26261\&\N__26513\&\N__26736\&\N__26946\;
    \this_spr_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22964\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33894\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus3_3\ <= \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus3_2\ <= \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__20805\&\N__21029\&\N__21440\&\N__21200\&\N__20335\&\N__31258\&\N__31486\&\N__34799\&\N__30888\&\N__31086\&\N__34088\;
    \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__27236\&\N__27438\&\N__27612\&\N__27852\&\N__25641\&\N__25857\&\N__26052\&\N__26312\&\N__26514\&\N__26671\&\N__26947\;
    \this_spr_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37161\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22744\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus4_1\ <= \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus4_0\ <= \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__20834\&\N__21030\&\N__21452\&\N__21196\&\N__20355\&\N__31277\&\N__31503\&\N__34800\&\N__30889\&\N__31087\&\N__34095\;
    \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__27243\&\N__27449\&\N__27662\&\N__27853\&\N__25639\&\N__25853\&\N__26061\&\N__26316\&\N__26523\&\N__26735\&\N__26958\;
    \this_spr_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22969\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33898\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus4_3\ <= \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus4_2\ <= \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__20833\&\N__21034\&\N__21453\&\N__21220\&\N__20364\&\N__31278\&\N__31504\&\N__34798\&\N__30839\&\N__31009\&\N__34096\;
    \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__27247\&\N__27454\&\N__27667\&\N__27854\&\N__25645\&\N__25792\&\N__26062\&\N__26317\&\N__26524\&\N__26747\&\N__26959\;
    \this_spr_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37165\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22735\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus5_1\ <= \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus5_0\ <= \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__20841\&\N__21012\&\N__21427\&\N__21221\&\N__20312\&\N__31265\&\N__31400\&\N__34795\&\N__30816\&\N__31035\&\N__34012\;
    \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__27194\&\N__27381\&\N__27619\&\N__27868\&\N__25577\&\N__25841\&\N__26007\&\N__26218\&\N__26456\&\N__26730\&\N__26897\;
    \this_spr_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22946\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33864\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus5_3\ <= \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus5_2\ <= \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__20842\&\N__21013\&\N__21428\&\N__21222\&\N__20342\&\N__31279\&\N__31493\&\N__34794\&\N__30840\&\N__31057\&\N__34037\;
    \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__27214\&\N__27410\&\N__27611\&\N__27880\&\N__25597\&\N__25842\&\N__26008\&\N__26274\&\N__26508\&\N__26672\&\N__26898\;
    \this_spr_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37125\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22743\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus6_1\ <= \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus6_0\ <= \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__20839\&\N__21014\&\N__21429\&\N__21235\&\N__20346\&\N__31291\&\N__31429\&\N__34808\&\N__30810\&\N__31076\&\N__34064\;
    \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__27209\&\N__27431\&\N__27643\&\N__27888\&\N__25614\&\N__25865\&\N__26041\&\N__26307\&\N__26489\&\N__26746\&\N__26936\;
    \this_spr_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22960\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33877\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus6_3\ <= \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus6_2\ <= \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__20840\&\N__21015\&\N__21447\&\N__21236\&\N__20362\&\N__31301\&\N__31505\&\N__34792\&\N__30811\&\N__31088\&\N__34065\;
    \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__27234\&\N__27445\&\N__27658\&\N__27893\&\N__25626\&\N__25866\&\N__26042\&\N__26299\&\N__26463\&\N__26749\&\N__26937\;
    \this_spr_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37140\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22734\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus7_1\ <= \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus7_0\ <= \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__20831\&\N__21016\&\N__21448\&\N__21243\&\N__20365\&\N__31308\&\N__31512\&\N__34793\&\N__30862\&\N__31095\&\N__34085\;
    \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__27193\&\N__27453\&\N__27666\&\N__27897\&\N__25637\&\N__25843\&\N__26059\&\N__26235\&\N__26512\&\N__26741\&\N__26956\;
    \this_spr_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22968\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__33887\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus7_3\ <= \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus7_2\ <= \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__20832\&\N__21017\&\N__21454\&\N__21244\&\N__20325\&\N__31309\&\N__31513\&\N__34807\&\N__30879\&\N__31096\&\N__34086\;
    \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__27233\&\N__27408\&\N__27613\&\N__27898\&\N__25640\&\N__25867\&\N__26060\&\N__26298\&\N__26464\&\N__26721\&\N__26957\;
    \this_spr_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__37153\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22742\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__14839\&\N__18778\&\N__18013\&\N__17188\&\N__17197\&\N__17215\&\N__17164\&\N__17206\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__31863\&\N__28087\&\N__28138\&\N__28213\&\N__28303\&\N__28381\&\N__27961\&\N__29356\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21544\&\N__19735\&\N__20092\&\N__21514\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40442\,
            RE => \N__23663\,
            WCLKE => \N__22177\,
            WCLK => \N__40443\,
            WE => \N__23667\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40452\,
            RE => \N__23712\,
            WCLKE => \N__22159\,
            WCLK => \N__40453\,
            WE => \N__23713\
        );

    \this_oam_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40462\,
            RE => \N__23753\,
            WCLKE => \N__39384\,
            WCLK => \N__40463\,
            WE => \N__23662\
        );

    \this_oam_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40464\,
            RE => \N__23595\,
            WCLKE => \N__39385\,
            WCLK => \N__40465\,
            WE => \N__23521\
        );

    \this_ppu.oam_cache.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40447\,
            RE => \N__23719\,
            WCLKE => \N__41601\,
            WCLK => \N__40448\,
            WE => \N__23751\
        );

    \this_ppu.oam_cache.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40457\,
            RE => \N__23752\,
            WCLKE => \N__41552\,
            WCLK => \N__40458\,
            WE => \N__23514\
        );

    \this_spr_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40434\,
            RE => \N__23718\,
            WCLKE => \N__36115\,
            WCLK => \N__40435\,
            WE => \N__23513\
        );

    \this_spr_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40417\,
            RE => \N__23676\,
            WCLKE => \N__36114\,
            WCLK => \N__40418\,
            WE => \N__23717\
        );

    \this_spr_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40396\,
            RE => \N__23675\,
            WCLKE => \N__37216\,
            WCLK => \N__40397\,
            WE => \N__23430\
        );

    \this_spr_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40376\,
            RE => \N__23614\,
            WCLKE => \N__37212\,
            WCLK => \N__40377\,
            WE => \N__23674\
        );

    \this_spr_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40388\,
            RE => \N__23596\,
            WCLKE => \N__22768\,
            WCLK => \N__40389\,
            WE => \N__23597\
        );

    \this_spr_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40369\,
            RE => \N__23525\,
            WCLKE => \N__22764\,
            WCLK => \N__40370\,
            WE => \N__23523\
        );

    \this_spr_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40342\,
            RE => \N__23524\,
            WCLKE => \N__22368\,
            WCLK => \N__40343\,
            WE => \N__23522\
        );

    \this_spr_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40325\,
            RE => \N__23456\,
            WCLKE => \N__22372\,
            WCLK => \N__40324\,
            WE => \N__23447\
        );

    \this_spr_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40310\,
            RE => \N__23455\,
            WCLKE => \N__22020\,
            WCLK => \N__40311\,
            WE => \N__23446\
        );

    \this_spr_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40302\,
            RE => \N__23445\,
            WCLKE => \N__22024\,
            WCLK => \N__40303\,
            WE => \N__23363\
        );

    \this_spr_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40351\,
            RE => \N__23613\,
            WCLKE => \N__36156\,
            WCLK => \N__40352\,
            WE => \N__23429\
        );

    \this_spr_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40332\,
            RE => \N__23548\,
            WCLKE => \N__36157\,
            WCLK => \N__40331\,
            WE => \N__23546\
        );

    \this_spr_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40319\,
            RE => \N__23547\,
            WCLKE => \N__36168\,
            WCLK => \N__40320\,
            WE => \N__23428\
        );

    \this_spr_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40306\,
            RE => \N__23476\,
            WCLKE => \N__36172\,
            WCLK => \N__40307\,
            WE => \N__23481\
        );

    \this_spr_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40298\,
            RE => \N__23477\,
            WCLKE => \N__34213\,
            WCLK => \N__40299\,
            WE => \N__23405\
        );

    \this_spr_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40288\,
            RE => \N__23545\,
            WCLKE => \N__34212\,
            WCLK => \N__40289\,
            WE => \N__23591\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__40293\,
            RE => \N__23475\,
            WCLKE => \N__20107\,
            WCLK => \N__40294\,
            WE => \N__23454\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__42116\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42118\,
            DIN => \N__42117\,
            DOUT => \N__42116\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__42118\,
            PADOUT => \N__42117\,
            PADIN => \N__42116\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42107\,
            DIN => \N__42106\,
            DOUT => \N__42105\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42107\,
            PADOUT => \N__42106\,
            PADIN => \N__42105\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42098\,
            DIN => \N__42097\,
            DOUT => \N__42096\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42098\,
            PADOUT => \N__42097\,
            PADIN => \N__42096\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42089\,
            DIN => \N__42088\,
            DOUT => \N__42087\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42089\,
            PADOUT => \N__42088\,
            PADIN => \N__42087\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17236\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42080\,
            DIN => \N__42079\,
            DOUT => \N__42078\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42080\,
            PADOUT => \N__42079\,
            PADIN => \N__42078\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15973\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42071\,
            DIN => \N__42070\,
            DOUT => \N__42069\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42071\,
            PADOUT => \N__42070\,
            PADIN => \N__42069\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__23636\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42062\,
            DIN => \N__42061\,
            DOUT => \N__42060\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42062\,
            PADOUT => \N__42061\,
            PADIN => \N__42060\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36904\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42053\,
            DIN => \N__42052\,
            DOUT => \N__42051\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42053\,
            PADOUT => \N__42052\,
            PADIN => \N__42051\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42044\,
            DIN => \N__42043\,
            DOUT => \N__42042\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42044\,
            PADOUT => \N__42043\,
            PADIN => \N__42042\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42035\,
            DIN => \N__42034\,
            DOUT => \N__42033\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42035\,
            PADOUT => \N__42034\,
            PADIN => \N__42033\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42026\,
            DIN => \N__42025\,
            DOUT => \N__42024\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42026\,
            PADOUT => \N__42025\,
            PADIN => \N__42024\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42017\,
            DIN => \N__42016\,
            DOUT => \N__42015\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42017\,
            PADOUT => \N__42016\,
            PADIN => \N__42015\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__42008\,
            DIN => \N__42007\,
            DOUT => \N__42006\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__42008\,
            PADOUT => \N__42007\,
            PADIN => \N__42006\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41999\,
            DIN => \N__41998\,
            DOUT => \N__41997\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41999\,
            PADOUT => \N__41998\,
            PADIN => \N__41997\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__37717\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19593\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41990\,
            DIN => \N__41989\,
            DOUT => \N__41988\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41990\,
            PADOUT => \N__41989\,
            PADIN => \N__41988\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__37681\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19620\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41981\,
            DIN => \N__41980\,
            DOUT => \N__41979\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41981\,
            PADOUT => \N__41980\,
            PADIN => \N__41979\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__37636\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19609\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41972\,
            DIN => \N__41971\,
            DOUT => \N__41970\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41972\,
            PADOUT => \N__41971\,
            PADIN => \N__41970\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__37600\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19607\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41963\,
            DIN => \N__41962\,
            DOUT => \N__41961\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41963\,
            PADOUT => \N__41962\,
            PADIN => \N__41961\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__38626\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19588\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41954\,
            DIN => \N__41953\,
            DOUT => \N__41952\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41954\,
            PADOUT => \N__41953\,
            PADIN => \N__41952\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__41233\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19536\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41945\,
            DIN => \N__41944\,
            DOUT => \N__41943\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41945\,
            PADOUT => \N__41944\,
            PADIN => \N__41943\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__41191\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19587\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41936\,
            DIN => \N__41935\,
            DOUT => \N__41934\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41936\,
            PADOUT => \N__41935\,
            PADIN => \N__41934\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__41146\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19585\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41927\,
            DIN => \N__41926\,
            DOUT => \N__41925\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41927\,
            PADOUT => \N__41926\,
            PADIN => \N__41925\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__38665\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19608\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41918\,
            DIN => \N__41917\,
            DOUT => \N__41916\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41918\,
            PADOUT => \N__41917\,
            PADIN => \N__41916\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__41092\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19624\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41909\,
            DIN => \N__41908\,
            DOUT => \N__41907\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41909\,
            PADOUT => \N__41908\,
            PADIN => \N__41907\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40936\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19589\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41900\,
            DIN => \N__41899\,
            DOUT => \N__41898\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41900\,
            PADOUT => \N__41899\,
            PADIN => \N__41898\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__40492\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19564\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41891\,
            DIN => \N__41890\,
            DOUT => \N__41889\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41891\,
            PADOUT => \N__41890\,
            PADIN => \N__41889\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__38011\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19586\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41882\,
            DIN => \N__41881\,
            DOUT => \N__41880\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41882\,
            PADOUT => \N__41881\,
            PADIN => \N__41880\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37975\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19554\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41873\,
            DIN => \N__41872\,
            DOUT => \N__41871\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41873\,
            PADOUT => \N__41872\,
            PADIN => \N__41871\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37837\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19521\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41864\,
            DIN => \N__41863\,
            DOUT => \N__41862\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41864\,
            PADOUT => \N__41863\,
            PADIN => \N__41862\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37801\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19619\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41855\,
            DIN => \N__41854\,
            DOUT => \N__41853\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41855\,
            PADOUT => \N__41854\,
            PADIN => \N__41853\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41846\,
            DIN => \N__41845\,
            DOUT => \N__41844\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41846\,
            PADOUT => \N__41845\,
            PADIN => \N__41844\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41837\,
            DIN => \N__41836\,
            DOUT => \N__41835\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41837\,
            PADOUT => \N__41836\,
            PADIN => \N__41835\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41828\,
            DIN => \N__41827\,
            DOUT => \N__41826\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41828\,
            PADOUT => \N__41827\,
            PADIN => \N__41826\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41819\,
            DIN => \N__41818\,
            DOUT => \N__41817\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41819\,
            PADOUT => \N__41818\,
            PADIN => \N__41817\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41810\,
            DIN => \N__41809\,
            DOUT => \N__41808\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41810\,
            PADOUT => \N__41809\,
            PADIN => \N__41808\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41801\,
            DIN => \N__41800\,
            DOUT => \N__41799\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41801\,
            PADOUT => \N__41800\,
            PADIN => \N__41799\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41792\,
            DIN => \N__41791\,
            DOUT => \N__41790\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41792\,
            PADOUT => \N__41791\,
            PADIN => \N__41790\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41783\,
            DIN => \N__41782\,
            DOUT => \N__41781\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41783\,
            PADOUT => \N__41782\,
            PADIN => \N__41781\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41774\,
            DIN => \N__41773\,
            DOUT => \N__41772\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41774\,
            PADOUT => \N__41773\,
            PADIN => \N__41772\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13423\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41765\,
            DIN => \N__41764\,
            DOUT => \N__41763\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41765\,
            PADOUT => \N__41764\,
            PADIN => \N__41763\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29239\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41756\,
            DIN => \N__41755\,
            DOUT => \N__41754\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41756\,
            PADOUT => \N__41755\,
            PADIN => \N__41754\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41747\,
            DIN => \N__41746\,
            DOUT => \N__41745\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41747\,
            PADOUT => \N__41746\,
            PADIN => \N__41745\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__18760\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41738\,
            DIN => \N__41737\,
            DOUT => \N__41736\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__41738\,
            PADOUT => \N__41737\,
            PADIN => \N__41736\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__23750\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__19488\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41729\,
            DIN => \N__41728\,
            DOUT => \N__41727\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41729\,
            PADOUT => \N__41728\,
            PADIN => \N__41727\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13399\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41720\,
            DIN => \N__41719\,
            DOUT => \N__41718\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41720\,
            PADOUT => \N__41719\,
            PADIN => \N__41718\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13387\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41711\,
            DIN => \N__41710\,
            DOUT => \N__41709\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41711\,
            PADOUT => \N__41710\,
            PADIN => \N__41709\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15094\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41702\,
            DIN => \N__41701\,
            DOUT => \N__41700\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41702\,
            PADOUT => \N__41701\,
            PADIN => \N__41700\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15031\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41693\,
            DIN => \N__41692\,
            DOUT => \N__41691\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41693\,
            PADOUT => \N__41692\,
            PADIN => \N__41691\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13342\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41684\,
            DIN => \N__41683\,
            DOUT => \N__41682\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41684\,
            PADOUT => \N__41683\,
            PADIN => \N__41682\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15955\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41675\,
            DIN => \N__41674\,
            DOUT => \N__41673\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__41675\,
            PADOUT => \N__41674\,
            PADIN => \N__41673\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41666\,
            DIN => \N__41665\,
            DOUT => \N__41664\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41666\,
            PADOUT => \N__41665\,
            PADIN => \N__41664\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__16441\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__41657\,
            DIN => \N__41656\,
            DOUT => \N__41655\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__41657\,
            PADOUT => \N__41656\,
            PADIN => \N__41655\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__15064\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__10490\ : InMux
    port map (
            O => \N__41638\,
            I => \N__41635\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__41635\,
            I => \N__41632\
        );

    \I__10488\ : Odrv4
    port map (
            O => \N__41632\,
            I => \M_this_oam_ram_read_data_28\
        );

    \I__10487\ : InMux
    port map (
            O => \N__41629\,
            I => \N__41626\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__41626\,
            I => \N__41623\
        );

    \I__10485\ : Span4Mux_h
    port map (
            O => \N__41623\,
            I => \N__41620\
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__41620\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_28\
        );

    \I__10483\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41614\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__41614\,
            I => \N__41611\
        );

    \I__10481\ : Span4Mux_v
    port map (
            O => \N__41611\,
            I => \N__41608\
        );

    \I__10480\ : Odrv4
    port map (
            O => \N__41608\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__10479\ : InMux
    port map (
            O => \N__41605\,
            I => \N__41598\
        );

    \I__10478\ : InMux
    port map (
            O => \N__41604\,
            I => \N__41593\
        );

    \I__10477\ : CascadeMux
    port map (
            O => \N__41603\,
            I => \N__41577\
        );

    \I__10476\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41570\
        );

    \I__10475\ : CEMux
    port map (
            O => \N__41601\,
            I => \N__41561\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__41598\,
            I => \N__41558\
        );

    \I__10473\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41555\
        );

    \I__10472\ : CascadeMux
    port map (
            O => \N__41596\,
            I => \N__41549\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__41593\,
            I => \N__41545\
        );

    \I__10470\ : InMux
    port map (
            O => \N__41592\,
            I => \N__41540\
        );

    \I__10469\ : InMux
    port map (
            O => \N__41591\,
            I => \N__41540\
        );

    \I__10468\ : InMux
    port map (
            O => \N__41590\,
            I => \N__41535\
        );

    \I__10467\ : InMux
    port map (
            O => \N__41589\,
            I => \N__41535\
        );

    \I__10466\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41526\
        );

    \I__10465\ : InMux
    port map (
            O => \N__41587\,
            I => \N__41526\
        );

    \I__10464\ : InMux
    port map (
            O => \N__41586\,
            I => \N__41526\
        );

    \I__10463\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41526\
        );

    \I__10462\ : InMux
    port map (
            O => \N__41584\,
            I => \N__41523\
        );

    \I__10461\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41510\
        );

    \I__10460\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41510\
        );

    \I__10459\ : InMux
    port map (
            O => \N__41581\,
            I => \N__41510\
        );

    \I__10458\ : InMux
    port map (
            O => \N__41580\,
            I => \N__41510\
        );

    \I__10457\ : InMux
    port map (
            O => \N__41577\,
            I => \N__41510\
        );

    \I__10456\ : InMux
    port map (
            O => \N__41576\,
            I => \N__41510\
        );

    \I__10455\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41503\
        );

    \I__10454\ : InMux
    port map (
            O => \N__41574\,
            I => \N__41503\
        );

    \I__10453\ : InMux
    port map (
            O => \N__41573\,
            I => \N__41503\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__41570\,
            I => \N__41500\
        );

    \I__10451\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41495\
        );

    \I__10450\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41495\
        );

    \I__10449\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41486\
        );

    \I__10448\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41486\
        );

    \I__10447\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41486\
        );

    \I__10446\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41486\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__41561\,
            I => \N__41483\
        );

    \I__10444\ : Span4Mux_v
    port map (
            O => \N__41558\,
            I => \N__41478\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__41555\,
            I => \N__41478\
        );

    \I__10442\ : InMux
    port map (
            O => \N__41554\,
            I => \N__41473\
        );

    \I__10441\ : InMux
    port map (
            O => \N__41553\,
            I => \N__41473\
        );

    \I__10440\ : CEMux
    port map (
            O => \N__41552\,
            I => \N__41470\
        );

    \I__10439\ : InMux
    port map (
            O => \N__41549\,
            I => \N__41465\
        );

    \I__10438\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41462\
        );

    \I__10437\ : Span4Mux_h
    port map (
            O => \N__41545\,
            I => \N__41459\
        );

    \I__10436\ : LocalMux
    port map (
            O => \N__41540\,
            I => \N__41448\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__41535\,
            I => \N__41448\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__41526\,
            I => \N__41448\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__41523\,
            I => \N__41448\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__41510\,
            I => \N__41448\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__41503\,
            I => \N__41439\
        );

    \I__10430\ : Span4Mux_v
    port map (
            O => \N__41500\,
            I => \N__41439\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__41495\,
            I => \N__41439\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__41486\,
            I => \N__41439\
        );

    \I__10427\ : Span4Mux_h
    port map (
            O => \N__41483\,
            I => \N__41433\
        );

    \I__10426\ : Span4Mux_v
    port map (
            O => \N__41478\,
            I => \N__41430\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__41473\,
            I => \N__41427\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__41470\,
            I => \N__41424\
        );

    \I__10423\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41419\
        );

    \I__10422\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41419\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__41465\,
            I => \N__41414\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__41462\,
            I => \N__41414\
        );

    \I__10419\ : Span4Mux_h
    port map (
            O => \N__41459\,
            I => \N__41407\
        );

    \I__10418\ : Span4Mux_v
    port map (
            O => \N__41448\,
            I => \N__41407\
        );

    \I__10417\ : Span4Mux_v
    port map (
            O => \N__41439\,
            I => \N__41407\
        );

    \I__10416\ : InMux
    port map (
            O => \N__41438\,
            I => \N__41402\
        );

    \I__10415\ : InMux
    port map (
            O => \N__41437\,
            I => \N__41402\
        );

    \I__10414\ : InMux
    port map (
            O => \N__41436\,
            I => \N__41399\
        );

    \I__10413\ : Span4Mux_h
    port map (
            O => \N__41433\,
            I => \N__41395\
        );

    \I__10412\ : Span4Mux_h
    port map (
            O => \N__41430\,
            I => \N__41390\
        );

    \I__10411\ : Span4Mux_v
    port map (
            O => \N__41427\,
            I => \N__41390\
        );

    \I__10410\ : Span12Mux_s11_v
    port map (
            O => \N__41424\,
            I => \N__41385\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__41419\,
            I => \N__41385\
        );

    \I__10408\ : Span4Mux_v
    port map (
            O => \N__41414\,
            I => \N__41382\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__41407\,
            I => \N__41377\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__41402\,
            I => \N__41377\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__41399\,
            I => \N__41374\
        );

    \I__10404\ : InMux
    port map (
            O => \N__41398\,
            I => \N__41371\
        );

    \I__10403\ : Odrv4
    port map (
            O => \N__41395\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__10402\ : Odrv4
    port map (
            O => \N__41390\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__10401\ : Odrv12
    port map (
            O => \N__41385\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__10400\ : Odrv4
    port map (
            O => \N__41382\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__10399\ : Odrv4
    port map (
            O => \N__41377\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__41374\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__41371\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__10396\ : InMux
    port map (
            O => \N__41356\,
            I => \N__41353\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__41353\,
            I => \N__41350\
        );

    \I__10394\ : Span4Mux_h
    port map (
            O => \N__41350\,
            I => \N__41347\
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__41347\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_14\
        );

    \I__10392\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41341\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41338\
        );

    \I__10390\ : Span4Mux_v
    port map (
            O => \N__41338\,
            I => \N__41335\
        );

    \I__10389\ : Sp12to4
    port map (
            O => \N__41335\,
            I => \N__41332\
        );

    \I__10388\ : Span12Mux_s10_h
    port map (
            O => \N__41332\,
            I => \N__41329\
        );

    \I__10387\ : Odrv12
    port map (
            O => \N__41329\,
            I => port_address_in_2
        );

    \I__10386\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41323\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__41323\,
            I => \N__41320\
        );

    \I__10384\ : Odrv4
    port map (
            O => \N__41320\,
            I => port_address_in_3
        );

    \I__10383\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41314\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__41314\,
            I => port_address_in_6
        );

    \I__10381\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41308\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__41308\,
            I => \N__41305\
        );

    \I__10379\ : Span12Mux_v
    port map (
            O => \N__41305\,
            I => \N__41302\
        );

    \I__10378\ : Odrv12
    port map (
            O => \N__41302\,
            I => port_address_in_5
        );

    \I__10377\ : CascadeMux
    port map (
            O => \N__41299\,
            I => \N__41296\
        );

    \I__10376\ : InMux
    port map (
            O => \N__41296\,
            I => \N__41293\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__41293\,
            I => \N__41290\
        );

    \I__10374\ : Span12Mux_s1_h
    port map (
            O => \N__41290\,
            I => \N__41287\
        );

    \I__10373\ : Odrv12
    port map (
            O => \N__41287\,
            I => \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1Z0Z_0\
        );

    \I__10372\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41281\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__41281\,
            I => \N__41278\
        );

    \I__10370\ : Span12Mux_s2_h
    port map (
            O => \N__41278\,
            I => \N__41275\
        );

    \I__10369\ : Span12Mux_v
    port map (
            O => \N__41275\,
            I => \N__41272\
        );

    \I__10368\ : Odrv12
    port map (
            O => \N__41272\,
            I => port_address_in_7
        );

    \I__10367\ : InMux
    port map (
            O => \N__41269\,
            I => \N__41266\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__41266\,
            I => \N__41263\
        );

    \I__10365\ : Span4Mux_v
    port map (
            O => \N__41263\,
            I => \N__41260\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__41260\,
            I => \N__41256\
        );

    \I__10363\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41253\
        );

    \I__10362\ : Sp12to4
    port map (
            O => \N__41256\,
            I => \N__41248\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41248\
        );

    \I__10360\ : Odrv12
    port map (
            O => \N__41248\,
            I => \this_ppu.N_173\
        );

    \I__10359\ : InMux
    port map (
            O => \N__41245\,
            I => \N__41242\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__41242\,
            I => \N__41239\
        );

    \I__10357\ : Span4Mux_v
    port map (
            O => \N__41239\,
            I => \N__41236\
        );

    \I__10356\ : Odrv4
    port map (
            O => \N__41236\,
            I => \un1_M_this_ext_address_q_cry_4_THRU_CO\
        );

    \I__10355\ : IoInMux
    port map (
            O => \N__41233\,
            I => \N__41230\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__41230\,
            I => \N__41226\
        );

    \I__10353\ : InMux
    port map (
            O => \N__41229\,
            I => \N__41223\
        );

    \I__10352\ : Span4Mux_s2_h
    port map (
            O => \N__41226\,
            I => \N__41219\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41216\
        );

    \I__10350\ : InMux
    port map (
            O => \N__41222\,
            I => \N__41213\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__41219\,
            I => \N__41208\
        );

    \I__10348\ : Span4Mux_h
    port map (
            O => \N__41216\,
            I => \N__41208\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__41213\,
            I => \M_this_ext_address_qZ0Z_5\
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__41208\,
            I => \M_this_ext_address_qZ0Z_5\
        );

    \I__10345\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41200\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__41200\,
            I => \N__41197\
        );

    \I__10343\ : Span4Mux_h
    port map (
            O => \N__41197\,
            I => \N__41194\
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__41194\,
            I => \un1_M_this_ext_address_q_cry_5_THRU_CO\
        );

    \I__10341\ : IoInMux
    port map (
            O => \N__41191\,
            I => \N__41188\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__41188\,
            I => \N__41185\
        );

    \I__10339\ : Span4Mux_s2_h
    port map (
            O => \N__41185\,
            I => \N__41181\
        );

    \I__10338\ : InMux
    port map (
            O => \N__41184\,
            I => \N__41178\
        );

    \I__10337\ : Span4Mux_v
    port map (
            O => \N__41181\,
            I => \N__41174\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__41178\,
            I => \N__41171\
        );

    \I__10335\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41168\
        );

    \I__10334\ : Span4Mux_h
    port map (
            O => \N__41174\,
            I => \N__41163\
        );

    \I__10333\ : Span4Mux_h
    port map (
            O => \N__41171\,
            I => \N__41163\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__41168\,
            I => \M_this_ext_address_qZ0Z_6\
        );

    \I__10331\ : Odrv4
    port map (
            O => \N__41163\,
            I => \M_this_ext_address_qZ0Z_6\
        );

    \I__10330\ : InMux
    port map (
            O => \N__41158\,
            I => \N__41155\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__41155\,
            I => \N__41152\
        );

    \I__10328\ : Span4Mux_h
    port map (
            O => \N__41152\,
            I => \N__41149\
        );

    \I__10327\ : Odrv4
    port map (
            O => \N__41149\,
            I => \un1_M_this_ext_address_q_cry_6_THRU_CO\
        );

    \I__10326\ : IoInMux
    port map (
            O => \N__41146\,
            I => \N__41143\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__41143\,
            I => \N__41140\
        );

    \I__10324\ : IoSpan4Mux
    port map (
            O => \N__41140\,
            I => \N__41137\
        );

    \I__10323\ : Span4Mux_s2_h
    port map (
            O => \N__41137\,
            I => \N__41133\
        );

    \I__10322\ : CascadeMux
    port map (
            O => \N__41136\,
            I => \N__41130\
        );

    \I__10321\ : Span4Mux_h
    port map (
            O => \N__41133\,
            I => \N__41127\
        );

    \I__10320\ : InMux
    port map (
            O => \N__41130\,
            I => \N__41124\
        );

    \I__10319\ : Sp12to4
    port map (
            O => \N__41127\,
            I => \N__41121\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__41124\,
            I => \N__41117\
        );

    \I__10317\ : Span12Mux_v
    port map (
            O => \N__41121\,
            I => \N__41114\
        );

    \I__10316\ : InMux
    port map (
            O => \N__41120\,
            I => \N__41111\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__41117\,
            I => \N__41108\
        );

    \I__10314\ : Odrv12
    port map (
            O => \N__41114\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__41111\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__10312\ : Odrv4
    port map (
            O => \N__41108\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__10311\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41098\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__41098\,
            I => \N__41095\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__41095\,
            I => \un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0\
        );

    \I__10308\ : IoInMux
    port map (
            O => \N__41092\,
            I => \N__41089\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__41089\,
            I => \N__41086\
        );

    \I__10306\ : Span4Mux_s3_v
    port map (
            O => \N__41086\,
            I => \N__41083\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__41083\,
            I => \N__41079\
        );

    \I__10304\ : InMux
    port map (
            O => \N__41082\,
            I => \N__41076\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__41079\,
            I => \N__41073\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__41076\,
            I => \N__41070\
        );

    \I__10301\ : Odrv4
    port map (
            O => \N__41073\,
            I => \M_this_ext_address_qZ0Z_11\
        );

    \I__10300\ : Odrv12
    port map (
            O => \N__41070\,
            I => \M_this_ext_address_qZ0Z_11\
        );

    \I__10299\ : InMux
    port map (
            O => \N__41065\,
            I => \N__41062\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__41062\,
            I => \N__41059\
        );

    \I__10297\ : Odrv4
    port map (
            O => \N__41059\,
            I => \un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0\
        );

    \I__10296\ : CascadeMux
    port map (
            O => \N__41056\,
            I => \N__41051\
        );

    \I__10295\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41048\
        );

    \I__10294\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41045\
        );

    \I__10293\ : InMux
    port map (
            O => \N__41051\,
            I => \N__41042\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__41048\,
            I => \N__41036\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__41045\,
            I => \N__41033\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__41042\,
            I => \N__41030\
        );

    \I__10289\ : InMux
    port map (
            O => \N__41041\,
            I => \N__41026\
        );

    \I__10288\ : CascadeMux
    port map (
            O => \N__41040\,
            I => \N__41023\
        );

    \I__10287\ : InMux
    port map (
            O => \N__41039\,
            I => \N__41020\
        );

    \I__10286\ : Span4Mux_v
    port map (
            O => \N__41036\,
            I => \N__41017\
        );

    \I__10285\ : Span4Mux_v
    port map (
            O => \N__41033\,
            I => \N__41013\
        );

    \I__10284\ : Span4Mux_v
    port map (
            O => \N__41030\,
            I => \N__41010\
        );

    \I__10283\ : InMux
    port map (
            O => \N__41029\,
            I => \N__41007\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__41026\,
            I => \N__41004\
        );

    \I__10281\ : InMux
    port map (
            O => \N__41023\,
            I => \N__41001\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__41020\,
            I => \N__40998\
        );

    \I__10279\ : Span4Mux_v
    port map (
            O => \N__41017\,
            I => \N__40995\
        );

    \I__10278\ : InMux
    port map (
            O => \N__41016\,
            I => \N__40992\
        );

    \I__10277\ : Span4Mux_h
    port map (
            O => \N__41013\,
            I => \N__40989\
        );

    \I__10276\ : Span4Mux_v
    port map (
            O => \N__41010\,
            I => \N__40984\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__41007\,
            I => \N__40984\
        );

    \I__10274\ : Span12Mux_h
    port map (
            O => \N__41004\,
            I => \N__40980\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__41001\,
            I => \N__40977\
        );

    \I__10272\ : Span12Mux_v
    port map (
            O => \N__40998\,
            I => \N__40974\
        );

    \I__10271\ : Span4Mux_h
    port map (
            O => \N__40995\,
            I => \N__40971\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__40992\,
            I => \N__40968\
        );

    \I__10269\ : Span4Mux_h
    port map (
            O => \N__40989\,
            I => \N__40963\
        );

    \I__10268\ : Span4Mux_v
    port map (
            O => \N__40984\,
            I => \N__40963\
        );

    \I__10267\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40960\
        );

    \I__10266\ : Span12Mux_v
    port map (
            O => \N__40980\,
            I => \N__40957\
        );

    \I__10265\ : Span12Mux_v
    port map (
            O => \N__40977\,
            I => \N__40954\
        );

    \I__10264\ : Span12Mux_h
    port map (
            O => \N__40974\,
            I => \N__40943\
        );

    \I__10263\ : Sp12to4
    port map (
            O => \N__40971\,
            I => \N__40943\
        );

    \I__10262\ : Span12Mux_v
    port map (
            O => \N__40968\,
            I => \N__40943\
        );

    \I__10261\ : Sp12to4
    port map (
            O => \N__40963\,
            I => \N__40943\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__40960\,
            I => \N__40943\
        );

    \I__10259\ : Odrv12
    port map (
            O => \N__40957\,
            I => port_data_c_4
        );

    \I__10258\ : Odrv12
    port map (
            O => \N__40954\,
            I => port_data_c_4
        );

    \I__10257\ : Odrv12
    port map (
            O => \N__40943\,
            I => port_data_c_4
        );

    \I__10256\ : IoInMux
    port map (
            O => \N__40936\,
            I => \N__40933\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__40933\,
            I => \N__40930\
        );

    \I__10254\ : Span4Mux_s2_h
    port map (
            O => \N__40930\,
            I => \N__40926\
        );

    \I__10253\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40923\
        );

    \I__10252\ : Span4Mux_h
    port map (
            O => \N__40926\,
            I => \N__40920\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__40923\,
            I => \N__40917\
        );

    \I__10250\ : Odrv4
    port map (
            O => \N__40920\,
            I => \M_this_ext_address_qZ0Z_12\
        );

    \I__10249\ : Odrv12
    port map (
            O => \N__40917\,
            I => \M_this_ext_address_qZ0Z_12\
        );

    \I__10248\ : InMux
    port map (
            O => \N__40912\,
            I => \N__40888\
        );

    \I__10247\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40888\
        );

    \I__10246\ : InMux
    port map (
            O => \N__40910\,
            I => \N__40888\
        );

    \I__10245\ : InMux
    port map (
            O => \N__40909\,
            I => \N__40888\
        );

    \I__10244\ : InMux
    port map (
            O => \N__40908\,
            I => \N__40888\
        );

    \I__10243\ : InMux
    port map (
            O => \N__40907\,
            I => \N__40888\
        );

    \I__10242\ : InMux
    port map (
            O => \N__40906\,
            I => \N__40888\
        );

    \I__10241\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40888\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__40888\,
            I => \N__40876\
        );

    \I__10239\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40869\
        );

    \I__10238\ : InMux
    port map (
            O => \N__40886\,
            I => \N__40869\
        );

    \I__10237\ : InMux
    port map (
            O => \N__40885\,
            I => \N__40869\
        );

    \I__10236\ : InMux
    port map (
            O => \N__40884\,
            I => \N__40856\
        );

    \I__10235\ : InMux
    port map (
            O => \N__40883\,
            I => \N__40856\
        );

    \I__10234\ : InMux
    port map (
            O => \N__40882\,
            I => \N__40856\
        );

    \I__10233\ : InMux
    port map (
            O => \N__40881\,
            I => \N__40856\
        );

    \I__10232\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40856\
        );

    \I__10231\ : InMux
    port map (
            O => \N__40879\,
            I => \N__40856\
        );

    \I__10230\ : Span4Mux_v
    port map (
            O => \N__40876\,
            I => \N__40852\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__40869\,
            I => \N__40849\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__40856\,
            I => \N__40840\
        );

    \I__10227\ : InMux
    port map (
            O => \N__40855\,
            I => \N__40837\
        );

    \I__10226\ : Span4Mux_h
    port map (
            O => \N__40852\,
            I => \N__40831\
        );

    \I__10225\ : Span4Mux_v
    port map (
            O => \N__40849\,
            I => \N__40831\
        );

    \I__10224\ : InMux
    port map (
            O => \N__40848\,
            I => \N__40828\
        );

    \I__10223\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40824\
        );

    \I__10222\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40821\
        );

    \I__10221\ : InMux
    port map (
            O => \N__40845\,
            I => \N__40814\
        );

    \I__10220\ : InMux
    port map (
            O => \N__40844\,
            I => \N__40814\
        );

    \I__10219\ : InMux
    port map (
            O => \N__40843\,
            I => \N__40811\
        );

    \I__10218\ : Span4Mux_v
    port map (
            O => \N__40840\,
            I => \N__40806\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__40837\,
            I => \N__40806\
        );

    \I__10216\ : InMux
    port map (
            O => \N__40836\,
            I => \N__40800\
        );

    \I__10215\ : Span4Mux_v
    port map (
            O => \N__40831\,
            I => \N__40795\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__40828\,
            I => \N__40795\
        );

    \I__10213\ : InMux
    port map (
            O => \N__40827\,
            I => \N__40790\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__40824\,
            I => \N__40785\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__40821\,
            I => \N__40785\
        );

    \I__10210\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40782\
        );

    \I__10209\ : InMux
    port map (
            O => \N__40819\,
            I => \N__40779\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__40814\,
            I => \N__40776\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__40811\,
            I => \N__40771\
        );

    \I__10206\ : Span4Mux_h
    port map (
            O => \N__40806\,
            I => \N__40771\
        );

    \I__10205\ : InMux
    port map (
            O => \N__40805\,
            I => \N__40766\
        );

    \I__10204\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40766\
        );

    \I__10203\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40763\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__40800\,
            I => \N__40760\
        );

    \I__10201\ : Span4Mux_h
    port map (
            O => \N__40795\,
            I => \N__40757\
        );

    \I__10200\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40752\
        );

    \I__10199\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40752\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__40790\,
            I => \N__40739\
        );

    \I__10197\ : Span4Mux_h
    port map (
            O => \N__40785\,
            I => \N__40739\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__40782\,
            I => \N__40739\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__40779\,
            I => \N__40739\
        );

    \I__10194\ : Span4Mux_v
    port map (
            O => \N__40776\,
            I => \N__40739\
        );

    \I__10193\ : Span4Mux_v
    port map (
            O => \N__40771\,
            I => \N__40739\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__40766\,
            I => \N_309_0\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__40763\,
            I => \N_309_0\
        );

    \I__10190\ : Odrv4
    port map (
            O => \N__40760\,
            I => \N_309_0\
        );

    \I__10189\ : Odrv4
    port map (
            O => \N__40757\,
            I => \N_309_0\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__40752\,
            I => \N_309_0\
        );

    \I__10187\ : Odrv4
    port map (
            O => \N__40739\,
            I => \N_309_0\
        );

    \I__10186\ : CascadeMux
    port map (
            O => \N__40726\,
            I => \N__40714\
        );

    \I__10185\ : CascadeMux
    port map (
            O => \N__40725\,
            I => \N__40711\
        );

    \I__10184\ : CascadeMux
    port map (
            O => \N__40724\,
            I => \N__40707\
        );

    \I__10183\ : CascadeMux
    port map (
            O => \N__40723\,
            I => \N__40704\
        );

    \I__10182\ : CascadeMux
    port map (
            O => \N__40722\,
            I => \N__40696\
        );

    \I__10181\ : CascadeMux
    port map (
            O => \N__40721\,
            I => \N__40693\
        );

    \I__10180\ : CascadeMux
    port map (
            O => \N__40720\,
            I => \N__40690\
        );

    \I__10179\ : InMux
    port map (
            O => \N__40719\,
            I => \N__40683\
        );

    \I__10178\ : InMux
    port map (
            O => \N__40718\,
            I => \N__40683\
        );

    \I__10177\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40683\
        );

    \I__10176\ : InMux
    port map (
            O => \N__40714\,
            I => \N__40676\
        );

    \I__10175\ : InMux
    port map (
            O => \N__40711\,
            I => \N__40676\
        );

    \I__10174\ : InMux
    port map (
            O => \N__40710\,
            I => \N__40676\
        );

    \I__10173\ : InMux
    port map (
            O => \N__40707\,
            I => \N__40665\
        );

    \I__10172\ : InMux
    port map (
            O => \N__40704\,
            I => \N__40665\
        );

    \I__10171\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40665\
        );

    \I__10170\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40665\
        );

    \I__10169\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40665\
        );

    \I__10168\ : InMux
    port map (
            O => \N__40700\,
            I => \N__40653\
        );

    \I__10167\ : InMux
    port map (
            O => \N__40699\,
            I => \N__40653\
        );

    \I__10166\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40653\
        );

    \I__10165\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40653\
        );

    \I__10164\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40653\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__40683\,
            I => \N__40650\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__40676\,
            I => \N__40645\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__40665\,
            I => \N__40645\
        );

    \I__10160\ : CascadeMux
    port map (
            O => \N__40664\,
            I => \N__40642\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__40653\,
            I => \N__40639\
        );

    \I__10158\ : Span4Mux_h
    port map (
            O => \N__40650\,
            I => \N__40636\
        );

    \I__10157\ : Span4Mux_v
    port map (
            O => \N__40645\,
            I => \N__40633\
        );

    \I__10156\ : InMux
    port map (
            O => \N__40642\,
            I => \N__40630\
        );

    \I__10155\ : Span4Mux_v
    port map (
            O => \N__40639\,
            I => \N__40627\
        );

    \I__10154\ : Span4Mux_v
    port map (
            O => \N__40636\,
            I => \N__40624\
        );

    \I__10153\ : Span4Mux_h
    port map (
            O => \N__40633\,
            I => \N__40621\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__40630\,
            I => \N__40618\
        );

    \I__10151\ : Odrv4
    port map (
            O => \N__40627\,
            I => \N_311_0\
        );

    \I__10150\ : Odrv4
    port map (
            O => \N__40624\,
            I => \N_311_0\
        );

    \I__10149\ : Odrv4
    port map (
            O => \N__40621\,
            I => \N_311_0\
        );

    \I__10148\ : Odrv4
    port map (
            O => \N__40618\,
            I => \N_311_0\
        );

    \I__10147\ : CascadeMux
    port map (
            O => \N__40609\,
            I => \N__40604\
        );

    \I__10146\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40601\
        );

    \I__10145\ : InMux
    port map (
            O => \N__40607\,
            I => \N__40595\
        );

    \I__10144\ : InMux
    port map (
            O => \N__40604\,
            I => \N__40592\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__40601\,
            I => \N__40589\
        );

    \I__10142\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40586\
        );

    \I__10141\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40583\
        );

    \I__10140\ : InMux
    port map (
            O => \N__40598\,
            I => \N__40579\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__40595\,
            I => \N__40576\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__40592\,
            I => \N__40571\
        );

    \I__10137\ : Span4Mux_h
    port map (
            O => \N__40589\,
            I => \N__40566\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__40586\,
            I => \N__40566\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__40583\,
            I => \N__40563\
        );

    \I__10134\ : CascadeMux
    port map (
            O => \N__40582\,
            I => \N__40560\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__40579\,
            I => \N__40557\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__40576\,
            I => \N__40554\
        );

    \I__10131\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40551\
        );

    \I__10130\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40548\
        );

    \I__10129\ : Span4Mux_v
    port map (
            O => \N__40571\,
            I => \N__40545\
        );

    \I__10128\ : Span4Mux_v
    port map (
            O => \N__40566\,
            I => \N__40540\
        );

    \I__10127\ : Span4Mux_v
    port map (
            O => \N__40563\,
            I => \N__40540\
        );

    \I__10126\ : InMux
    port map (
            O => \N__40560\,
            I => \N__40537\
        );

    \I__10125\ : Span12Mux_v
    port map (
            O => \N__40557\,
            I => \N__40534\
        );

    \I__10124\ : Sp12to4
    port map (
            O => \N__40554\,
            I => \N__40527\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__40551\,
            I => \N__40527\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__40548\,
            I => \N__40527\
        );

    \I__10121\ : Sp12to4
    port map (
            O => \N__40545\,
            I => \N__40522\
        );

    \I__10120\ : Sp12to4
    port map (
            O => \N__40540\,
            I => \N__40522\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__40537\,
            I => \N__40519\
        );

    \I__10118\ : Span12Mux_h
    port map (
            O => \N__40534\,
            I => \N__40516\
        );

    \I__10117\ : Span12Mux_v
    port map (
            O => \N__40527\,
            I => \N__40513\
        );

    \I__10116\ : Span12Mux_h
    port map (
            O => \N__40522\,
            I => \N__40508\
        );

    \I__10115\ : Span12Mux_v
    port map (
            O => \N__40519\,
            I => \N__40508\
        );

    \I__10114\ : Odrv12
    port map (
            O => \N__40516\,
            I => port_data_c_5
        );

    \I__10113\ : Odrv12
    port map (
            O => \N__40513\,
            I => port_data_c_5
        );

    \I__10112\ : Odrv12
    port map (
            O => \N__40508\,
            I => port_data_c_5
        );

    \I__10111\ : InMux
    port map (
            O => \N__40501\,
            I => \N__40498\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__40498\,
            I => \N__40495\
        );

    \I__10109\ : Odrv4
    port map (
            O => \N__40495\,
            I => \un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0\
        );

    \I__10108\ : IoInMux
    port map (
            O => \N__40492\,
            I => \N__40489\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__40489\,
            I => \N__40485\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__40488\,
            I => \N__40482\
        );

    \I__10105\ : IoSpan4Mux
    port map (
            O => \N__40485\,
            I => \N__40479\
        );

    \I__10104\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40476\
        );

    \I__10103\ : Span4Mux_s3_h
    port map (
            O => \N__40479\,
            I => \N__40473\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__40476\,
            I => \N__40470\
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__40473\,
            I => \M_this_ext_address_qZ0Z_13\
        );

    \I__10100\ : Odrv4
    port map (
            O => \N__40470\,
            I => \M_this_ext_address_qZ0Z_13\
        );

    \I__10099\ : ClkMux
    port map (
            O => \N__40465\,
            I => \N__39928\
        );

    \I__10098\ : ClkMux
    port map (
            O => \N__40464\,
            I => \N__39928\
        );

    \I__10097\ : ClkMux
    port map (
            O => \N__40463\,
            I => \N__39928\
        );

    \I__10096\ : ClkMux
    port map (
            O => \N__40462\,
            I => \N__39928\
        );

    \I__10095\ : ClkMux
    port map (
            O => \N__40461\,
            I => \N__39928\
        );

    \I__10094\ : ClkMux
    port map (
            O => \N__40460\,
            I => \N__39928\
        );

    \I__10093\ : ClkMux
    port map (
            O => \N__40459\,
            I => \N__39928\
        );

    \I__10092\ : ClkMux
    port map (
            O => \N__40458\,
            I => \N__39928\
        );

    \I__10091\ : ClkMux
    port map (
            O => \N__40457\,
            I => \N__39928\
        );

    \I__10090\ : ClkMux
    port map (
            O => \N__40456\,
            I => \N__39928\
        );

    \I__10089\ : ClkMux
    port map (
            O => \N__40455\,
            I => \N__39928\
        );

    \I__10088\ : ClkMux
    port map (
            O => \N__40454\,
            I => \N__39928\
        );

    \I__10087\ : ClkMux
    port map (
            O => \N__40453\,
            I => \N__39928\
        );

    \I__10086\ : ClkMux
    port map (
            O => \N__40452\,
            I => \N__39928\
        );

    \I__10085\ : ClkMux
    port map (
            O => \N__40451\,
            I => \N__39928\
        );

    \I__10084\ : ClkMux
    port map (
            O => \N__40450\,
            I => \N__39928\
        );

    \I__10083\ : ClkMux
    port map (
            O => \N__40449\,
            I => \N__39928\
        );

    \I__10082\ : ClkMux
    port map (
            O => \N__40448\,
            I => \N__39928\
        );

    \I__10081\ : ClkMux
    port map (
            O => \N__40447\,
            I => \N__39928\
        );

    \I__10080\ : ClkMux
    port map (
            O => \N__40446\,
            I => \N__39928\
        );

    \I__10079\ : ClkMux
    port map (
            O => \N__40445\,
            I => \N__39928\
        );

    \I__10078\ : ClkMux
    port map (
            O => \N__40444\,
            I => \N__39928\
        );

    \I__10077\ : ClkMux
    port map (
            O => \N__40443\,
            I => \N__39928\
        );

    \I__10076\ : ClkMux
    port map (
            O => \N__40442\,
            I => \N__39928\
        );

    \I__10075\ : ClkMux
    port map (
            O => \N__40441\,
            I => \N__39928\
        );

    \I__10074\ : ClkMux
    port map (
            O => \N__40440\,
            I => \N__39928\
        );

    \I__10073\ : ClkMux
    port map (
            O => \N__40439\,
            I => \N__39928\
        );

    \I__10072\ : ClkMux
    port map (
            O => \N__40438\,
            I => \N__39928\
        );

    \I__10071\ : ClkMux
    port map (
            O => \N__40437\,
            I => \N__39928\
        );

    \I__10070\ : ClkMux
    port map (
            O => \N__40436\,
            I => \N__39928\
        );

    \I__10069\ : ClkMux
    port map (
            O => \N__40435\,
            I => \N__39928\
        );

    \I__10068\ : ClkMux
    port map (
            O => \N__40434\,
            I => \N__39928\
        );

    \I__10067\ : ClkMux
    port map (
            O => \N__40433\,
            I => \N__39928\
        );

    \I__10066\ : ClkMux
    port map (
            O => \N__40432\,
            I => \N__39928\
        );

    \I__10065\ : ClkMux
    port map (
            O => \N__40431\,
            I => \N__39928\
        );

    \I__10064\ : ClkMux
    port map (
            O => \N__40430\,
            I => \N__39928\
        );

    \I__10063\ : ClkMux
    port map (
            O => \N__40429\,
            I => \N__39928\
        );

    \I__10062\ : ClkMux
    port map (
            O => \N__40428\,
            I => \N__39928\
        );

    \I__10061\ : ClkMux
    port map (
            O => \N__40427\,
            I => \N__39928\
        );

    \I__10060\ : ClkMux
    port map (
            O => \N__40426\,
            I => \N__39928\
        );

    \I__10059\ : ClkMux
    port map (
            O => \N__40425\,
            I => \N__39928\
        );

    \I__10058\ : ClkMux
    port map (
            O => \N__40424\,
            I => \N__39928\
        );

    \I__10057\ : ClkMux
    port map (
            O => \N__40423\,
            I => \N__39928\
        );

    \I__10056\ : ClkMux
    port map (
            O => \N__40422\,
            I => \N__39928\
        );

    \I__10055\ : ClkMux
    port map (
            O => \N__40421\,
            I => \N__39928\
        );

    \I__10054\ : ClkMux
    port map (
            O => \N__40420\,
            I => \N__39928\
        );

    \I__10053\ : ClkMux
    port map (
            O => \N__40419\,
            I => \N__39928\
        );

    \I__10052\ : ClkMux
    port map (
            O => \N__40418\,
            I => \N__39928\
        );

    \I__10051\ : ClkMux
    port map (
            O => \N__40417\,
            I => \N__39928\
        );

    \I__10050\ : ClkMux
    port map (
            O => \N__40416\,
            I => \N__39928\
        );

    \I__10049\ : ClkMux
    port map (
            O => \N__40415\,
            I => \N__39928\
        );

    \I__10048\ : ClkMux
    port map (
            O => \N__40414\,
            I => \N__39928\
        );

    \I__10047\ : ClkMux
    port map (
            O => \N__40413\,
            I => \N__39928\
        );

    \I__10046\ : ClkMux
    port map (
            O => \N__40412\,
            I => \N__39928\
        );

    \I__10045\ : ClkMux
    port map (
            O => \N__40411\,
            I => \N__39928\
        );

    \I__10044\ : ClkMux
    port map (
            O => \N__40410\,
            I => \N__39928\
        );

    \I__10043\ : ClkMux
    port map (
            O => \N__40409\,
            I => \N__39928\
        );

    \I__10042\ : ClkMux
    port map (
            O => \N__40408\,
            I => \N__39928\
        );

    \I__10041\ : ClkMux
    port map (
            O => \N__40407\,
            I => \N__39928\
        );

    \I__10040\ : ClkMux
    port map (
            O => \N__40406\,
            I => \N__39928\
        );

    \I__10039\ : ClkMux
    port map (
            O => \N__40405\,
            I => \N__39928\
        );

    \I__10038\ : ClkMux
    port map (
            O => \N__40404\,
            I => \N__39928\
        );

    \I__10037\ : ClkMux
    port map (
            O => \N__40403\,
            I => \N__39928\
        );

    \I__10036\ : ClkMux
    port map (
            O => \N__40402\,
            I => \N__39928\
        );

    \I__10035\ : ClkMux
    port map (
            O => \N__40401\,
            I => \N__39928\
        );

    \I__10034\ : ClkMux
    port map (
            O => \N__40400\,
            I => \N__39928\
        );

    \I__10033\ : ClkMux
    port map (
            O => \N__40399\,
            I => \N__39928\
        );

    \I__10032\ : ClkMux
    port map (
            O => \N__40398\,
            I => \N__39928\
        );

    \I__10031\ : ClkMux
    port map (
            O => \N__40397\,
            I => \N__39928\
        );

    \I__10030\ : ClkMux
    port map (
            O => \N__40396\,
            I => \N__39928\
        );

    \I__10029\ : ClkMux
    port map (
            O => \N__40395\,
            I => \N__39928\
        );

    \I__10028\ : ClkMux
    port map (
            O => \N__40394\,
            I => \N__39928\
        );

    \I__10027\ : ClkMux
    port map (
            O => \N__40393\,
            I => \N__39928\
        );

    \I__10026\ : ClkMux
    port map (
            O => \N__40392\,
            I => \N__39928\
        );

    \I__10025\ : ClkMux
    port map (
            O => \N__40391\,
            I => \N__39928\
        );

    \I__10024\ : ClkMux
    port map (
            O => \N__40390\,
            I => \N__39928\
        );

    \I__10023\ : ClkMux
    port map (
            O => \N__40389\,
            I => \N__39928\
        );

    \I__10022\ : ClkMux
    port map (
            O => \N__40388\,
            I => \N__39928\
        );

    \I__10021\ : ClkMux
    port map (
            O => \N__40387\,
            I => \N__39928\
        );

    \I__10020\ : ClkMux
    port map (
            O => \N__40386\,
            I => \N__39928\
        );

    \I__10019\ : ClkMux
    port map (
            O => \N__40385\,
            I => \N__39928\
        );

    \I__10018\ : ClkMux
    port map (
            O => \N__40384\,
            I => \N__39928\
        );

    \I__10017\ : ClkMux
    port map (
            O => \N__40383\,
            I => \N__39928\
        );

    \I__10016\ : ClkMux
    port map (
            O => \N__40382\,
            I => \N__39928\
        );

    \I__10015\ : ClkMux
    port map (
            O => \N__40381\,
            I => \N__39928\
        );

    \I__10014\ : ClkMux
    port map (
            O => \N__40380\,
            I => \N__39928\
        );

    \I__10013\ : ClkMux
    port map (
            O => \N__40379\,
            I => \N__39928\
        );

    \I__10012\ : ClkMux
    port map (
            O => \N__40378\,
            I => \N__39928\
        );

    \I__10011\ : ClkMux
    port map (
            O => \N__40377\,
            I => \N__39928\
        );

    \I__10010\ : ClkMux
    port map (
            O => \N__40376\,
            I => \N__39928\
        );

    \I__10009\ : ClkMux
    port map (
            O => \N__40375\,
            I => \N__39928\
        );

    \I__10008\ : ClkMux
    port map (
            O => \N__40374\,
            I => \N__39928\
        );

    \I__10007\ : ClkMux
    port map (
            O => \N__40373\,
            I => \N__39928\
        );

    \I__10006\ : ClkMux
    port map (
            O => \N__40372\,
            I => \N__39928\
        );

    \I__10005\ : ClkMux
    port map (
            O => \N__40371\,
            I => \N__39928\
        );

    \I__10004\ : ClkMux
    port map (
            O => \N__40370\,
            I => \N__39928\
        );

    \I__10003\ : ClkMux
    port map (
            O => \N__40369\,
            I => \N__39928\
        );

    \I__10002\ : ClkMux
    port map (
            O => \N__40368\,
            I => \N__39928\
        );

    \I__10001\ : ClkMux
    port map (
            O => \N__40367\,
            I => \N__39928\
        );

    \I__10000\ : ClkMux
    port map (
            O => \N__40366\,
            I => \N__39928\
        );

    \I__9999\ : ClkMux
    port map (
            O => \N__40365\,
            I => \N__39928\
        );

    \I__9998\ : ClkMux
    port map (
            O => \N__40364\,
            I => \N__39928\
        );

    \I__9997\ : ClkMux
    port map (
            O => \N__40363\,
            I => \N__39928\
        );

    \I__9996\ : ClkMux
    port map (
            O => \N__40362\,
            I => \N__39928\
        );

    \I__9995\ : ClkMux
    port map (
            O => \N__40361\,
            I => \N__39928\
        );

    \I__9994\ : ClkMux
    port map (
            O => \N__40360\,
            I => \N__39928\
        );

    \I__9993\ : ClkMux
    port map (
            O => \N__40359\,
            I => \N__39928\
        );

    \I__9992\ : ClkMux
    port map (
            O => \N__40358\,
            I => \N__39928\
        );

    \I__9991\ : ClkMux
    port map (
            O => \N__40357\,
            I => \N__39928\
        );

    \I__9990\ : ClkMux
    port map (
            O => \N__40356\,
            I => \N__39928\
        );

    \I__9989\ : ClkMux
    port map (
            O => \N__40355\,
            I => \N__39928\
        );

    \I__9988\ : ClkMux
    port map (
            O => \N__40354\,
            I => \N__39928\
        );

    \I__9987\ : ClkMux
    port map (
            O => \N__40353\,
            I => \N__39928\
        );

    \I__9986\ : ClkMux
    port map (
            O => \N__40352\,
            I => \N__39928\
        );

    \I__9985\ : ClkMux
    port map (
            O => \N__40351\,
            I => \N__39928\
        );

    \I__9984\ : ClkMux
    port map (
            O => \N__40350\,
            I => \N__39928\
        );

    \I__9983\ : ClkMux
    port map (
            O => \N__40349\,
            I => \N__39928\
        );

    \I__9982\ : ClkMux
    port map (
            O => \N__40348\,
            I => \N__39928\
        );

    \I__9981\ : ClkMux
    port map (
            O => \N__40347\,
            I => \N__39928\
        );

    \I__9980\ : ClkMux
    port map (
            O => \N__40346\,
            I => \N__39928\
        );

    \I__9979\ : ClkMux
    port map (
            O => \N__40345\,
            I => \N__39928\
        );

    \I__9978\ : ClkMux
    port map (
            O => \N__40344\,
            I => \N__39928\
        );

    \I__9977\ : ClkMux
    port map (
            O => \N__40343\,
            I => \N__39928\
        );

    \I__9976\ : ClkMux
    port map (
            O => \N__40342\,
            I => \N__39928\
        );

    \I__9975\ : ClkMux
    port map (
            O => \N__40341\,
            I => \N__39928\
        );

    \I__9974\ : ClkMux
    port map (
            O => \N__40340\,
            I => \N__39928\
        );

    \I__9973\ : ClkMux
    port map (
            O => \N__40339\,
            I => \N__39928\
        );

    \I__9972\ : ClkMux
    port map (
            O => \N__40338\,
            I => \N__39928\
        );

    \I__9971\ : ClkMux
    port map (
            O => \N__40337\,
            I => \N__39928\
        );

    \I__9970\ : ClkMux
    port map (
            O => \N__40336\,
            I => \N__39928\
        );

    \I__9969\ : ClkMux
    port map (
            O => \N__40335\,
            I => \N__39928\
        );

    \I__9968\ : ClkMux
    port map (
            O => \N__40334\,
            I => \N__39928\
        );

    \I__9967\ : ClkMux
    port map (
            O => \N__40333\,
            I => \N__39928\
        );

    \I__9966\ : ClkMux
    port map (
            O => \N__40332\,
            I => \N__39928\
        );

    \I__9965\ : ClkMux
    port map (
            O => \N__40331\,
            I => \N__39928\
        );

    \I__9964\ : ClkMux
    port map (
            O => \N__40330\,
            I => \N__39928\
        );

    \I__9963\ : ClkMux
    port map (
            O => \N__40329\,
            I => \N__39928\
        );

    \I__9962\ : ClkMux
    port map (
            O => \N__40328\,
            I => \N__39928\
        );

    \I__9961\ : ClkMux
    port map (
            O => \N__40327\,
            I => \N__39928\
        );

    \I__9960\ : ClkMux
    port map (
            O => \N__40326\,
            I => \N__39928\
        );

    \I__9959\ : ClkMux
    port map (
            O => \N__40325\,
            I => \N__39928\
        );

    \I__9958\ : ClkMux
    port map (
            O => \N__40324\,
            I => \N__39928\
        );

    \I__9957\ : ClkMux
    port map (
            O => \N__40323\,
            I => \N__39928\
        );

    \I__9956\ : ClkMux
    port map (
            O => \N__40322\,
            I => \N__39928\
        );

    \I__9955\ : ClkMux
    port map (
            O => \N__40321\,
            I => \N__39928\
        );

    \I__9954\ : ClkMux
    port map (
            O => \N__40320\,
            I => \N__39928\
        );

    \I__9953\ : ClkMux
    port map (
            O => \N__40319\,
            I => \N__39928\
        );

    \I__9952\ : ClkMux
    port map (
            O => \N__40318\,
            I => \N__39928\
        );

    \I__9951\ : ClkMux
    port map (
            O => \N__40317\,
            I => \N__39928\
        );

    \I__9950\ : ClkMux
    port map (
            O => \N__40316\,
            I => \N__39928\
        );

    \I__9949\ : ClkMux
    port map (
            O => \N__40315\,
            I => \N__39928\
        );

    \I__9948\ : ClkMux
    port map (
            O => \N__40314\,
            I => \N__39928\
        );

    \I__9947\ : ClkMux
    port map (
            O => \N__40313\,
            I => \N__39928\
        );

    \I__9946\ : ClkMux
    port map (
            O => \N__40312\,
            I => \N__39928\
        );

    \I__9945\ : ClkMux
    port map (
            O => \N__40311\,
            I => \N__39928\
        );

    \I__9944\ : ClkMux
    port map (
            O => \N__40310\,
            I => \N__39928\
        );

    \I__9943\ : ClkMux
    port map (
            O => \N__40309\,
            I => \N__39928\
        );

    \I__9942\ : ClkMux
    port map (
            O => \N__40308\,
            I => \N__39928\
        );

    \I__9941\ : ClkMux
    port map (
            O => \N__40307\,
            I => \N__39928\
        );

    \I__9940\ : ClkMux
    port map (
            O => \N__40306\,
            I => \N__39928\
        );

    \I__9939\ : ClkMux
    port map (
            O => \N__40305\,
            I => \N__39928\
        );

    \I__9938\ : ClkMux
    port map (
            O => \N__40304\,
            I => \N__39928\
        );

    \I__9937\ : ClkMux
    port map (
            O => \N__40303\,
            I => \N__39928\
        );

    \I__9936\ : ClkMux
    port map (
            O => \N__40302\,
            I => \N__39928\
        );

    \I__9935\ : ClkMux
    port map (
            O => \N__40301\,
            I => \N__39928\
        );

    \I__9934\ : ClkMux
    port map (
            O => \N__40300\,
            I => \N__39928\
        );

    \I__9933\ : ClkMux
    port map (
            O => \N__40299\,
            I => \N__39928\
        );

    \I__9932\ : ClkMux
    port map (
            O => \N__40298\,
            I => \N__39928\
        );

    \I__9931\ : ClkMux
    port map (
            O => \N__40297\,
            I => \N__39928\
        );

    \I__9930\ : ClkMux
    port map (
            O => \N__40296\,
            I => \N__39928\
        );

    \I__9929\ : ClkMux
    port map (
            O => \N__40295\,
            I => \N__39928\
        );

    \I__9928\ : ClkMux
    port map (
            O => \N__40294\,
            I => \N__39928\
        );

    \I__9927\ : ClkMux
    port map (
            O => \N__40293\,
            I => \N__39928\
        );

    \I__9926\ : ClkMux
    port map (
            O => \N__40292\,
            I => \N__39928\
        );

    \I__9925\ : ClkMux
    port map (
            O => \N__40291\,
            I => \N__39928\
        );

    \I__9924\ : ClkMux
    port map (
            O => \N__40290\,
            I => \N__39928\
        );

    \I__9923\ : ClkMux
    port map (
            O => \N__40289\,
            I => \N__39928\
        );

    \I__9922\ : ClkMux
    port map (
            O => \N__40288\,
            I => \N__39928\
        );

    \I__9921\ : ClkMux
    port map (
            O => \N__40287\,
            I => \N__39928\
        );

    \I__9920\ : GlobalMux
    port map (
            O => \N__39928\,
            I => \N__39925\
        );

    \I__9919\ : gio2CtrlBuf
    port map (
            O => \N__39925\,
            I => clk_0_c_g
        );

    \I__9918\ : CascadeMux
    port map (
            O => \N__39922\,
            I => \N__39916\
        );

    \I__9917\ : CascadeMux
    port map (
            O => \N__39921\,
            I => \N__39905\
        );

    \I__9916\ : CascadeMux
    port map (
            O => \N__39920\,
            I => \N__39898\
        );

    \I__9915\ : CascadeMux
    port map (
            O => \N__39919\,
            I => \N__39886\
        );

    \I__9914\ : InMux
    port map (
            O => \N__39916\,
            I => \N__39878\
        );

    \I__9913\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39875\
        );

    \I__9912\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39872\
        );

    \I__9911\ : InMux
    port map (
            O => \N__39913\,
            I => \N__39869\
        );

    \I__9910\ : InMux
    port map (
            O => \N__39912\,
            I => \N__39866\
        );

    \I__9909\ : InMux
    port map (
            O => \N__39911\,
            I => \N__39863\
        );

    \I__9908\ : InMux
    port map (
            O => \N__39910\,
            I => \N__39858\
        );

    \I__9907\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39858\
        );

    \I__9906\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39855\
        );

    \I__9905\ : InMux
    port map (
            O => \N__39905\,
            I => \N__39852\
        );

    \I__9904\ : InMux
    port map (
            O => \N__39904\,
            I => \N__39849\
        );

    \I__9903\ : InMux
    port map (
            O => \N__39903\,
            I => \N__39846\
        );

    \I__9902\ : InMux
    port map (
            O => \N__39902\,
            I => \N__39841\
        );

    \I__9901\ : InMux
    port map (
            O => \N__39901\,
            I => \N__39841\
        );

    \I__9900\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39838\
        );

    \I__9899\ : InMux
    port map (
            O => \N__39897\,
            I => \N__39835\
        );

    \I__9898\ : InMux
    port map (
            O => \N__39896\,
            I => \N__39832\
        );

    \I__9897\ : InMux
    port map (
            O => \N__39895\,
            I => \N__39829\
        );

    \I__9896\ : InMux
    port map (
            O => \N__39894\,
            I => \N__39826\
        );

    \I__9895\ : InMux
    port map (
            O => \N__39893\,
            I => \N__39821\
        );

    \I__9894\ : InMux
    port map (
            O => \N__39892\,
            I => \N__39821\
        );

    \I__9893\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39818\
        );

    \I__9892\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39815\
        );

    \I__9891\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39812\
        );

    \I__9890\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39809\
        );

    \I__9889\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39804\
        );

    \I__9888\ : InMux
    port map (
            O => \N__39884\,
            I => \N__39804\
        );

    \I__9887\ : InMux
    port map (
            O => \N__39883\,
            I => \N__39801\
        );

    \I__9886\ : InMux
    port map (
            O => \N__39882\,
            I => \N__39796\
        );

    \I__9885\ : InMux
    port map (
            O => \N__39881\,
            I => \N__39796\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__39878\,
            I => \N__39751\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39748\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__39872\,
            I => \N__39745\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__39869\,
            I => \N__39742\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__39866\,
            I => \N__39739\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__39863\,
            I => \N__39736\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__39858\,
            I => \N__39733\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__39855\,
            I => \N__39730\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__39852\,
            I => \N__39727\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__39849\,
            I => \N__39724\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__39846\,
            I => \N__39721\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__39841\,
            I => \N__39718\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__39838\,
            I => \N__39715\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__39835\,
            I => \N__39712\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__39832\,
            I => \N__39709\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__39829\,
            I => \N__39706\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__39826\,
            I => \N__39703\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__39821\,
            I => \N__39700\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__39818\,
            I => \N__39697\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39694\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__39812\,
            I => \N__39691\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__39809\,
            I => \N__39688\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__39804\,
            I => \N__39685\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__39801\,
            I => \N__39682\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__39796\,
            I => \N__39679\
        );

    \I__9859\ : SRMux
    port map (
            O => \N__39795\,
            I => \N__39544\
        );

    \I__9858\ : SRMux
    port map (
            O => \N__39794\,
            I => \N__39544\
        );

    \I__9857\ : SRMux
    port map (
            O => \N__39793\,
            I => \N__39544\
        );

    \I__9856\ : SRMux
    port map (
            O => \N__39792\,
            I => \N__39544\
        );

    \I__9855\ : SRMux
    port map (
            O => \N__39791\,
            I => \N__39544\
        );

    \I__9854\ : SRMux
    port map (
            O => \N__39790\,
            I => \N__39544\
        );

    \I__9853\ : SRMux
    port map (
            O => \N__39789\,
            I => \N__39544\
        );

    \I__9852\ : SRMux
    port map (
            O => \N__39788\,
            I => \N__39544\
        );

    \I__9851\ : SRMux
    port map (
            O => \N__39787\,
            I => \N__39544\
        );

    \I__9850\ : SRMux
    port map (
            O => \N__39786\,
            I => \N__39544\
        );

    \I__9849\ : SRMux
    port map (
            O => \N__39785\,
            I => \N__39544\
        );

    \I__9848\ : SRMux
    port map (
            O => \N__39784\,
            I => \N__39544\
        );

    \I__9847\ : SRMux
    port map (
            O => \N__39783\,
            I => \N__39544\
        );

    \I__9846\ : SRMux
    port map (
            O => \N__39782\,
            I => \N__39544\
        );

    \I__9845\ : SRMux
    port map (
            O => \N__39781\,
            I => \N__39544\
        );

    \I__9844\ : SRMux
    port map (
            O => \N__39780\,
            I => \N__39544\
        );

    \I__9843\ : SRMux
    port map (
            O => \N__39779\,
            I => \N__39544\
        );

    \I__9842\ : SRMux
    port map (
            O => \N__39778\,
            I => \N__39544\
        );

    \I__9841\ : SRMux
    port map (
            O => \N__39777\,
            I => \N__39544\
        );

    \I__9840\ : SRMux
    port map (
            O => \N__39776\,
            I => \N__39544\
        );

    \I__9839\ : SRMux
    port map (
            O => \N__39775\,
            I => \N__39544\
        );

    \I__9838\ : SRMux
    port map (
            O => \N__39774\,
            I => \N__39544\
        );

    \I__9837\ : SRMux
    port map (
            O => \N__39773\,
            I => \N__39544\
        );

    \I__9836\ : SRMux
    port map (
            O => \N__39772\,
            I => \N__39544\
        );

    \I__9835\ : SRMux
    port map (
            O => \N__39771\,
            I => \N__39544\
        );

    \I__9834\ : SRMux
    port map (
            O => \N__39770\,
            I => \N__39544\
        );

    \I__9833\ : SRMux
    port map (
            O => \N__39769\,
            I => \N__39544\
        );

    \I__9832\ : SRMux
    port map (
            O => \N__39768\,
            I => \N__39544\
        );

    \I__9831\ : SRMux
    port map (
            O => \N__39767\,
            I => \N__39544\
        );

    \I__9830\ : SRMux
    port map (
            O => \N__39766\,
            I => \N__39544\
        );

    \I__9829\ : SRMux
    port map (
            O => \N__39765\,
            I => \N__39544\
        );

    \I__9828\ : SRMux
    port map (
            O => \N__39764\,
            I => \N__39544\
        );

    \I__9827\ : SRMux
    port map (
            O => \N__39763\,
            I => \N__39544\
        );

    \I__9826\ : SRMux
    port map (
            O => \N__39762\,
            I => \N__39544\
        );

    \I__9825\ : SRMux
    port map (
            O => \N__39761\,
            I => \N__39544\
        );

    \I__9824\ : SRMux
    port map (
            O => \N__39760\,
            I => \N__39544\
        );

    \I__9823\ : SRMux
    port map (
            O => \N__39759\,
            I => \N__39544\
        );

    \I__9822\ : SRMux
    port map (
            O => \N__39758\,
            I => \N__39544\
        );

    \I__9821\ : SRMux
    port map (
            O => \N__39757\,
            I => \N__39544\
        );

    \I__9820\ : SRMux
    port map (
            O => \N__39756\,
            I => \N__39544\
        );

    \I__9819\ : SRMux
    port map (
            O => \N__39755\,
            I => \N__39544\
        );

    \I__9818\ : SRMux
    port map (
            O => \N__39754\,
            I => \N__39544\
        );

    \I__9817\ : Glb2LocalMux
    port map (
            O => \N__39751\,
            I => \N__39544\
        );

    \I__9816\ : Glb2LocalMux
    port map (
            O => \N__39748\,
            I => \N__39544\
        );

    \I__9815\ : Glb2LocalMux
    port map (
            O => \N__39745\,
            I => \N__39544\
        );

    \I__9814\ : Glb2LocalMux
    port map (
            O => \N__39742\,
            I => \N__39544\
        );

    \I__9813\ : Glb2LocalMux
    port map (
            O => \N__39739\,
            I => \N__39544\
        );

    \I__9812\ : Glb2LocalMux
    port map (
            O => \N__39736\,
            I => \N__39544\
        );

    \I__9811\ : Glb2LocalMux
    port map (
            O => \N__39733\,
            I => \N__39544\
        );

    \I__9810\ : Glb2LocalMux
    port map (
            O => \N__39730\,
            I => \N__39544\
        );

    \I__9809\ : Glb2LocalMux
    port map (
            O => \N__39727\,
            I => \N__39544\
        );

    \I__9808\ : Glb2LocalMux
    port map (
            O => \N__39724\,
            I => \N__39544\
        );

    \I__9807\ : Glb2LocalMux
    port map (
            O => \N__39721\,
            I => \N__39544\
        );

    \I__9806\ : Glb2LocalMux
    port map (
            O => \N__39718\,
            I => \N__39544\
        );

    \I__9805\ : Glb2LocalMux
    port map (
            O => \N__39715\,
            I => \N__39544\
        );

    \I__9804\ : Glb2LocalMux
    port map (
            O => \N__39712\,
            I => \N__39544\
        );

    \I__9803\ : Glb2LocalMux
    port map (
            O => \N__39709\,
            I => \N__39544\
        );

    \I__9802\ : Glb2LocalMux
    port map (
            O => \N__39706\,
            I => \N__39544\
        );

    \I__9801\ : Glb2LocalMux
    port map (
            O => \N__39703\,
            I => \N__39544\
        );

    \I__9800\ : Glb2LocalMux
    port map (
            O => \N__39700\,
            I => \N__39544\
        );

    \I__9799\ : Glb2LocalMux
    port map (
            O => \N__39697\,
            I => \N__39544\
        );

    \I__9798\ : Glb2LocalMux
    port map (
            O => \N__39694\,
            I => \N__39544\
        );

    \I__9797\ : Glb2LocalMux
    port map (
            O => \N__39691\,
            I => \N__39544\
        );

    \I__9796\ : Glb2LocalMux
    port map (
            O => \N__39688\,
            I => \N__39544\
        );

    \I__9795\ : Glb2LocalMux
    port map (
            O => \N__39685\,
            I => \N__39544\
        );

    \I__9794\ : Glb2LocalMux
    port map (
            O => \N__39682\,
            I => \N__39544\
        );

    \I__9793\ : Glb2LocalMux
    port map (
            O => \N__39679\,
            I => \N__39544\
        );

    \I__9792\ : GlobalMux
    port map (
            O => \N__39544\,
            I => \N__39541\
        );

    \I__9791\ : gio2CtrlBuf
    port map (
            O => \N__39541\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__9790\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39535\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__39535\,
            I => \N__39532\
        );

    \I__9788\ : Odrv4
    port map (
            O => \N__39532\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__9787\ : InMux
    port map (
            O => \N__39529\,
            I => \N__39526\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__39526\,
            I => \N__39523\
        );

    \I__9785\ : Span4Mux_v
    port map (
            O => \N__39523\,
            I => \N__39520\
        );

    \I__9784\ : Odrv4
    port map (
            O => \N__39520\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_12\
        );

    \I__9783\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39513\
        );

    \I__9782\ : CascadeMux
    port map (
            O => \N__39516\,
            I => \N__39510\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__39513\,
            I => \N__39507\
        );

    \I__9780\ : InMux
    port map (
            O => \N__39510\,
            I => \N__39502\
        );

    \I__9779\ : Span4Mux_h
    port map (
            O => \N__39507\,
            I => \N__39499\
        );

    \I__9778\ : InMux
    port map (
            O => \N__39506\,
            I => \N__39494\
        );

    \I__9777\ : CascadeMux
    port map (
            O => \N__39505\,
            I => \N__39491\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__39502\,
            I => \N__39488\
        );

    \I__9775\ : Span4Mux_v
    port map (
            O => \N__39499\,
            I => \N__39485\
        );

    \I__9774\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39482\
        );

    \I__9773\ : InMux
    port map (
            O => \N__39497\,
            I => \N__39479\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__39494\,
            I => \N__39475\
        );

    \I__9771\ : InMux
    port map (
            O => \N__39491\,
            I => \N__39472\
        );

    \I__9770\ : Span4Mux_v
    port map (
            O => \N__39488\,
            I => \N__39469\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__39485\,
            I => \N__39464\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__39482\,
            I => \N__39464\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__39479\,
            I => \N__39461\
        );

    \I__9766\ : InMux
    port map (
            O => \N__39478\,
            I => \N__39458\
        );

    \I__9765\ : Span4Mux_v
    port map (
            O => \N__39475\,
            I => \N__39455\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__39472\,
            I => \N__39451\
        );

    \I__9763\ : Span4Mux_v
    port map (
            O => \N__39469\,
            I => \N__39448\
        );

    \I__9762\ : Span4Mux_h
    port map (
            O => \N__39464\,
            I => \N__39441\
        );

    \I__9761\ : Span4Mux_v
    port map (
            O => \N__39461\,
            I => \N__39441\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__39458\,
            I => \N__39441\
        );

    \I__9759\ : Sp12to4
    port map (
            O => \N__39455\,
            I => \N__39437\
        );

    \I__9758\ : InMux
    port map (
            O => \N__39454\,
            I => \N__39434\
        );

    \I__9757\ : Span4Mux_h
    port map (
            O => \N__39451\,
            I => \N__39431\
        );

    \I__9756\ : Span4Mux_v
    port map (
            O => \N__39448\,
            I => \N__39426\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__39441\,
            I => \N__39426\
        );

    \I__9754\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39423\
        );

    \I__9753\ : Span12Mux_h
    port map (
            O => \N__39437\,
            I => \N__39420\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__39434\,
            I => \N__39417\
        );

    \I__9751\ : Span4Mux_v
    port map (
            O => \N__39431\,
            I => \N__39414\
        );

    \I__9750\ : Span4Mux_h
    port map (
            O => \N__39426\,
            I => \N__39411\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__39423\,
            I => \N__39408\
        );

    \I__9748\ : Span12Mux_v
    port map (
            O => \N__39420\,
            I => \N__39405\
        );

    \I__9747\ : Span12Mux_h
    port map (
            O => \N__39417\,
            I => \N__39402\
        );

    \I__9746\ : Span4Mux_v
    port map (
            O => \N__39414\,
            I => \N__39399\
        );

    \I__9745\ : Span4Mux_v
    port map (
            O => \N__39411\,
            I => \N__39394\
        );

    \I__9744\ : Span4Mux_h
    port map (
            O => \N__39408\,
            I => \N__39394\
        );

    \I__9743\ : Odrv12
    port map (
            O => \N__39405\,
            I => port_data_c_3
        );

    \I__9742\ : Odrv12
    port map (
            O => \N__39402\,
            I => port_data_c_3
        );

    \I__9741\ : Odrv4
    port map (
            O => \N__39399\,
            I => port_data_c_3
        );

    \I__9740\ : Odrv4
    port map (
            O => \N__39394\,
            I => port_data_c_3
        );

    \I__9739\ : CEMux
    port map (
            O => \N__39385\,
            I => \N__39381\
        );

    \I__9738\ : CEMux
    port map (
            O => \N__39384\,
            I => \N__39378\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__39381\,
            I => \N__39365\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__39378\,
            I => \N__39362\
        );

    \I__9735\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39355\
        );

    \I__9734\ : InMux
    port map (
            O => \N__39376\,
            I => \N__39355\
        );

    \I__9733\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39355\
        );

    \I__9732\ : InMux
    port map (
            O => \N__39374\,
            I => \N__39350\
        );

    \I__9731\ : InMux
    port map (
            O => \N__39373\,
            I => \N__39350\
        );

    \I__9730\ : InMux
    port map (
            O => \N__39372\,
            I => \N__39343\
        );

    \I__9729\ : InMux
    port map (
            O => \N__39371\,
            I => \N__39336\
        );

    \I__9728\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39336\
        );

    \I__9727\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39336\
        );

    \I__9726\ : InMux
    port map (
            O => \N__39368\,
            I => \N__39330\
        );

    \I__9725\ : Span4Mux_h
    port map (
            O => \N__39365\,
            I => \N__39325\
        );

    \I__9724\ : Span4Mux_v
    port map (
            O => \N__39362\,
            I => \N__39320\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__39355\,
            I => \N__39320\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__39350\,
            I => \N__39309\
        );

    \I__9721\ : InMux
    port map (
            O => \N__39349\,
            I => \N__39298\
        );

    \I__9720\ : InMux
    port map (
            O => \N__39348\,
            I => \N__39298\
        );

    \I__9719\ : InMux
    port map (
            O => \N__39347\,
            I => \N__39298\
        );

    \I__9718\ : InMux
    port map (
            O => \N__39346\,
            I => \N__39298\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__39343\,
            I => \N__39293\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__39336\,
            I => \N__39293\
        );

    \I__9715\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39286\
        );

    \I__9714\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39286\
        );

    \I__9713\ : InMux
    port map (
            O => \N__39333\,
            I => \N__39286\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__39330\,
            I => \N__39283\
        );

    \I__9711\ : InMux
    port map (
            O => \N__39329\,
            I => \N__39280\
        );

    \I__9710\ : InMux
    port map (
            O => \N__39328\,
            I => \N__39277\
        );

    \I__9709\ : Span4Mux_v
    port map (
            O => \N__39325\,
            I => \N__39272\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__39320\,
            I => \N__39272\
        );

    \I__9707\ : InMux
    port map (
            O => \N__39319\,
            I => \N__39266\
        );

    \I__9706\ : InMux
    port map (
            O => \N__39318\,
            I => \N__39263\
        );

    \I__9705\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39258\
        );

    \I__9704\ : InMux
    port map (
            O => \N__39316\,
            I => \N__39258\
        );

    \I__9703\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39255\
        );

    \I__9702\ : InMux
    port map (
            O => \N__39314\,
            I => \N__39252\
        );

    \I__9701\ : InMux
    port map (
            O => \N__39313\,
            I => \N__39247\
        );

    \I__9700\ : InMux
    port map (
            O => \N__39312\,
            I => \N__39247\
        );

    \I__9699\ : Span4Mux_h
    port map (
            O => \N__39309\,
            I => \N__39244\
        );

    \I__9698\ : InMux
    port map (
            O => \N__39308\,
            I => \N__39241\
        );

    \I__9697\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39238\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__39298\,
            I => \N__39231\
        );

    \I__9695\ : Span4Mux_v
    port map (
            O => \N__39293\,
            I => \N__39231\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__39286\,
            I => \N__39231\
        );

    \I__9693\ : Span4Mux_v
    port map (
            O => \N__39283\,
            I => \N__39224\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__39280\,
            I => \N__39224\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__39277\,
            I => \N__39224\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__39272\,
            I => \N__39221\
        );

    \I__9689\ : InMux
    port map (
            O => \N__39271\,
            I => \N__39216\
        );

    \I__9688\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39216\
        );

    \I__9687\ : InMux
    port map (
            O => \N__39269\,
            I => \N__39213\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__39266\,
            I => \N__39210\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__39263\,
            I => \N__39193\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__39258\,
            I => \N__39193\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__39255\,
            I => \N__39193\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__39252\,
            I => \N__39193\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__39247\,
            I => \N__39193\
        );

    \I__9680\ : Sp12to4
    port map (
            O => \N__39244\,
            I => \N__39193\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__39241\,
            I => \N__39193\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__39238\,
            I => \N__39193\
        );

    \I__9677\ : Span4Mux_v
    port map (
            O => \N__39231\,
            I => \N__39190\
        );

    \I__9676\ : Span4Mux_v
    port map (
            O => \N__39224\,
            I => \N__39187\
        );

    \I__9675\ : Sp12to4
    port map (
            O => \N__39221\,
            I => \N__39178\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__39216\,
            I => \N__39178\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__39213\,
            I => \N__39178\
        );

    \I__9672\ : Span12Mux_h
    port map (
            O => \N__39210\,
            I => \N__39178\
        );

    \I__9671\ : Span12Mux_v
    port map (
            O => \N__39193\,
            I => \N__39175\
        );

    \I__9670\ : Span4Mux_h
    port map (
            O => \N__39190\,
            I => \N__39172\
        );

    \I__9669\ : Odrv4
    port map (
            O => \N__39187\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__9668\ : Odrv12
    port map (
            O => \N__39178\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__9667\ : Odrv12
    port map (
            O => \N__39175\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__9666\ : Odrv4
    port map (
            O => \N__39172\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__9665\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39160\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39157\
        );

    \I__9663\ : Odrv4
    port map (
            O => \N__39157\,
            I => \N_436\
        );

    \I__9662\ : InMux
    port map (
            O => \N__39154\,
            I => \N__39151\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__39151\,
            I => \M_this_oam_ram_read_data_30\
        );

    \I__9660\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39145\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__39145\,
            I => \N__39142\
        );

    \I__9658\ : Span4Mux_h
    port map (
            O => \N__39142\,
            I => \N__39139\
        );

    \I__9657\ : Span4Mux_h
    port map (
            O => \N__39139\,
            I => \N__39136\
        );

    \I__9656\ : Odrv4
    port map (
            O => \N__39136\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_30\
        );

    \I__9655\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39130\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__39130\,
            I => \N__39127\
        );

    \I__9653\ : Span4Mux_h
    port map (
            O => \N__39127\,
            I => \N__39124\
        );

    \I__9652\ : Odrv4
    port map (
            O => \N__39124\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__9651\ : InMux
    port map (
            O => \N__39121\,
            I => \N__39118\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__39118\,
            I => \N__39115\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__39115\,
            I => \N__39112\
        );

    \I__9648\ : Odrv4
    port map (
            O => \N__39112\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_9\
        );

    \I__9647\ : InMux
    port map (
            O => \N__39109\,
            I => \N__39106\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__39106\,
            I => \N_435\
        );

    \I__9645\ : InMux
    port map (
            O => \N__39103\,
            I => \N__39099\
        );

    \I__9644\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39096\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__39099\,
            I => \N__39093\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__39096\,
            I => \N__39087\
        );

    \I__9641\ : Span4Mux_h
    port map (
            O => \N__39093\,
            I => \N__39087\
        );

    \I__9640\ : InMux
    port map (
            O => \N__39092\,
            I => \N__39084\
        );

    \I__9639\ : Span4Mux_v
    port map (
            O => \N__39087\,
            I => \N__39078\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__39084\,
            I => \N__39075\
        );

    \I__9637\ : InMux
    port map (
            O => \N__39083\,
            I => \N__39068\
        );

    \I__9636\ : InMux
    port map (
            O => \N__39082\,
            I => \N__39068\
        );

    \I__9635\ : InMux
    port map (
            O => \N__39081\,
            I => \N__39068\
        );

    \I__9634\ : Odrv4
    port map (
            O => \N__39078\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__39075\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__39068\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__9631\ : InMux
    port map (
            O => \N__39061\,
            I => \N__39058\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__39058\,
            I => \N__39053\
        );

    \I__9629\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39050\
        );

    \I__9628\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39047\
        );

    \I__9627\ : Sp12to4
    port map (
            O => \N__39053\,
            I => \N__39041\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__39050\,
            I => \N__39041\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__39047\,
            I => \N__39038\
        );

    \I__9624\ : InMux
    port map (
            O => \N__39046\,
            I => \N__39035\
        );

    \I__9623\ : Span12Mux_v
    port map (
            O => \N__39041\,
            I => \N__39029\
        );

    \I__9622\ : Span4Mux_v
    port map (
            O => \N__39038\,
            I => \N__39024\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__39035\,
            I => \N__39024\
        );

    \I__9620\ : InMux
    port map (
            O => \N__39034\,
            I => \N__39017\
        );

    \I__9619\ : InMux
    port map (
            O => \N__39033\,
            I => \N__39017\
        );

    \I__9618\ : InMux
    port map (
            O => \N__39032\,
            I => \N__39017\
        );

    \I__9617\ : Odrv12
    port map (
            O => \N__39029\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__9616\ : Odrv4
    port map (
            O => \N__39024\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__39017\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__9614\ : InMux
    port map (
            O => \N__39010\,
            I => \N__39007\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__39007\,
            I => \N__39004\
        );

    \I__9612\ : Span12Mux_v
    port map (
            O => \N__39004\,
            I => \N__39001\
        );

    \I__9611\ : Odrv12
    port map (
            O => \N__39001\,
            I => \this_ppu.un1_oam_data_1_1\
        );

    \I__9610\ : InMux
    port map (
            O => \N__38998\,
            I => \N__38995\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__38995\,
            I => \this_spr_ram.mem_out_bus5_2\
        );

    \I__9608\ : InMux
    port map (
            O => \N__38992\,
            I => \N__38989\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__38989\,
            I => \N__38986\
        );

    \I__9606\ : Span4Mux_v
    port map (
            O => \N__38986\,
            I => \N__38983\
        );

    \I__9605\ : Odrv4
    port map (
            O => \N__38983\,
            I => \this_spr_ram.mem_out_bus1_2\
        );

    \I__9604\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38977\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__38977\,
            I => \N__38974\
        );

    \I__9602\ : Span4Mux_h
    port map (
            O => \N__38974\,
            I => \N__38971\
        );

    \I__9601\ : Sp12to4
    port map (
            O => \N__38971\,
            I => \N__38968\
        );

    \I__9600\ : Odrv12
    port map (
            O => \N__38968\,
            I => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\
        );

    \I__9599\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38962\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__38962\,
            I => \N__38959\
        );

    \I__9597\ : Odrv4
    port map (
            O => \N__38959\,
            I => \this_spr_ram.mem_out_bus5_0\
        );

    \I__9596\ : InMux
    port map (
            O => \N__38956\,
            I => \N__38953\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__38953\,
            I => \N__38950\
        );

    \I__9594\ : Span4Mux_v
    port map (
            O => \N__38950\,
            I => \N__38947\
        );

    \I__9593\ : Odrv4
    port map (
            O => \N__38947\,
            I => \this_spr_ram.mem_out_bus1_0\
        );

    \I__9592\ : InMux
    port map (
            O => \N__38944\,
            I => \N__38938\
        );

    \I__9591\ : InMux
    port map (
            O => \N__38943\,
            I => \N__38938\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__38938\,
            I => \N__38925\
        );

    \I__9589\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38920\
        );

    \I__9588\ : InMux
    port map (
            O => \N__38936\,
            I => \N__38920\
        );

    \I__9587\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38915\
        );

    \I__9586\ : InMux
    port map (
            O => \N__38934\,
            I => \N__38915\
        );

    \I__9585\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38911\
        );

    \I__9584\ : InMux
    port map (
            O => \N__38932\,
            I => \N__38908\
        );

    \I__9583\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38905\
        );

    \I__9582\ : InMux
    port map (
            O => \N__38930\,
            I => \N__38902\
        );

    \I__9581\ : InMux
    port map (
            O => \N__38929\,
            I => \N__38896\
        );

    \I__9580\ : InMux
    port map (
            O => \N__38928\,
            I => \N__38893\
        );

    \I__9579\ : Span4Mux_v
    port map (
            O => \N__38925\,
            I => \N__38886\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__38920\,
            I => \N__38886\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__38915\,
            I => \N__38886\
        );

    \I__9576\ : InMux
    port map (
            O => \N__38914\,
            I => \N__38883\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__38911\,
            I => \N__38880\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__38908\,
            I => \N__38873\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__38905\,
            I => \N__38873\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__38902\,
            I => \N__38873\
        );

    \I__9571\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38870\
        );

    \I__9570\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38867\
        );

    \I__9569\ : InMux
    port map (
            O => \N__38899\,
            I => \N__38864\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__38896\,
            I => \N__38859\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__38893\,
            I => \N__38859\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__38886\,
            I => \N__38856\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__38883\,
            I => \N__38853\
        );

    \I__9564\ : Span4Mux_h
    port map (
            O => \N__38880\,
            I => \N__38848\
        );

    \I__9563\ : Span4Mux_v
    port map (
            O => \N__38873\,
            I => \N__38848\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__38870\,
            I => \N__38845\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__38867\,
            I => \N__38842\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__38864\,
            I => \N__38837\
        );

    \I__9559\ : Span4Mux_v
    port map (
            O => \N__38859\,
            I => \N__38837\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__38856\,
            I => \N__38834\
        );

    \I__9557\ : Span12Mux_h
    port map (
            O => \N__38853\,
            I => \N__38831\
        );

    \I__9556\ : Span4Mux_h
    port map (
            O => \N__38848\,
            I => \N__38828\
        );

    \I__9555\ : Span12Mux_h
    port map (
            O => \N__38845\,
            I => \N__38825\
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__38842\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9553\ : Odrv4
    port map (
            O => \N__38837\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9552\ : Odrv4
    port map (
            O => \N__38834\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9551\ : Odrv12
    port map (
            O => \N__38831\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9550\ : Odrv4
    port map (
            O => \N__38828\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9549\ : Odrv12
    port map (
            O => \N__38825\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__9548\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38809\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__38809\,
            I => \N__38806\
        );

    \I__9546\ : Span12Mux_h
    port map (
            O => \N__38806\,
            I => \N__38803\
        );

    \I__9545\ : Odrv12
    port map (
            O => \N__38803\,
            I => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\
        );

    \I__9544\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38797\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__38797\,
            I => \N__38794\
        );

    \I__9542\ : Odrv4
    port map (
            O => \N__38794\,
            I => \un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0\
        );

    \I__9541\ : InMux
    port map (
            O => \N__38791\,
            I => \N__38788\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__38788\,
            I => \N__38785\
        );

    \I__9539\ : Span4Mux_v
    port map (
            O => \N__38785\,
            I => \N__38781\
        );

    \I__9538\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38776\
        );

    \I__9537\ : Span4Mux_v
    port map (
            O => \N__38781\,
            I => \N__38773\
        );

    \I__9536\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38770\
        );

    \I__9535\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38766\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__38776\,
            I => \N__38761\
        );

    \I__9533\ : Span4Mux_v
    port map (
            O => \N__38773\,
            I => \N__38755\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__38770\,
            I => \N__38755\
        );

    \I__9531\ : InMux
    port map (
            O => \N__38769\,
            I => \N__38751\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__38766\,
            I => \N__38748\
        );

    \I__9529\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38745\
        );

    \I__9528\ : InMux
    port map (
            O => \N__38764\,
            I => \N__38742\
        );

    \I__9527\ : Span4Mux_v
    port map (
            O => \N__38761\,
            I => \N__38739\
        );

    \I__9526\ : CascadeMux
    port map (
            O => \N__38760\,
            I => \N__38736\
        );

    \I__9525\ : Span4Mux_v
    port map (
            O => \N__38755\,
            I => \N__38733\
        );

    \I__9524\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38730\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__38751\,
            I => \N__38727\
        );

    \I__9522\ : Span4Mux_h
    port map (
            O => \N__38748\,
            I => \N__38722\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__38745\,
            I => \N__38722\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__38742\,
            I => \N__38719\
        );

    \I__9519\ : Span4Mux_h
    port map (
            O => \N__38739\,
            I => \N__38716\
        );

    \I__9518\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38713\
        );

    \I__9517\ : Span4Mux_h
    port map (
            O => \N__38733\,
            I => \N__38710\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__38730\,
            I => \N__38707\
        );

    \I__9515\ : Span12Mux_v
    port map (
            O => \N__38727\,
            I => \N__38704\
        );

    \I__9514\ : Span4Mux_v
    port map (
            O => \N__38722\,
            I => \N__38701\
        );

    \I__9513\ : Span12Mux_h
    port map (
            O => \N__38719\,
            I => \N__38698\
        );

    \I__9512\ : Span4Mux_h
    port map (
            O => \N__38716\,
            I => \N__38693\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__38713\,
            I => \N__38693\
        );

    \I__9510\ : Span4Mux_h
    port map (
            O => \N__38710\,
            I => \N__38688\
        );

    \I__9509\ : Span4Mux_v
    port map (
            O => \N__38707\,
            I => \N__38688\
        );

    \I__9508\ : Span12Mux_h
    port map (
            O => \N__38704\,
            I => \N__38685\
        );

    \I__9507\ : Span4Mux_h
    port map (
            O => \N__38701\,
            I => \N__38682\
        );

    \I__9506\ : Span12Mux_h
    port map (
            O => \N__38698\,
            I => \N__38677\
        );

    \I__9505\ : Sp12to4
    port map (
            O => \N__38693\,
            I => \N__38677\
        );

    \I__9504\ : IoSpan4Mux
    port map (
            O => \N__38688\,
            I => \N__38674\
        );

    \I__9503\ : Odrv12
    port map (
            O => \N__38685\,
            I => port_data_c_2
        );

    \I__9502\ : Odrv4
    port map (
            O => \N__38682\,
            I => port_data_c_2
        );

    \I__9501\ : Odrv12
    port map (
            O => \N__38677\,
            I => port_data_c_2
        );

    \I__9500\ : Odrv4
    port map (
            O => \N__38674\,
            I => port_data_c_2
        );

    \I__9499\ : IoInMux
    port map (
            O => \N__38665\,
            I => \N__38662\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__38662\,
            I => \N__38659\
        );

    \I__9497\ : IoSpan4Mux
    port map (
            O => \N__38659\,
            I => \N__38656\
        );

    \I__9496\ : Span4Mux_s2_v
    port map (
            O => \N__38656\,
            I => \N__38653\
        );

    \I__9495\ : Sp12to4
    port map (
            O => \N__38653\,
            I => \N__38649\
        );

    \I__9494\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38646\
        );

    \I__9493\ : Span12Mux_s10_v
    port map (
            O => \N__38649\,
            I => \N__38641\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__38646\,
            I => \N__38641\
        );

    \I__9491\ : Odrv12
    port map (
            O => \N__38641\,
            I => \M_this_ext_address_qZ0Z_10\
        );

    \I__9490\ : InMux
    port map (
            O => \N__38638\,
            I => \N__38635\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__38635\,
            I => \N__38632\
        );

    \I__9488\ : Span4Mux_v
    port map (
            O => \N__38632\,
            I => \N__38629\
        );

    \I__9487\ : Odrv4
    port map (
            O => \N__38629\,
            I => \un1_M_this_ext_address_q_cry_3_THRU_CO\
        );

    \I__9486\ : IoInMux
    port map (
            O => \N__38626\,
            I => \N__38622\
        );

    \I__9485\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38619\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__38622\,
            I => \N__38616\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__38619\,
            I => \N__38612\
        );

    \I__9482\ : Span12Mux_s6_h
    port map (
            O => \N__38616\,
            I => \N__38609\
        );

    \I__9481\ : InMux
    port map (
            O => \N__38615\,
            I => \N__38606\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__38612\,
            I => \N__38603\
        );

    \I__9479\ : Odrv12
    port map (
            O => \N__38609\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__38606\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__9477\ : Odrv4
    port map (
            O => \N__38603\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__9476\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38593\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__38593\,
            I => \N__38590\
        );

    \I__9474\ : Span4Mux_v
    port map (
            O => \N__38590\,
            I => \N__38587\
        );

    \I__9473\ : Span4Mux_h
    port map (
            O => \N__38587\,
            I => \N__38584\
        );

    \I__9472\ : Odrv4
    port map (
            O => \N__38584\,
            I => \this_ppu.un1_oam_data_1_4\
        );

    \I__9471\ : InMux
    port map (
            O => \N__38581\,
            I => \N__38578\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__38578\,
            I => \M_this_oam_ram_read_data_31\
        );

    \I__9469\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38572\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__38572\,
            I => \N__38569\
        );

    \I__9467\ : Odrv4
    port map (
            O => \N__38569\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_31\
        );

    \I__9466\ : InMux
    port map (
            O => \N__38566\,
            I => \N__38560\
        );

    \I__9465\ : InMux
    port map (
            O => \N__38565\,
            I => \N__38557\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__38564\,
            I => \N__38553\
        );

    \I__9463\ : CascadeMux
    port map (
            O => \N__38563\,
            I => \N__38550\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__38560\,
            I => \N__38547\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__38557\,
            I => \N__38544\
        );

    \I__9460\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38537\
        );

    \I__9459\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38537\
        );

    \I__9458\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38537\
        );

    \I__9457\ : Span4Mux_v
    port map (
            O => \N__38547\,
            I => \N__38534\
        );

    \I__9456\ : Span4Mux_h
    port map (
            O => \N__38544\,
            I => \N__38529\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__38537\,
            I => \N__38529\
        );

    \I__9454\ : Span4Mux_v
    port map (
            O => \N__38534\,
            I => \N__38526\
        );

    \I__9453\ : Odrv4
    port map (
            O => \N__38529\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__9452\ : Odrv4
    port map (
            O => \N__38526\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__9451\ : InMux
    port map (
            O => \N__38521\,
            I => \N__38518\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__38518\,
            I => \N__38515\
        );

    \I__9449\ : Odrv4
    port map (
            O => \N__38515\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_19\
        );

    \I__9448\ : CascadeMux
    port map (
            O => \N__38512\,
            I => \N__38509\
        );

    \I__9447\ : InMux
    port map (
            O => \N__38509\,
            I => \N__38505\
        );

    \I__9446\ : InMux
    port map (
            O => \N__38508\,
            I => \N__38502\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__38505\,
            I => \N__38497\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__38502\,
            I => \N__38494\
        );

    \I__9443\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38489\
        );

    \I__9442\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38489\
        );

    \I__9441\ : Span4Mux_h
    port map (
            O => \N__38497\,
            I => \N__38486\
        );

    \I__9440\ : Span4Mux_h
    port map (
            O => \N__38494\,
            I => \N__38481\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__38489\,
            I => \N__38481\
        );

    \I__9438\ : Span4Mux_v
    port map (
            O => \N__38486\,
            I => \N__38478\
        );

    \I__9437\ : Odrv4
    port map (
            O => \N__38481\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__9436\ : Odrv4
    port map (
            O => \N__38478\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__9435\ : InMux
    port map (
            O => \N__38473\,
            I => \N__38470\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__38470\,
            I => \N__38467\
        );

    \I__9433\ : Span4Mux_h
    port map (
            O => \N__38467\,
            I => \N__38464\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__38464\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_20\
        );

    \I__9431\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38458\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__38458\,
            I => \M_this_oam_ram_read_data_24\
        );

    \I__9429\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38452\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__38452\,
            I => \N__38449\
        );

    \I__9427\ : Span4Mux_h
    port map (
            O => \N__38449\,
            I => \N__38446\
        );

    \I__9426\ : Odrv4
    port map (
            O => \N__38446\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_24\
        );

    \I__9425\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38438\
        );

    \I__9424\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38435\
        );

    \I__9423\ : InMux
    port map (
            O => \N__38441\,
            I => \N__38432\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__38438\,
            I => \N__38427\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__38435\,
            I => \N__38424\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__38432\,
            I => \N__38421\
        );

    \I__9419\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38416\
        );

    \I__9418\ : InMux
    port map (
            O => \N__38430\,
            I => \N__38416\
        );

    \I__9417\ : Span4Mux_v
    port map (
            O => \N__38427\,
            I => \N__38412\
        );

    \I__9416\ : Span12Mux_v
    port map (
            O => \N__38424\,
            I => \N__38409\
        );

    \I__9415\ : Span4Mux_h
    port map (
            O => \N__38421\,
            I => \N__38404\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38404\
        );

    \I__9413\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38401\
        );

    \I__9412\ : Span4Mux_v
    port map (
            O => \N__38412\,
            I => \N__38398\
        );

    \I__9411\ : Odrv12
    port map (
            O => \N__38409\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__38404\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__38401\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__9408\ : Odrv4
    port map (
            O => \N__38398\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__9407\ : InMux
    port map (
            O => \N__38389\,
            I => \N__38386\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__38386\,
            I => \N__38383\
        );

    \I__9405\ : Span4Mux_h
    port map (
            O => \N__38383\,
            I => \N__38380\
        );

    \I__9404\ : Span4Mux_v
    port map (
            O => \N__38380\,
            I => \N__38377\
        );

    \I__9403\ : Odrv4
    port map (
            O => \N__38377\,
            I => \this_ppu.un1_oam_data_1_2\
        );

    \I__9402\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38371\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38368\
        );

    \I__9400\ : Odrv12
    port map (
            O => \N__38368\,
            I => \M_this_data_tmp_qZ0Z_17\
        );

    \I__9399\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38362\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__38362\,
            I => \M_this_oam_ram_write_data_17\
        );

    \I__9397\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38356\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__38356\,
            I => \N__38352\
        );

    \I__9395\ : InMux
    port map (
            O => \N__38355\,
            I => \N__38349\
        );

    \I__9394\ : Span4Mux_v
    port map (
            O => \N__38352\,
            I => \N__38346\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__38349\,
            I => \this_ppu.un1_oam_data_1_4_c2\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__38346\,
            I => \this_ppu.un1_oam_data_1_4_c2\
        );

    \I__9391\ : InMux
    port map (
            O => \N__38341\,
            I => \N__38335\
        );

    \I__9390\ : InMux
    port map (
            O => \N__38340\,
            I => \N__38335\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__38335\,
            I => \M_this_oam_ram_read_data_5\
        );

    \I__9388\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38329\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__38329\,
            I => \N__38326\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__38326\,
            I => \N__38323\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__38323\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_5\
        );

    \I__9384\ : InMux
    port map (
            O => \N__38320\,
            I => \N__38314\
        );

    \I__9383\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38314\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__38314\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__9381\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38308\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__38308\,
            I => \N__38305\
        );

    \I__9379\ : Odrv4
    port map (
            O => \N__38305\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_6\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__38302\,
            I => \N__38298\
        );

    \I__9377\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38293\
        );

    \I__9376\ : InMux
    port map (
            O => \N__38298\,
            I => \N__38293\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__38293\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__9374\ : InMux
    port map (
            O => \N__38290\,
            I => \N__38287\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__38287\,
            I => \N__38284\
        );

    \I__9372\ : Odrv4
    port map (
            O => \N__38284\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_7\
        );

    \I__9371\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38278\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__38278\,
            I => \N__38275\
        );

    \I__9369\ : Odrv4
    port map (
            O => \N__38275\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_0\
        );

    \I__9368\ : InMux
    port map (
            O => \N__38272\,
            I => \N__38269\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__38269\,
            I => \N__38266\
        );

    \I__9366\ : Span4Mux_h
    port map (
            O => \N__38266\,
            I => \N__38263\
        );

    \I__9365\ : Odrv4
    port map (
            O => \N__38263\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_1\
        );

    \I__9364\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38257\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__38257\,
            I => \N__38253\
        );

    \I__9362\ : InMux
    port map (
            O => \N__38256\,
            I => \N__38250\
        );

    \I__9361\ : Odrv4
    port map (
            O => \N__38253\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__38250\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__9359\ : InMux
    port map (
            O => \N__38245\,
            I => \N__38239\
        );

    \I__9358\ : InMux
    port map (
            O => \N__38244\,
            I => \N__38239\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__38239\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__9356\ : InMux
    port map (
            O => \N__38236\,
            I => \N__38232\
        );

    \I__9355\ : CascadeMux
    port map (
            O => \N__38235\,
            I => \N__38229\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__38232\,
            I => \N__38226\
        );

    \I__9353\ : InMux
    port map (
            O => \N__38229\,
            I => \N__38223\
        );

    \I__9352\ : Odrv4
    port map (
            O => \N__38226\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__38223\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__9350\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38212\
        );

    \I__9349\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38212\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__38212\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__9347\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38206\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__38206\,
            I => \N__38203\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__38203\,
            I => \this_ppu.un12lto7Z0Z_5\
        );

    \I__9344\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38197\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__38197\,
            I => \M_this_oam_ram_read_data_27\
        );

    \I__9342\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38191\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__38191\,
            I => \N__38188\
        );

    \I__9340\ : Span4Mux_h
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__9339\ : Odrv4
    port map (
            O => \N__38185\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_27\
        );

    \I__9338\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38179\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__38179\,
            I => \N__38176\
        );

    \I__9336\ : Span4Mux_h
    port map (
            O => \N__38176\,
            I => \N__38173\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__38173\,
            I => \N__38170\
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__38170\,
            I => \this_ppu.un1_oam_data_1_3\
        );

    \I__9333\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38164\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__38164\,
            I => \M_this_oam_ram_read_data_29\
        );

    \I__9331\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38158\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__38158\,
            I => \N__38155\
        );

    \I__9329\ : Span4Mux_h
    port map (
            O => \N__38155\,
            I => \N__38152\
        );

    \I__9328\ : Odrv4
    port map (
            O => \N__38152\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_29\
        );

    \I__9327\ : InMux
    port map (
            O => \N__38149\,
            I => \N__38146\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__38146\,
            I => \N__38143\
        );

    \I__9325\ : Span4Mux_h
    port map (
            O => \N__38143\,
            I => \N__38140\
        );

    \I__9324\ : Odrv4
    port map (
            O => \N__38140\,
            I => \M_this_oam_ram_read_data_25\
        );

    \I__9323\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38134\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__38134\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_25\
        );

    \I__9321\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38128\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__38128\,
            I => \N__38125\
        );

    \I__9319\ : Span4Mux_v
    port map (
            O => \N__38125\,
            I => \N__38122\
        );

    \I__9318\ : Odrv4
    port map (
            O => \N__38122\,
            I => \M_this_oam_ram_read_data_26\
        );

    \I__9317\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__38116\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_26\
        );

    \I__9315\ : InMux
    port map (
            O => \N__38113\,
            I => \N__38110\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__38110\,
            I => \N__38107\
        );

    \I__9313\ : Span12Mux_s9_h
    port map (
            O => \N__38107\,
            I => \N__38104\
        );

    \I__9312\ : Odrv12
    port map (
            O => \N__38104\,
            I => \M_this_data_tmp_qZ0Z_10\
        );

    \I__9311\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38098\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__38098\,
            I => \M_this_oam_ram_write_data_10\
        );

    \I__9309\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38092\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__38092\,
            I => \M_this_data_tmp_qZ0Z_6\
        );

    \I__9307\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38086\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__38086\,
            I => \N__38083\
        );

    \I__9305\ : Odrv4
    port map (
            O => \N__38083\,
            I => \M_this_oam_ram_write_data_6\
        );

    \I__9304\ : InMux
    port map (
            O => \N__38080\,
            I => \N__38077\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__38077\,
            I => \N__38074\
        );

    \I__9302\ : Span4Mux_h
    port map (
            O => \N__38074\,
            I => \N__38071\
        );

    \I__9301\ : Span4Mux_h
    port map (
            O => \N__38071\,
            I => \N__38068\
        );

    \I__9300\ : Odrv4
    port map (
            O => \N__38068\,
            I => \M_this_data_tmp_qZ0Z_11\
        );

    \I__9299\ : InMux
    port map (
            O => \N__38065\,
            I => \N__38062\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__38062\,
            I => \N__38059\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__38059\,
            I => \M_this_oam_ram_write_data_11\
        );

    \I__9296\ : InMux
    port map (
            O => \N__38056\,
            I => \N__38053\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__38053\,
            I => \N__38050\
        );

    \I__9294\ : Span4Mux_h
    port map (
            O => \N__38050\,
            I => \N__38047\
        );

    \I__9293\ : Odrv4
    port map (
            O => \N__38047\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_2\
        );

    \I__9292\ : InMux
    port map (
            O => \N__38044\,
            I => \N__38041\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__38041\,
            I => \N__38038\
        );

    \I__9290\ : Odrv4
    port map (
            O => \N__38038\,
            I => \this_ppu.un12lto7Z0Z_4\
        );

    \I__9289\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38029\
        );

    \I__9288\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38029\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__38029\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__9286\ : InMux
    port map (
            O => \N__38026\,
            I => \N__38023\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__38023\,
            I => \N__38020\
        );

    \I__9284\ : Span4Mux_h
    port map (
            O => \N__38020\,
            I => \N__38017\
        );

    \I__9283\ : Odrv4
    port map (
            O => \N__38017\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_4\
        );

    \I__9282\ : InMux
    port map (
            O => \N__38014\,
            I => \un1_M_this_ext_address_q_cry_12\
        );

    \I__9281\ : IoInMux
    port map (
            O => \N__38011\,
            I => \N__38008\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__38008\,
            I => \N__38005\
        );

    \I__9279\ : Span4Mux_s1_h
    port map (
            O => \N__38005\,
            I => \N__38002\
        );

    \I__9278\ : Sp12to4
    port map (
            O => \N__38002\,
            I => \N__37998\
        );

    \I__9277\ : CascadeMux
    port map (
            O => \N__38001\,
            I => \N__37995\
        );

    \I__9276\ : Span12Mux_v
    port map (
            O => \N__37998\,
            I => \N__37992\
        );

    \I__9275\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37989\
        );

    \I__9274\ : Odrv12
    port map (
            O => \N__37992\,
            I => \M_this_ext_address_qZ0Z_14\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__37989\,
            I => \M_this_ext_address_qZ0Z_14\
        );

    \I__9272\ : InMux
    port map (
            O => \N__37984\,
            I => \N__37981\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__37981\,
            I => \un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0\
        );

    \I__9270\ : InMux
    port map (
            O => \N__37978\,
            I => \un1_M_this_ext_address_q_cry_13\
        );

    \I__9269\ : IoInMux
    port map (
            O => \N__37975\,
            I => \N__37972\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__37972\,
            I => \N__37969\
        );

    \I__9267\ : Span4Mux_s0_h
    port map (
            O => \N__37969\,
            I => \N__37966\
        );

    \I__9266\ : Sp12to4
    port map (
            O => \N__37966\,
            I => \N__37962\
        );

    \I__9265\ : InMux
    port map (
            O => \N__37965\,
            I => \N__37959\
        );

    \I__9264\ : Span12Mux_v
    port map (
            O => \N__37962\,
            I => \N__37956\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__37959\,
            I => \N__37953\
        );

    \I__9262\ : Odrv12
    port map (
            O => \N__37956\,
            I => \M_this_ext_address_qZ0Z_15\
        );

    \I__9261\ : Odrv4
    port map (
            O => \N__37953\,
            I => \M_this_ext_address_qZ0Z_15\
        );

    \I__9260\ : InMux
    port map (
            O => \N__37948\,
            I => \un1_M_this_ext_address_q_cry_14\
        );

    \I__9259\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37942\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__37942\,
            I => \N__37939\
        );

    \I__9257\ : Odrv4
    port map (
            O => \N__37939\,
            I => \un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0\
        );

    \I__9256\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37933\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__37933\,
            I => \N__37930\
        );

    \I__9254\ : Odrv4
    port map (
            O => \N__37930\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__9253\ : InMux
    port map (
            O => \N__37927\,
            I => \N__37924\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__37924\,
            I => \N__37921\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__37921\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_13\
        );

    \I__9250\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37915\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__37915\,
            I => \N__37912\
        );

    \I__9248\ : Odrv4
    port map (
            O => \N__37912\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__9247\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37906\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__37906\,
            I => \N__37903\
        );

    \I__9245\ : Odrv4
    port map (
            O => \N__37903\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_15\
        );

    \I__9244\ : InMux
    port map (
            O => \N__37900\,
            I => \N__37897\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__37897\,
            I => \N__37894\
        );

    \I__9242\ : Odrv4
    port map (
            O => \N__37894\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_3\
        );

    \I__9241\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37888\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__37888\,
            I => \N__37885\
        );

    \I__9239\ : Odrv4
    port map (
            O => \N__37885\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__9238\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37879\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__37879\,
            I => \N__37876\
        );

    \I__9236\ : Odrv4
    port map (
            O => \N__37876\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_8\
        );

    \I__9235\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37870\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__37870\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_16\
        );

    \I__9233\ : InMux
    port map (
            O => \N__37867\,
            I => \N__37864\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__37864\,
            I => \N__37861\
        );

    \I__9231\ : Odrv4
    port map (
            O => \N__37861\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__9230\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37855\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__37855\,
            I => \N__37852\
        );

    \I__9228\ : Odrv4
    port map (
            O => \N__37852\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_10\
        );

    \I__9227\ : InMux
    port map (
            O => \N__37849\,
            I => \un1_M_this_ext_address_q_cry_3\
        );

    \I__9226\ : InMux
    port map (
            O => \N__37846\,
            I => \un1_M_this_ext_address_q_cry_4\
        );

    \I__9225\ : InMux
    port map (
            O => \N__37843\,
            I => \un1_M_this_ext_address_q_cry_5\
        );

    \I__9224\ : InMux
    port map (
            O => \N__37840\,
            I => \un1_M_this_ext_address_q_cry_6\
        );

    \I__9223\ : IoInMux
    port map (
            O => \N__37837\,
            I => \N__37834\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__37834\,
            I => \N__37831\
        );

    \I__9221\ : IoSpan4Mux
    port map (
            O => \N__37831\,
            I => \N__37828\
        );

    \I__9220\ : IoSpan4Mux
    port map (
            O => \N__37828\,
            I => \N__37825\
        );

    \I__9219\ : Span4Mux_s2_v
    port map (
            O => \N__37825\,
            I => \N__37822\
        );

    \I__9218\ : Sp12to4
    port map (
            O => \N__37822\,
            I => \N__37818\
        );

    \I__9217\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37815\
        );

    \I__9216\ : Odrv12
    port map (
            O => \N__37818\,
            I => \M_this_ext_address_qZ0Z_8\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__37815\,
            I => \M_this_ext_address_qZ0Z_8\
        );

    \I__9214\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37807\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__37807\,
            I => \un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0\
        );

    \I__9212\ : InMux
    port map (
            O => \N__37804\,
            I => \bfn_24_22_0_\
        );

    \I__9211\ : IoInMux
    port map (
            O => \N__37801\,
            I => \N__37798\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__37798\,
            I => \N__37795\
        );

    \I__9209\ : IoSpan4Mux
    port map (
            O => \N__37795\,
            I => \N__37792\
        );

    \I__9208\ : Span4Mux_s3_v
    port map (
            O => \N__37792\,
            I => \N__37789\
        );

    \I__9207\ : Span4Mux_v
    port map (
            O => \N__37789\,
            I => \N__37785\
        );

    \I__9206\ : InMux
    port map (
            O => \N__37788\,
            I => \N__37782\
        );

    \I__9205\ : Odrv4
    port map (
            O => \N__37785\,
            I => \M_this_ext_address_qZ0Z_9\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__37782\,
            I => \M_this_ext_address_qZ0Z_9\
        );

    \I__9203\ : CascadeMux
    port map (
            O => \N__37777\,
            I => \N__37774\
        );

    \I__9202\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37771\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__37771\,
            I => \N__37768\
        );

    \I__9200\ : Odrv4
    port map (
            O => \N__37768\,
            I => \un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0\
        );

    \I__9199\ : InMux
    port map (
            O => \N__37765\,
            I => \un1_M_this_ext_address_q_cry_8\
        );

    \I__9198\ : InMux
    port map (
            O => \N__37762\,
            I => \un1_M_this_ext_address_q_cry_9\
        );

    \I__9197\ : InMux
    port map (
            O => \N__37759\,
            I => \un1_M_this_ext_address_q_cry_10\
        );

    \I__9196\ : InMux
    port map (
            O => \N__37756\,
            I => \un1_M_this_ext_address_q_cry_11\
        );

    \I__9195\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37750\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37747\
        );

    \I__9193\ : Span12Mux_v
    port map (
            O => \N__37747\,
            I => \N__37744\
        );

    \I__9192\ : Span12Mux_h
    port map (
            O => \N__37744\,
            I => \N__37740\
        );

    \I__9191\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37737\
        );

    \I__9190\ : Odrv12
    port map (
            O => \N__37740\,
            I => \M_this_ctrl_flags_qZ0Z_7\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__37737\,
            I => \M_this_ctrl_flags_qZ0Z_7\
        );

    \I__9188\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37728\
        );

    \I__9187\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37725\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37722\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__37725\,
            I => \N_312_0\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__37722\,
            I => \N_312_0\
        );

    \I__9183\ : IoInMux
    port map (
            O => \N__37717\,
            I => \N__37714\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__37714\,
            I => \N__37711\
        );

    \I__9181\ : Span4Mux_s0_v
    port map (
            O => \N__37711\,
            I => \N__37708\
        );

    \I__9180\ : Sp12to4
    port map (
            O => \N__37708\,
            I => \N__37705\
        );

    \I__9179\ : Span12Mux_h
    port map (
            O => \N__37705\,
            I => \N__37701\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__37704\,
            I => \N__37697\
        );

    \I__9177\ : Span12Mux_v
    port map (
            O => \N__37701\,
            I => \N__37694\
        );

    \I__9176\ : InMux
    port map (
            O => \N__37700\,
            I => \N__37691\
        );

    \I__9175\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37688\
        );

    \I__9174\ : Odrv12
    port map (
            O => \N__37694\,
            I => \M_this_ext_address_qZ0Z_0\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__37691\,
            I => \M_this_ext_address_qZ0Z_0\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__37688\,
            I => \M_this_ext_address_qZ0Z_0\
        );

    \I__9171\ : IoInMux
    port map (
            O => \N__37681\,
            I => \N__37678\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__37678\,
            I => \N__37675\
        );

    \I__9169\ : IoSpan4Mux
    port map (
            O => \N__37675\,
            I => \N__37672\
        );

    \I__9168\ : Sp12to4
    port map (
            O => \N__37672\,
            I => \N__37669\
        );

    \I__9167\ : Span12Mux_v
    port map (
            O => \N__37669\,
            I => \N__37664\
        );

    \I__9166\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37661\
        );

    \I__9165\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37658\
        );

    \I__9164\ : Odrv12
    port map (
            O => \N__37664\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__37661\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__37658\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__9161\ : CascadeMux
    port map (
            O => \N__37651\,
            I => \N__37648\
        );

    \I__9160\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37645\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__37645\,
            I => \N__37642\
        );

    \I__9158\ : Odrv4
    port map (
            O => \N__37642\,
            I => \un1_M_this_ext_address_q_cry_0_THRU_CO\
        );

    \I__9157\ : InMux
    port map (
            O => \N__37639\,
            I => \un1_M_this_ext_address_q_cry_0\
        );

    \I__9156\ : IoInMux
    port map (
            O => \N__37636\,
            I => \N__37633\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__37633\,
            I => \N__37630\
        );

    \I__9154\ : Span12Mux_s0_v
    port map (
            O => \N__37630\,
            I => \N__37627\
        );

    \I__9153\ : Span12Mux_v
    port map (
            O => \N__37627\,
            I => \N__37622\
        );

    \I__9152\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37619\
        );

    \I__9151\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37616\
        );

    \I__9150\ : Odrv12
    port map (
            O => \N__37622\,
            I => \M_this_ext_address_qZ0Z_2\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__37619\,
            I => \M_this_ext_address_qZ0Z_2\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__37616\,
            I => \M_this_ext_address_qZ0Z_2\
        );

    \I__9147\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37606\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__37606\,
            I => \un1_M_this_ext_address_q_cry_1_THRU_CO\
        );

    \I__9145\ : InMux
    port map (
            O => \N__37603\,
            I => \un1_M_this_ext_address_q_cry_1\
        );

    \I__9144\ : IoInMux
    port map (
            O => \N__37600\,
            I => \N__37597\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__37597\,
            I => \N__37594\
        );

    \I__9142\ : Span4Mux_s1_h
    port map (
            O => \N__37594\,
            I => \N__37591\
        );

    \I__9141\ : Span4Mux_h
    port map (
            O => \N__37591\,
            I => \N__37588\
        );

    \I__9140\ : Span4Mux_v
    port map (
            O => \N__37588\,
            I => \N__37585\
        );

    \I__9139\ : Span4Mux_v
    port map (
            O => \N__37585\,
            I => \N__37580\
        );

    \I__9138\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37577\
        );

    \I__9137\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37574\
        );

    \I__9136\ : Odrv4
    port map (
            O => \N__37580\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__37577\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__37574\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__9133\ : CascadeMux
    port map (
            O => \N__37567\,
            I => \N__37564\
        );

    \I__9132\ : InMux
    port map (
            O => \N__37564\,
            I => \N__37561\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__37561\,
            I => \un1_M_this_ext_address_q_cry_2_THRU_CO\
        );

    \I__9130\ : InMux
    port map (
            O => \N__37558\,
            I => \un1_M_this_ext_address_q_cry_2\
        );

    \I__9129\ : InMux
    port map (
            O => \N__37555\,
            I => \N__37552\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__37552\,
            I => \N__37544\
        );

    \I__9127\ : InMux
    port map (
            O => \N__37551\,
            I => \N__37541\
        );

    \I__9126\ : InMux
    port map (
            O => \N__37550\,
            I => \N__37538\
        );

    \I__9125\ : InMux
    port map (
            O => \N__37549\,
            I => \N__37535\
        );

    \I__9124\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37530\
        );

    \I__9123\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37530\
        );

    \I__9122\ : Span4Mux_v
    port map (
            O => \N__37544\,
            I => \N__37522\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37522\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__37538\,
            I => \N__37522\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__37535\,
            I => \N__37519\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__37530\,
            I => \N__37516\
        );

    \I__9117\ : InMux
    port map (
            O => \N__37529\,
            I => \N__37513\
        );

    \I__9116\ : Span4Mux_h
    port map (
            O => \N__37522\,
            I => \N__37510\
        );

    \I__9115\ : Span4Mux_h
    port map (
            O => \N__37519\,
            I => \N__37507\
        );

    \I__9114\ : Span4Mux_h
    port map (
            O => \N__37516\,
            I => \N__37504\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__37513\,
            I => \N__37501\
        );

    \I__9112\ : Span4Mux_v
    port map (
            O => \N__37510\,
            I => \N__37497\
        );

    \I__9111\ : Span4Mux_v
    port map (
            O => \N__37507\,
            I => \N__37492\
        );

    \I__9110\ : Span4Mux_h
    port map (
            O => \N__37504\,
            I => \N__37492\
        );

    \I__9109\ : Span4Mux_h
    port map (
            O => \N__37501\,
            I => \N__37489\
        );

    \I__9108\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37486\
        );

    \I__9107\ : Odrv4
    port map (
            O => \N__37497\,
            I => \N_260_0\
        );

    \I__9106\ : Odrv4
    port map (
            O => \N__37492\,
            I => \N_260_0\
        );

    \I__9105\ : Odrv4
    port map (
            O => \N__37489\,
            I => \N_260_0\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__37486\,
            I => \N_260_0\
        );

    \I__9103\ : CascadeMux
    port map (
            O => \N__37477\,
            I => \N__37471\
        );

    \I__9102\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37468\
        );

    \I__9101\ : CascadeMux
    port map (
            O => \N__37475\,
            I => \N__37463\
        );

    \I__9100\ : CascadeMux
    port map (
            O => \N__37474\,
            I => \N__37459\
        );

    \I__9099\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37456\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__37468\,
            I => \N__37453\
        );

    \I__9097\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37450\
        );

    \I__9096\ : InMux
    port map (
            O => \N__37466\,
            I => \N__37445\
        );

    \I__9095\ : InMux
    port map (
            O => \N__37463\,
            I => \N__37445\
        );

    \I__9094\ : CascadeMux
    port map (
            O => \N__37462\,
            I => \N__37442\
        );

    \I__9093\ : InMux
    port map (
            O => \N__37459\,
            I => \N__37438\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__37456\,
            I => \N__37435\
        );

    \I__9091\ : Span4Mux_v
    port map (
            O => \N__37453\,
            I => \N__37428\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__37450\,
            I => \N__37428\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__37445\,
            I => \N__37428\
        );

    \I__9088\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37425\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__37441\,
            I => \N__37422\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__37438\,
            I => \N__37418\
        );

    \I__9085\ : Span4Mux_v
    port map (
            O => \N__37435\,
            I => \N__37415\
        );

    \I__9084\ : Span4Mux_v
    port map (
            O => \N__37428\,
            I => \N__37412\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__37425\,
            I => \N__37409\
        );

    \I__9082\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37406\
        );

    \I__9081\ : InMux
    port map (
            O => \N__37421\,
            I => \N__37403\
        );

    \I__9080\ : Span4Mux_v
    port map (
            O => \N__37418\,
            I => \N__37400\
        );

    \I__9079\ : Span4Mux_v
    port map (
            O => \N__37415\,
            I => \N__37391\
        );

    \I__9078\ : Span4Mux_h
    port map (
            O => \N__37412\,
            I => \N__37391\
        );

    \I__9077\ : Span4Mux_v
    port map (
            O => \N__37409\,
            I => \N__37391\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__37406\,
            I => \N__37391\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__37403\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__37400\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__9073\ : Odrv4
    port map (
            O => \N__37391\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__9072\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37380\
        );

    \I__9071\ : CascadeMux
    port map (
            O => \N__37383\,
            I => \N__37376\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__37380\,
            I => \N__37370\
        );

    \I__9069\ : InMux
    port map (
            O => \N__37379\,
            I => \N__37367\
        );

    \I__9068\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37362\
        );

    \I__9067\ : InMux
    port map (
            O => \N__37375\,
            I => \N__37362\
        );

    \I__9066\ : InMux
    port map (
            O => \N__37374\,
            I => \N__37359\
        );

    \I__9065\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37355\
        );

    \I__9064\ : Span4Mux_v
    port map (
            O => \N__37370\,
            I => \N__37348\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__37367\,
            I => \N__37348\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__37362\,
            I => \N__37348\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__37359\,
            I => \N__37345\
        );

    \I__9060\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37342\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37337\
        );

    \I__9058\ : Span4Mux_v
    port map (
            O => \N__37348\,
            I => \N__37334\
        );

    \I__9057\ : Span4Mux_v
    port map (
            O => \N__37345\,
            I => \N__37329\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__37342\,
            I => \N__37329\
        );

    \I__9055\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37326\
        );

    \I__9054\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37323\
        );

    \I__9053\ : Span4Mux_v
    port map (
            O => \N__37337\,
            I => \N__37320\
        );

    \I__9052\ : Span4Mux_h
    port map (
            O => \N__37334\,
            I => \N__37313\
        );

    \I__9051\ : Span4Mux_v
    port map (
            O => \N__37329\,
            I => \N__37313\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__37326\,
            I => \N__37313\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__37323\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__9048\ : Odrv4
    port map (
            O => \N__37320\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__9047\ : Odrv4
    port map (
            O => \N__37313\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__9046\ : CascadeMux
    port map (
            O => \N__37306\,
            I => \N__37297\
        );

    \I__9045\ : CascadeMux
    port map (
            O => \N__37305\,
            I => \N__37294\
        );

    \I__9044\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37291\
        );

    \I__9043\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37288\
        );

    \I__9042\ : InMux
    port map (
            O => \N__37302\,
            I => \N__37283\
        );

    \I__9041\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37283\
        );

    \I__9040\ : InMux
    port map (
            O => \N__37300\,
            I => \N__37280\
        );

    \I__9039\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37277\
        );

    \I__9038\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37274\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__37291\,
            I => \N__37270\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__37288\,
            I => \N__37267\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__37283\,
            I => \N__37264\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__37280\,
            I => \N__37261\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__37277\,
            I => \N__37255\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__37274\,
            I => \N__37255\
        );

    \I__9031\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37252\
        );

    \I__9030\ : Span4Mux_v
    port map (
            O => \N__37270\,
            I => \N__37249\
        );

    \I__9029\ : Span4Mux_v
    port map (
            O => \N__37267\,
            I => \N__37244\
        );

    \I__9028\ : Span4Mux_h
    port map (
            O => \N__37264\,
            I => \N__37244\
        );

    \I__9027\ : Span4Mux_h
    port map (
            O => \N__37261\,
            I => \N__37241\
        );

    \I__9026\ : InMux
    port map (
            O => \N__37260\,
            I => \N__37238\
        );

    \I__9025\ : Span12Mux_v
    port map (
            O => \N__37255\,
            I => \N__37233\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__37252\,
            I => \N__37233\
        );

    \I__9023\ : Span4Mux_h
    port map (
            O => \N__37249\,
            I => \N__37230\
        );

    \I__9022\ : Span4Mux_h
    port map (
            O => \N__37244\,
            I => \N__37225\
        );

    \I__9021\ : Span4Mux_v
    port map (
            O => \N__37241\,
            I => \N__37225\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__37238\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__9019\ : Odrv12
    port map (
            O => \N__37233\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__37230\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__37225\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__9016\ : CEMux
    port map (
            O => \N__37216\,
            I => \N__37213\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__37213\,
            I => \N__37209\
        );

    \I__9014\ : CEMux
    port map (
            O => \N__37212\,
            I => \N__37206\
        );

    \I__9013\ : Odrv4
    port map (
            O => \N__37209\,
            I => \this_spr_ram.mem_WE_12\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__37206\,
            I => \this_spr_ram.mem_WE_12\
        );

    \I__9011\ : InMux
    port map (
            O => \N__37201\,
            I => \N__37198\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__37198\,
            I => \N__37195\
        );

    \I__9009\ : Span4Mux_v
    port map (
            O => \N__37195\,
            I => \N__37190\
        );

    \I__9008\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37187\
        );

    \I__9007\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37184\
        );

    \I__9006\ : Sp12to4
    port map (
            O => \N__37190\,
            I => \N__37178\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__37187\,
            I => \N__37178\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__37184\,
            I => \N__37175\
        );

    \I__9003\ : InMux
    port map (
            O => \N__37183\,
            I => \N__37172\
        );

    \I__9002\ : Odrv12
    port map (
            O => \N__37178\,
            I => \this_ppu.N_545\
        );

    \I__9001\ : Odrv4
    port map (
            O => \N__37175\,
            I => \this_ppu.N_545\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__37172\,
            I => \this_ppu.N_545\
        );

    \I__8999\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37162\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__37162\,
            I => \N__37158\
        );

    \I__8997\ : InMux
    port map (
            O => \N__37161\,
            I => \N__37155\
        );

    \I__8996\ : Span4Mux_h
    port map (
            O => \N__37158\,
            I => \N__37150\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__37155\,
            I => \N__37147\
        );

    \I__8994\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37144\
        );

    \I__8993\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37141\
        );

    \I__8992\ : Span4Mux_v
    port map (
            O => \N__37150\,
            I => \N__37135\
        );

    \I__8991\ : Span4Mux_h
    port map (
            O => \N__37147\,
            I => \N__37135\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__37144\,
            I => \N__37132\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__37141\,
            I => \N__37129\
        );

    \I__8988\ : InMux
    port map (
            O => \N__37140\,
            I => \N__37126\
        );

    \I__8987\ : Span4Mux_v
    port map (
            O => \N__37135\,
            I => \N__37120\
        );

    \I__8986\ : Span4Mux_h
    port map (
            O => \N__37132\,
            I => \N__37120\
        );

    \I__8985\ : Span4Mux_s2_v
    port map (
            O => \N__37129\,
            I => \N__37115\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__37126\,
            I => \N__37115\
        );

    \I__8983\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37112\
        );

    \I__8982\ : Sp12to4
    port map (
            O => \N__37120\,
            I => \N__37108\
        );

    \I__8981\ : Span4Mux_v
    port map (
            O => \N__37115\,
            I => \N__37103\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__37112\,
            I => \N__37103\
        );

    \I__8979\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37100\
        );

    \I__8978\ : Span12Mux_h
    port map (
            O => \N__37108\,
            I => \N__37096\
        );

    \I__8977\ : Span4Mux_v
    port map (
            O => \N__37103\,
            I => \N__37093\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37090\
        );

    \I__8975\ : InMux
    port map (
            O => \N__37099\,
            I => \N__37087\
        );

    \I__8974\ : Odrv12
    port map (
            O => \N__37096\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__8973\ : Odrv4
    port map (
            O => \N__37093\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__8972\ : Odrv4
    port map (
            O => \N__37090\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__37087\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__8970\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37071\
        );

    \I__8969\ : CascadeMux
    port map (
            O => \N__37077\,
            I => \N__37068\
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__37076\,
            I => \N__37065\
        );

    \I__8967\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37058\
        );

    \I__8966\ : InMux
    port map (
            O => \N__37074\,
            I => \N__37058\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__37071\,
            I => \N__37055\
        );

    \I__8964\ : InMux
    port map (
            O => \N__37068\,
            I => \N__37052\
        );

    \I__8963\ : InMux
    port map (
            O => \N__37065\,
            I => \N__37049\
        );

    \I__8962\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37046\
        );

    \I__8961\ : InMux
    port map (
            O => \N__37063\,
            I => \N__37043\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__37058\,
            I => \N__37040\
        );

    \I__8959\ : Span4Mux_v
    port map (
            O => \N__37055\,
            I => \N__37033\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__37052\,
            I => \N__37033\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__37049\,
            I => \N__37033\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__37046\,
            I => \N__37030\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__37043\,
            I => \N__37027\
        );

    \I__8954\ : Span4Mux_v
    port map (
            O => \N__37040\,
            I => \N__37024\
        );

    \I__8953\ : Span4Mux_h
    port map (
            O => \N__37033\,
            I => \N__37021\
        );

    \I__8952\ : Span4Mux_v
    port map (
            O => \N__37030\,
            I => \N__37018\
        );

    \I__8951\ : Span4Mux_v
    port map (
            O => \N__37027\,
            I => \N__37015\
        );

    \I__8950\ : Span4Mux_v
    port map (
            O => \N__37024\,
            I => \N__37012\
        );

    \I__8949\ : Sp12to4
    port map (
            O => \N__37021\,
            I => \N__37009\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__37018\,
            I => \N__37004\
        );

    \I__8947\ : Span4Mux_v
    port map (
            O => \N__37015\,
            I => \N__37004\
        );

    \I__8946\ : Sp12to4
    port map (
            O => \N__37012\,
            I => \N__37001\
        );

    \I__8945\ : Span12Mux_v
    port map (
            O => \N__37009\,
            I => \N__36998\
        );

    \I__8944\ : Span4Mux_h
    port map (
            O => \N__37004\,
            I => \N__36995\
        );

    \I__8943\ : Odrv12
    port map (
            O => \N__37001\,
            I => port_address_in_4
        );

    \I__8942\ : Odrv12
    port map (
            O => \N__36998\,
            I => port_address_in_4
        );

    \I__8941\ : Odrv4
    port map (
            O => \N__36995\,
            I => port_address_in_4
        );

    \I__8940\ : InMux
    port map (
            O => \N__36988\,
            I => \N__36982\
        );

    \I__8939\ : InMux
    port map (
            O => \N__36987\,
            I => \N__36977\
        );

    \I__8938\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36977\
        );

    \I__8937\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36974\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__36982\,
            I => \N__36968\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36968\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__36974\,
            I => \N__36963\
        );

    \I__8933\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36960\
        );

    \I__8932\ : Span4Mux_v
    port map (
            O => \N__36968\,
            I => \N__36957\
        );

    \I__8931\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36954\
        );

    \I__8930\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36951\
        );

    \I__8929\ : Span4Mux_v
    port map (
            O => \N__36963\,
            I => \N__36946\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__36960\,
            I => \N__36946\
        );

    \I__8927\ : Sp12to4
    port map (
            O => \N__36957\,
            I => \N__36939\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__36954\,
            I => \N__36939\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__36951\,
            I => \N__36939\
        );

    \I__8924\ : Span4Mux_v
    port map (
            O => \N__36946\,
            I => \N__36936\
        );

    \I__8923\ : Span12Mux_h
    port map (
            O => \N__36939\,
            I => \N__36933\
        );

    \I__8922\ : Span4Mux_h
    port map (
            O => \N__36936\,
            I => \N__36930\
        );

    \I__8921\ : Span12Mux_v
    port map (
            O => \N__36933\,
            I => \N__36927\
        );

    \I__8920\ : Sp12to4
    port map (
            O => \N__36930\,
            I => \N__36924\
        );

    \I__8919\ : Odrv12
    port map (
            O => \N__36927\,
            I => port_address_in_0
        );

    \I__8918\ : Odrv12
    port map (
            O => \N__36924\,
            I => port_address_in_0
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__36919\,
            I => \N__36916\
        );

    \I__8916\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36913\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__36913\,
            I => \this_ppu.N_610\
        );

    \I__8914\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36907\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__36907\,
            I => \M_this_state_d_0_sqmuxa_2\
        );

    \I__8912\ : IoInMux
    port map (
            O => \N__36904\,
            I => \N__36901\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__36901\,
            I => \N__36898\
        );

    \I__8910\ : IoSpan4Mux
    port map (
            O => \N__36898\,
            I => \N__36895\
        );

    \I__8909\ : Span4Mux_s0_h
    port map (
            O => \N__36895\,
            I => \N__36890\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__36894\,
            I => \N__36887\
        );

    \I__8907\ : CascadeMux
    port map (
            O => \N__36893\,
            I => \N__36882\
        );

    \I__8906\ : Sp12to4
    port map (
            O => \N__36890\,
            I => \N__36879\
        );

    \I__8905\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36876\
        );

    \I__8904\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36872\
        );

    \I__8903\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36867\
        );

    \I__8902\ : InMux
    port map (
            O => \N__36882\,
            I => \N__36867\
        );

    \I__8901\ : Span12Mux_v
    port map (
            O => \N__36879\,
            I => \N__36864\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__36876\,
            I => \N__36861\
        );

    \I__8899\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36858\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__36872\,
            I => \N__36853\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__36867\,
            I => \N__36853\
        );

    \I__8896\ : Odrv12
    port map (
            O => \N__36864\,
            I => led_c_1
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__36861\,
            I => led_c_1
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__36858\,
            I => led_c_1
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__36853\,
            I => led_c_1
        );

    \I__8892\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36840\
        );

    \I__8891\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36837\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__36840\,
            I => \N_608\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__36837\,
            I => \N_608\
        );

    \I__8888\ : InMux
    port map (
            O => \N__36832\,
            I => \N__36826\
        );

    \I__8887\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36821\
        );

    \I__8886\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36821\
        );

    \I__8885\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36818\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__36826\,
            I => \M_this_substate_qZ0\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__36821\,
            I => \M_this_substate_qZ0\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__36818\,
            I => \M_this_substate_qZ0\
        );

    \I__8881\ : CascadeMux
    port map (
            O => \N__36811\,
            I => \N__36807\
        );

    \I__8880\ : InMux
    port map (
            O => \N__36810\,
            I => \N__36803\
        );

    \I__8879\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36800\
        );

    \I__8878\ : CascadeMux
    port map (
            O => \N__36806\,
            I => \N__36793\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__36803\,
            I => \N__36790\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__36800\,
            I => \N__36787\
        );

    \I__8875\ : InMux
    port map (
            O => \N__36799\,
            I => \N__36784\
        );

    \I__8874\ : CascadeMux
    port map (
            O => \N__36798\,
            I => \N__36781\
        );

    \I__8873\ : CascadeMux
    port map (
            O => \N__36797\,
            I => \N__36778\
        );

    \I__8872\ : InMux
    port map (
            O => \N__36796\,
            I => \N__36770\
        );

    \I__8871\ : InMux
    port map (
            O => \N__36793\,
            I => \N__36770\
        );

    \I__8870\ : Span4Mux_v
    port map (
            O => \N__36790\,
            I => \N__36767\
        );

    \I__8869\ : Span12Mux_v
    port map (
            O => \N__36787\,
            I => \N__36762\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__36784\,
            I => \N__36762\
        );

    \I__8867\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36757\
        );

    \I__8866\ : InMux
    port map (
            O => \N__36778\,
            I => \N__36757\
        );

    \I__8865\ : InMux
    port map (
            O => \N__36777\,
            I => \N__36750\
        );

    \I__8864\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36750\
        );

    \I__8863\ : InMux
    port map (
            O => \N__36775\,
            I => \N__36750\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__36770\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8861\ : Odrv4
    port map (
            O => \N__36767\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8860\ : Odrv12
    port map (
            O => \N__36762\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__36757\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__36750\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8857\ : InMux
    port map (
            O => \N__36739\,
            I => \N__36735\
        );

    \I__8856\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36732\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__36735\,
            I => \N__36728\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__36732\,
            I => \N__36723\
        );

    \I__8853\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36718\
        );

    \I__8852\ : Span4Mux_h
    port map (
            O => \N__36728\,
            I => \N__36715\
        );

    \I__8851\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36710\
        );

    \I__8850\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36710\
        );

    \I__8849\ : Span4Mux_v
    port map (
            O => \N__36723\,
            I => \N__36707\
        );

    \I__8848\ : InMux
    port map (
            O => \N__36722\,
            I => \N__36704\
        );

    \I__8847\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36701\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__36718\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8845\ : Odrv4
    port map (
            O => \N__36715\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__36710\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8843\ : Odrv4
    port map (
            O => \N__36707\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__36704\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__36701\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8840\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36684\
        );

    \I__8839\ : CascadeMux
    port map (
            O => \N__36687\,
            I => \N__36680\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__36684\,
            I => \N__36674\
        );

    \I__8837\ : InMux
    port map (
            O => \N__36683\,
            I => \N__36671\
        );

    \I__8836\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36664\
        );

    \I__8835\ : InMux
    port map (
            O => \N__36679\,
            I => \N__36661\
        );

    \I__8834\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36658\
        );

    \I__8833\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36653\
        );

    \I__8832\ : Span4Mux_h
    port map (
            O => \N__36674\,
            I => \N__36648\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36648\
        );

    \I__8830\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36643\
        );

    \I__8829\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36643\
        );

    \I__8828\ : InMux
    port map (
            O => \N__36668\,
            I => \N__36638\
        );

    \I__8827\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36638\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__36664\,
            I => \N__36635\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__36661\,
            I => \N__36632\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__36658\,
            I => \N__36629\
        );

    \I__8823\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36626\
        );

    \I__8822\ : InMux
    port map (
            O => \N__36656\,
            I => \N__36623\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__36653\,
            I => \N__36618\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__36648\,
            I => \N__36618\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__36643\,
            I => \N__36613\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__36638\,
            I => \N__36613\
        );

    \I__8817\ : Span12Mux_h
    port map (
            O => \N__36635\,
            I => \N__36610\
        );

    \I__8816\ : Odrv12
    port map (
            O => \N__36632\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__36629\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__36626\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__36623\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__36618\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__8811\ : Odrv4
    port map (
            O => \N__36613\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__8810\ : Odrv12
    port map (
            O => \N__36610\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__8809\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36592\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__36592\,
            I => \N__36589\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__36589\,
            I => \this_ppu.oam_cache.mem_10\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__36586\,
            I => \N__36583\
        );

    \I__8805\ : InMux
    port map (
            O => \N__36583\,
            I => \N__36578\
        );

    \I__8804\ : InMux
    port map (
            O => \N__36582\,
            I => \N__36575\
        );

    \I__8803\ : InMux
    port map (
            O => \N__36581\,
            I => \N__36572\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__36578\,
            I => \N__36569\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__36575\,
            I => \N__36563\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__36572\,
            I => \N__36563\
        );

    \I__8799\ : Span4Mux_h
    port map (
            O => \N__36569\,
            I => \N__36557\
        );

    \I__8798\ : InMux
    port map (
            O => \N__36568\,
            I => \N__36554\
        );

    \I__8797\ : Span4Mux_h
    port map (
            O => \N__36563\,
            I => \N__36551\
        );

    \I__8796\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36544\
        );

    \I__8795\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36544\
        );

    \I__8794\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36544\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__36557\,
            I => \this_ppu.un1_M_hoffset_q_5\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__36554\,
            I => \this_ppu.un1_M_hoffset_q_5\
        );

    \I__8791\ : Odrv4
    port map (
            O => \N__36551\,
            I => \this_ppu.un1_M_hoffset_q_5\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__36544\,
            I => \this_ppu.un1_M_hoffset_q_5\
        );

    \I__8789\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36532\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36529\
        );

    \I__8787\ : Span4Mux_v
    port map (
            O => \N__36529\,
            I => \N__36526\
        );

    \I__8786\ : Odrv4
    port map (
            O => \N__36526\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_18\
        );

    \I__8785\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36520\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__36520\,
            I => \N__36515\
        );

    \I__8783\ : InMux
    port map (
            O => \N__36519\,
            I => \N__36512\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__36518\,
            I => \N__36509\
        );

    \I__8781\ : Span4Mux_h
    port map (
            O => \N__36515\,
            I => \N__36505\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__36512\,
            I => \N__36502\
        );

    \I__8779\ : InMux
    port map (
            O => \N__36509\,
            I => \N__36499\
        );

    \I__8778\ : InMux
    port map (
            O => \N__36508\,
            I => \N__36496\
        );

    \I__8777\ : Odrv4
    port map (
            O => \N__36505\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8776\ : Odrv4
    port map (
            O => \N__36502\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__36499\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__36496\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8773\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36482\
        );

    \I__8772\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36479\
        );

    \I__8771\ : CascadeMux
    port map (
            O => \N__36485\,
            I => \N__36473\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__36482\,
            I => \N__36469\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36466\
        );

    \I__8768\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36463\
        );

    \I__8767\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36459\
        );

    \I__8766\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36453\
        );

    \I__8765\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36453\
        );

    \I__8764\ : InMux
    port map (
            O => \N__36472\,
            I => \N__36450\
        );

    \I__8763\ : Span4Mux_h
    port map (
            O => \N__36469\,
            I => \N__36445\
        );

    \I__8762\ : Span4Mux_v
    port map (
            O => \N__36466\,
            I => \N__36445\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__36463\,
            I => \N__36442\
        );

    \I__8760\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36439\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__36459\,
            I => \N__36436\
        );

    \I__8758\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36433\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__36453\,
            I => \N__36430\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__36450\,
            I => \N__36426\
        );

    \I__8755\ : Span4Mux_v
    port map (
            O => \N__36445\,
            I => \N__36423\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__36442\,
            I => \N__36420\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__36439\,
            I => \N__36415\
        );

    \I__8752\ : Span4Mux_h
    port map (
            O => \N__36436\,
            I => \N__36415\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__36433\,
            I => \N__36412\
        );

    \I__8750\ : Span4Mux_v
    port map (
            O => \N__36430\,
            I => \N__36409\
        );

    \I__8749\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36406\
        );

    \I__8748\ : Span12Mux_s10_v
    port map (
            O => \N__36426\,
            I => \N__36403\
        );

    \I__8747\ : Sp12to4
    port map (
            O => \N__36423\,
            I => \N__36400\
        );

    \I__8746\ : Sp12to4
    port map (
            O => \N__36420\,
            I => \N__36397\
        );

    \I__8745\ : Span4Mux_v
    port map (
            O => \N__36415\,
            I => \N__36394\
        );

    \I__8744\ : Span4Mux_h
    port map (
            O => \N__36412\,
            I => \N__36391\
        );

    \I__8743\ : Span4Mux_v
    port map (
            O => \N__36409\,
            I => \N__36388\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__36406\,
            I => \N__36385\
        );

    \I__8741\ : Span12Mux_v
    port map (
            O => \N__36403\,
            I => \N__36382\
        );

    \I__8740\ : Span12Mux_h
    port map (
            O => \N__36400\,
            I => \N__36379\
        );

    \I__8739\ : Span12Mux_h
    port map (
            O => \N__36397\,
            I => \N__36372\
        );

    \I__8738\ : Sp12to4
    port map (
            O => \N__36394\,
            I => \N__36372\
        );

    \I__8737\ : Sp12to4
    port map (
            O => \N__36391\,
            I => \N__36372\
        );

    \I__8736\ : Span4Mux_v
    port map (
            O => \N__36388\,
            I => \N__36367\
        );

    \I__8735\ : Span4Mux_v
    port map (
            O => \N__36385\,
            I => \N__36367\
        );

    \I__8734\ : Span12Mux_h
    port map (
            O => \N__36382\,
            I => \N__36362\
        );

    \I__8733\ : Span12Mux_v
    port map (
            O => \N__36379\,
            I => \N__36362\
        );

    \I__8732\ : Span12Mux_v
    port map (
            O => \N__36372\,
            I => \N__36359\
        );

    \I__8731\ : Span4Mux_h
    port map (
            O => \N__36367\,
            I => \N__36356\
        );

    \I__8730\ : Odrv12
    port map (
            O => \N__36362\,
            I => port_data_c_7
        );

    \I__8729\ : Odrv12
    port map (
            O => \N__36359\,
            I => port_data_c_7
        );

    \I__8728\ : Odrv4
    port map (
            O => \N__36356\,
            I => port_data_c_7
        );

    \I__8727\ : InMux
    port map (
            O => \N__36349\,
            I => \N__36346\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__36346\,
            I => \N__36343\
        );

    \I__8725\ : Odrv4
    port map (
            O => \N__36343\,
            I => \N_440\
        );

    \I__8724\ : InMux
    port map (
            O => \N__36340\,
            I => \N__36337\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__36337\,
            I => \N__36334\
        );

    \I__8722\ : Odrv4
    port map (
            O => \N__36334\,
            I => \N_437\
        );

    \I__8721\ : InMux
    port map (
            O => \N__36331\,
            I => \N__36328\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__36328\,
            I => \N__36325\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__36325\,
            I => \M_this_data_tmp_qZ0Z_22\
        );

    \I__8718\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36319\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__36319\,
            I => \N__36316\
        );

    \I__8716\ : Odrv12
    port map (
            O => \N__36316\,
            I => \M_this_oam_ram_write_data_22\
        );

    \I__8715\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36310\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__36310\,
            I => \N__36304\
        );

    \I__8713\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36301\
        );

    \I__8712\ : CascadeMux
    port map (
            O => \N__36308\,
            I => \N__36298\
        );

    \I__8711\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36295\
        );

    \I__8710\ : Span4Mux_v
    port map (
            O => \N__36304\,
            I => \N__36288\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__36301\,
            I => \N__36288\
        );

    \I__8708\ : InMux
    port map (
            O => \N__36298\,
            I => \N__36285\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__36295\,
            I => \N__36282\
        );

    \I__8706\ : CascadeMux
    port map (
            O => \N__36294\,
            I => \N__36279\
        );

    \I__8705\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36275\
        );

    \I__8704\ : Span4Mux_v
    port map (
            O => \N__36288\,
            I => \N__36270\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__36285\,
            I => \N__36270\
        );

    \I__8702\ : Span4Mux_v
    port map (
            O => \N__36282\,
            I => \N__36266\
        );

    \I__8701\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36263\
        );

    \I__8700\ : InMux
    port map (
            O => \N__36278\,
            I => \N__36259\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__36275\,
            I => \N__36256\
        );

    \I__8698\ : Span4Mux_v
    port map (
            O => \N__36270\,
            I => \N__36253\
        );

    \I__8697\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36250\
        );

    \I__8696\ : Span4Mux_v
    port map (
            O => \N__36266\,
            I => \N__36247\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__36263\,
            I => \N__36244\
        );

    \I__8694\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36241\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__36259\,
            I => \N__36238\
        );

    \I__8692\ : Sp12to4
    port map (
            O => \N__36256\,
            I => \N__36235\
        );

    \I__8691\ : Span4Mux_h
    port map (
            O => \N__36253\,
            I => \N__36230\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__36250\,
            I => \N__36230\
        );

    \I__8689\ : Sp12to4
    port map (
            O => \N__36247\,
            I => \N__36227\
        );

    \I__8688\ : Span4Mux_v
    port map (
            O => \N__36244\,
            I => \N__36224\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__36241\,
            I => \N__36221\
        );

    \I__8686\ : Span12Mux_h
    port map (
            O => \N__36238\,
            I => \N__36214\
        );

    \I__8685\ : Span12Mux_s9_v
    port map (
            O => \N__36235\,
            I => \N__36214\
        );

    \I__8684\ : Sp12to4
    port map (
            O => \N__36230\,
            I => \N__36214\
        );

    \I__8683\ : Span12Mux_h
    port map (
            O => \N__36227\,
            I => \N__36211\
        );

    \I__8682\ : Sp12to4
    port map (
            O => \N__36224\,
            I => \N__36208\
        );

    \I__8681\ : Span12Mux_h
    port map (
            O => \N__36221\,
            I => \N__36205\
        );

    \I__8680\ : Span12Mux_v
    port map (
            O => \N__36214\,
            I => \N__36202\
        );

    \I__8679\ : Span12Mux_v
    port map (
            O => \N__36211\,
            I => \N__36199\
        );

    \I__8678\ : Span12Mux_h
    port map (
            O => \N__36208\,
            I => \N__36196\
        );

    \I__8677\ : Span12Mux_v
    port map (
            O => \N__36205\,
            I => \N__36191\
        );

    \I__8676\ : Span12Mux_h
    port map (
            O => \N__36202\,
            I => \N__36191\
        );

    \I__8675\ : Odrv12
    port map (
            O => \N__36199\,
            I => port_data_c_6
        );

    \I__8674\ : Odrv12
    port map (
            O => \N__36196\,
            I => port_data_c_6
        );

    \I__8673\ : Odrv12
    port map (
            O => \N__36191\,
            I => port_data_c_6
        );

    \I__8672\ : InMux
    port map (
            O => \N__36184\,
            I => \N__36181\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__36181\,
            I => \N__36178\
        );

    \I__8670\ : Span4Mux_h
    port map (
            O => \N__36178\,
            I => \N__36175\
        );

    \I__8669\ : Odrv4
    port map (
            O => \N__36175\,
            I => \N_439\
        );

    \I__8668\ : CEMux
    port map (
            O => \N__36172\,
            I => \N__36169\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__36169\,
            I => \N__36165\
        );

    \I__8666\ : CEMux
    port map (
            O => \N__36168\,
            I => \N__36162\
        );

    \I__8665\ : Odrv4
    port map (
            O => \N__36165\,
            I => \this_spr_ram.mem_WE_2\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__36162\,
            I => \this_spr_ram.mem_WE_2\
        );

    \I__8663\ : CEMux
    port map (
            O => \N__36157\,
            I => \N__36153\
        );

    \I__8662\ : CEMux
    port map (
            O => \N__36156\,
            I => \N__36150\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__36153\,
            I => \this_spr_ram.mem_WE_4\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__36150\,
            I => \this_spr_ram.mem_WE_4\
        );

    \I__8659\ : InMux
    port map (
            O => \N__36145\,
            I => \N__36142\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__36142\,
            I => \this_spr_ram.mem_out_bus5_1\
        );

    \I__8657\ : InMux
    port map (
            O => \N__36139\,
            I => \N__36136\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__36136\,
            I => \N__36133\
        );

    \I__8655\ : Span4Mux_h
    port map (
            O => \N__36133\,
            I => \N__36130\
        );

    \I__8654\ : Odrv4
    port map (
            O => \N__36130\,
            I => \this_spr_ram.mem_out_bus1_1\
        );

    \I__8653\ : InMux
    port map (
            O => \N__36127\,
            I => \N__36124\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__36124\,
            I => \N__36121\
        );

    \I__8651\ : Span12Mux_s10_v
    port map (
            O => \N__36121\,
            I => \N__36118\
        );

    \I__8650\ : Odrv12
    port map (
            O => \N__36118\,
            I => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\
        );

    \I__8649\ : CEMux
    port map (
            O => \N__36115\,
            I => \N__36111\
        );

    \I__8648\ : CEMux
    port map (
            O => \N__36114\,
            I => \N__36108\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__36111\,
            I => \N__36105\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__36108\,
            I => \N__36102\
        );

    \I__8645\ : Span4Mux_v
    port map (
            O => \N__36105\,
            I => \N__36099\
        );

    \I__8644\ : Span4Mux_h
    port map (
            O => \N__36102\,
            I => \N__36096\
        );

    \I__8643\ : Span4Mux_v
    port map (
            O => \N__36099\,
            I => \N__36093\
        );

    \I__8642\ : Span4Mux_v
    port map (
            O => \N__36096\,
            I => \N__36090\
        );

    \I__8641\ : Odrv4
    port map (
            O => \N__36093\,
            I => \this_spr_ram.mem_WE_14\
        );

    \I__8640\ : Odrv4
    port map (
            O => \N__36090\,
            I => \this_spr_ram.mem_WE_14\
        );

    \I__8639\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36082\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__36082\,
            I => \N__36079\
        );

    \I__8637\ : Span4Mux_v
    port map (
            O => \N__36079\,
            I => \N__36076\
        );

    \I__8636\ : Odrv4
    port map (
            O => \N__36076\,
            I => \M_this_oam_ram_write_data_7\
        );

    \I__8635\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36070\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__36070\,
            I => \M_this_data_tmp_qZ0Z_7\
        );

    \I__8633\ : InMux
    port map (
            O => \N__36067\,
            I => \N__36064\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__36064\,
            I => \N__36061\
        );

    \I__8631\ : Span4Mux_h
    port map (
            O => \N__36061\,
            I => \N__36058\
        );

    \I__8630\ : Odrv4
    port map (
            O => \N__36058\,
            I => \M_this_oam_ram_write_data_3\
        );

    \I__8629\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36052\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__36052\,
            I => \M_this_data_tmp_qZ0Z_3\
        );

    \I__8627\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36046\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36043\
        );

    \I__8625\ : Span4Mux_h
    port map (
            O => \N__36043\,
            I => \N__36040\
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__36040\,
            I => \M_this_oam_ram_write_data_4\
        );

    \I__8623\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36034\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__36034\,
            I => \M_this_data_tmp_qZ0Z_4\
        );

    \I__8621\ : CEMux
    port map (
            O => \N__36031\,
            I => \N__36025\
        );

    \I__8620\ : CEMux
    port map (
            O => \N__36030\,
            I => \N__36022\
        );

    \I__8619\ : CEMux
    port map (
            O => \N__36029\,
            I => \N__36019\
        );

    \I__8618\ : CEMux
    port map (
            O => \N__36028\,
            I => \N__36016\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__36025\,
            I => \N__36012\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__36022\,
            I => \N__36009\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__36019\,
            I => \N__36004\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__36016\,
            I => \N__36004\
        );

    \I__8613\ : CEMux
    port map (
            O => \N__36015\,
            I => \N__36001\
        );

    \I__8612\ : Span4Mux_v
    port map (
            O => \N__36012\,
            I => \N__35998\
        );

    \I__8611\ : Span4Mux_h
    port map (
            O => \N__36009\,
            I => \N__35995\
        );

    \I__8610\ : Span4Mux_v
    port map (
            O => \N__36004\,
            I => \N__35990\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__36001\,
            I => \N__35990\
        );

    \I__8608\ : Span4Mux_h
    port map (
            O => \N__35998\,
            I => \N__35987\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__35995\,
            I => \N__35984\
        );

    \I__8606\ : Span4Mux_h
    port map (
            O => \N__35990\,
            I => \N__35981\
        );

    \I__8605\ : Odrv4
    port map (
            O => \N__35987\,
            I => \N_1302_0\
        );

    \I__8604\ : Odrv4
    port map (
            O => \N__35984\,
            I => \N_1302_0\
        );

    \I__8603\ : Odrv4
    port map (
            O => \N__35981\,
            I => \N_1302_0\
        );

    \I__8602\ : InMux
    port map (
            O => \N__35974\,
            I => \N__35971\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__35971\,
            I => \N__35968\
        );

    \I__8600\ : Odrv12
    port map (
            O => \N__35968\,
            I => \M_this_data_tmp_qZ0Z_23\
        );

    \I__8599\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35962\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__35962\,
            I => \N__35959\
        );

    \I__8597\ : Span4Mux_v
    port map (
            O => \N__35959\,
            I => \N__35956\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__35956\,
            I => \M_this_oam_ram_write_data_23\
        );

    \I__8595\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35950\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__35950\,
            I => \N__35947\
        );

    \I__8593\ : Span4Mux_v
    port map (
            O => \N__35947\,
            I => \N__35944\
        );

    \I__8592\ : Odrv4
    port map (
            O => \N__35944\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_17\
        );

    \I__8591\ : InMux
    port map (
            O => \N__35941\,
            I => \N__35938\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35935\
        );

    \I__8589\ : Odrv12
    port map (
            O => \N__35935\,
            I => \this_ppu.oam_cache.mem_11\
        );

    \I__8588\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35928\
        );

    \I__8587\ : InMux
    port map (
            O => \N__35931\,
            I => \N__35925\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__35928\,
            I => \N__35918\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__35925\,
            I => \N__35918\
        );

    \I__8584\ : CascadeMux
    port map (
            O => \N__35924\,
            I => \N__35915\
        );

    \I__8583\ : CascadeMux
    port map (
            O => \N__35923\,
            I => \N__35912\
        );

    \I__8582\ : Span4Mux_h
    port map (
            O => \N__35918\,
            I => \N__35909\
        );

    \I__8581\ : InMux
    port map (
            O => \N__35915\,
            I => \N__35904\
        );

    \I__8580\ : InMux
    port map (
            O => \N__35912\,
            I => \N__35904\
        );

    \I__8579\ : Odrv4
    port map (
            O => \N__35909\,
            I => \this_ppu.un1_M_hoffset_q_6\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__35904\,
            I => \this_ppu.un1_M_hoffset_q_6\
        );

    \I__8577\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35894\
        );

    \I__8576\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35891\
        );

    \I__8575\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35888\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35878\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__35891\,
            I => \N__35878\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__35888\,
            I => \N__35878\
        );

    \I__8571\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35875\
        );

    \I__8570\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35872\
        );

    \I__8569\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35869\
        );

    \I__8568\ : Span4Mux_v
    port map (
            O => \N__35878\,
            I => \N__35864\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__35875\,
            I => \N__35864\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__35872\,
            I => \N__35861\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__35869\,
            I => \N__35858\
        );

    \I__8564\ : Span4Mux_h
    port map (
            O => \N__35864\,
            I => \N__35855\
        );

    \I__8563\ : Odrv4
    port map (
            O => \N__35861\,
            I => \this_ppu.M_hoffset_qZ0Z_1\
        );

    \I__8562\ : Odrv4
    port map (
            O => \N__35858\,
            I => \this_ppu.M_hoffset_qZ0Z_1\
        );

    \I__8561\ : Odrv4
    port map (
            O => \N__35855\,
            I => \this_ppu.M_hoffset_qZ0Z_1\
        );

    \I__8560\ : InMux
    port map (
            O => \N__35848\,
            I => \N__35843\
        );

    \I__8559\ : InMux
    port map (
            O => \N__35847\,
            I => \N__35840\
        );

    \I__8558\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35837\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35833\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__35840\,
            I => \N__35827\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__35837\,
            I => \N__35827\
        );

    \I__8554\ : CascadeMux
    port map (
            O => \N__35836\,
            I => \N__35821\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__35833\,
            I => \N__35817\
        );

    \I__8552\ : InMux
    port map (
            O => \N__35832\,
            I => \N__35814\
        );

    \I__8551\ : Span4Mux_h
    port map (
            O => \N__35827\,
            I => \N__35811\
        );

    \I__8550\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35808\
        );

    \I__8549\ : InMux
    port map (
            O => \N__35825\,
            I => \N__35805\
        );

    \I__8548\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35798\
        );

    \I__8547\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35798\
        );

    \I__8546\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35798\
        );

    \I__8545\ : Odrv4
    port map (
            O => \N__35817\,
            I => \this_ppu.un1_M_hoffset_q_4\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__35814\,
            I => \this_ppu.un1_M_hoffset_q_4\
        );

    \I__8543\ : Odrv4
    port map (
            O => \N__35811\,
            I => \this_ppu.un1_M_hoffset_q_4\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__35808\,
            I => \this_ppu.un1_M_hoffset_q_4\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__35805\,
            I => \this_ppu.un1_M_hoffset_q_4\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__35798\,
            I => \this_ppu.un1_M_hoffset_q_4\
        );

    \I__8539\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35778\
        );

    \I__8538\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35775\
        );

    \I__8537\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35772\
        );

    \I__8536\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35769\
        );

    \I__8535\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35766\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35763\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35754\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__35772\,
            I => \N__35754\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__35769\,
            I => \N__35754\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__35766\,
            I => \N__35746\
        );

    \I__8529\ : Span4Mux_h
    port map (
            O => \N__35763\,
            I => \N__35743\
        );

    \I__8528\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35740\
        );

    \I__8527\ : InMux
    port map (
            O => \N__35761\,
            I => \N__35737\
        );

    \I__8526\ : Span4Mux_v
    port map (
            O => \N__35754\,
            I => \N__35734\
        );

    \I__8525\ : InMux
    port map (
            O => \N__35753\,
            I => \N__35731\
        );

    \I__8524\ : InMux
    port map (
            O => \N__35752\,
            I => \N__35728\
        );

    \I__8523\ : InMux
    port map (
            O => \N__35751\,
            I => \N__35721\
        );

    \I__8522\ : InMux
    port map (
            O => \N__35750\,
            I => \N__35721\
        );

    \I__8521\ : InMux
    port map (
            O => \N__35749\,
            I => \N__35721\
        );

    \I__8520\ : Odrv12
    port map (
            O => \N__35746\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8519\ : Odrv4
    port map (
            O => \N__35743\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__35740\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__35737\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__35734\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__35731\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__35728\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__35721\,
            I => \this_ppu.un1_M_hoffset_q_0\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__35704\,
            I => \N__35701\
        );

    \I__8511\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35698\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__35698\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNOZ0\
        );

    \I__8509\ : InMux
    port map (
            O => \N__35695\,
            I => \N__35683\
        );

    \I__8508\ : InMux
    port map (
            O => \N__35694\,
            I => \N__35683\
        );

    \I__8507\ : InMux
    port map (
            O => \N__35693\,
            I => \N__35683\
        );

    \I__8506\ : InMux
    port map (
            O => \N__35692\,
            I => \N__35683\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__35683\,
            I => \this_ppu.un1_oam_data_1_4_c5_0\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__35680\,
            I => \N__35676\
        );

    \I__8503\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35672\
        );

    \I__8502\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35666\
        );

    \I__8501\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35666\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__35672\,
            I => \N__35663\
        );

    \I__8499\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35660\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__35666\,
            I => \N__35657\
        );

    \I__8497\ : Span4Mux_h
    port map (
            O => \N__35663\,
            I => \N__35654\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__35660\,
            I => \N__35651\
        );

    \I__8495\ : Span4Mux_h
    port map (
            O => \N__35657\,
            I => \N__35648\
        );

    \I__8494\ : Span4Mux_v
    port map (
            O => \N__35654\,
            I => \N__35645\
        );

    \I__8493\ : Span4Mux_h
    port map (
            O => \N__35651\,
            I => \N__35640\
        );

    \I__8492\ : Span4Mux_v
    port map (
            O => \N__35648\,
            I => \N__35640\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__35645\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__35640\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__8489\ : InMux
    port map (
            O => \N__35635\,
            I => \N__35632\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__35632\,
            I => \N__35629\
        );

    \I__8487\ : Span4Mux_h
    port map (
            O => \N__35629\,
            I => \N__35626\
        );

    \I__8486\ : Odrv4
    port map (
            O => \N__35626\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_23\
        );

    \I__8485\ : InMux
    port map (
            O => \N__35623\,
            I => \N__35620\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__35620\,
            I => \N__35615\
        );

    \I__8483\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35612\
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__35618\,
            I => \N__35609\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__35615\,
            I => \N__35603\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__35612\,
            I => \N__35603\
        );

    \I__8479\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35599\
        );

    \I__8478\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35595\
        );

    \I__8477\ : Span4Mux_h
    port map (
            O => \N__35603\,
            I => \N__35592\
        );

    \I__8476\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35589\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__35599\,
            I => \N__35585\
        );

    \I__8474\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35582\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__35595\,
            I => \N__35579\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__35592\,
            I => \N__35576\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__35589\,
            I => \N__35573\
        );

    \I__8470\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35570\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__35585\,
            I => \N__35564\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__35582\,
            I => \N__35564\
        );

    \I__8467\ : Span4Mux_h
    port map (
            O => \N__35579\,
            I => \N__35560\
        );

    \I__8466\ : Span4Mux_v
    port map (
            O => \N__35576\,
            I => \N__35553\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__35573\,
            I => \N__35553\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__35570\,
            I => \N__35553\
        );

    \I__8463\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35550\
        );

    \I__8462\ : Span4Mux_v
    port map (
            O => \N__35564\,
            I => \N__35547\
        );

    \I__8461\ : InMux
    port map (
            O => \N__35563\,
            I => \N__35544\
        );

    \I__8460\ : Span4Mux_v
    port map (
            O => \N__35560\,
            I => \N__35539\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__35553\,
            I => \N__35539\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__35550\,
            I => \N__35536\
        );

    \I__8457\ : Sp12to4
    port map (
            O => \N__35547\,
            I => \N__35531\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__35544\,
            I => \N__35531\
        );

    \I__8455\ : Span4Mux_v
    port map (
            O => \N__35539\,
            I => \N__35528\
        );

    \I__8454\ : Span12Mux_h
    port map (
            O => \N__35536\,
            I => \N__35525\
        );

    \I__8453\ : Span12Mux_h
    port map (
            O => \N__35531\,
            I => \N__35522\
        );

    \I__8452\ : Span4Mux_v
    port map (
            O => \N__35528\,
            I => \N__35519\
        );

    \I__8451\ : Odrv12
    port map (
            O => \N__35525\,
            I => port_data_c_0
        );

    \I__8450\ : Odrv12
    port map (
            O => \N__35522\,
            I => port_data_c_0
        );

    \I__8449\ : Odrv4
    port map (
            O => \N__35519\,
            I => port_data_c_0
        );

    \I__8448\ : InMux
    port map (
            O => \N__35512\,
            I => \N__35508\
        );

    \I__8447\ : InMux
    port map (
            O => \N__35511\,
            I => \N__35505\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35499\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__35505\,
            I => \N__35499\
        );

    \I__8444\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35495\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__35499\,
            I => \N__35492\
        );

    \I__8442\ : InMux
    port map (
            O => \N__35498\,
            I => \N__35488\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__35495\,
            I => \N__35485\
        );

    \I__8440\ : Span4Mux_v
    port map (
            O => \N__35492\,
            I => \N__35482\
        );

    \I__8439\ : InMux
    port map (
            O => \N__35491\,
            I => \N__35479\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__35488\,
            I => \N__35476\
        );

    \I__8437\ : Span4Mux_v
    port map (
            O => \N__35485\,
            I => \N__35472\
        );

    \I__8436\ : Span4Mux_v
    port map (
            O => \N__35482\,
            I => \N__35464\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__35479\,
            I => \N__35464\
        );

    \I__8434\ : Span4Mux_v
    port map (
            O => \N__35476\,
            I => \N__35461\
        );

    \I__8433\ : InMux
    port map (
            O => \N__35475\,
            I => \N__35458\
        );

    \I__8432\ : Span4Mux_v
    port map (
            O => \N__35472\,
            I => \N__35455\
        );

    \I__8431\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35450\
        );

    \I__8430\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35450\
        );

    \I__8429\ : InMux
    port map (
            O => \N__35469\,
            I => \N__35447\
        );

    \I__8428\ : Span4Mux_v
    port map (
            O => \N__35464\,
            I => \N__35444\
        );

    \I__8427\ : Sp12to4
    port map (
            O => \N__35461\,
            I => \N__35439\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__35458\,
            I => \N__35439\
        );

    \I__8425\ : Sp12to4
    port map (
            O => \N__35455\,
            I => \N__35432\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__35450\,
            I => \N__35432\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35432\
        );

    \I__8422\ : Span4Mux_v
    port map (
            O => \N__35444\,
            I => \N__35429\
        );

    \I__8421\ : Span12Mux_h
    port map (
            O => \N__35439\,
            I => \N__35426\
        );

    \I__8420\ : Span12Mux_h
    port map (
            O => \N__35432\,
            I => \N__35423\
        );

    \I__8419\ : IoSpan4Mux
    port map (
            O => \N__35429\,
            I => \N__35420\
        );

    \I__8418\ : Odrv12
    port map (
            O => \N__35426\,
            I => port_data_c_1
        );

    \I__8417\ : Odrv12
    port map (
            O => \N__35423\,
            I => port_data_c_1
        );

    \I__8416\ : Odrv4
    port map (
            O => \N__35420\,
            I => port_data_c_1
        );

    \I__8415\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35410\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__35410\,
            I => \N__35407\
        );

    \I__8413\ : Span4Mux_h
    port map (
            O => \N__35407\,
            I => \N__35404\
        );

    \I__8412\ : Odrv4
    port map (
            O => \N__35404\,
            I => \this_ppu.oam_cache.mem_16\
        );

    \I__8411\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35397\
        );

    \I__8410\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35394\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__35397\,
            I => \N__35391\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__35394\,
            I => \N__35388\
        );

    \I__8407\ : Span4Mux_h
    port map (
            O => \N__35391\,
            I => \N__35385\
        );

    \I__8406\ : Odrv12
    port map (
            O => \N__35388\,
            I => \this_ppu.M_oam_cache_read_data_16\
        );

    \I__8405\ : Odrv4
    port map (
            O => \N__35385\,
            I => \this_ppu.M_oam_cache_read_data_16\
        );

    \I__8404\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35377\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35374\
        );

    \I__8402\ : Span4Mux_v
    port map (
            O => \N__35374\,
            I => \N__35371\
        );

    \I__8401\ : Span4Mux_h
    port map (
            O => \N__35371\,
            I => \N__35368\
        );

    \I__8400\ : Odrv4
    port map (
            O => \N__35368\,
            I => \M_this_data_tmp_qZ0Z_20\
        );

    \I__8399\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35362\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__35362\,
            I => \N__35359\
        );

    \I__8397\ : Span4Mux_h
    port map (
            O => \N__35359\,
            I => \N__35356\
        );

    \I__8396\ : Span4Mux_v
    port map (
            O => \N__35356\,
            I => \N__35353\
        );

    \I__8395\ : Odrv4
    port map (
            O => \N__35353\,
            I => \M_this_oam_ram_write_data_20\
        );

    \I__8394\ : InMux
    port map (
            O => \N__35350\,
            I => \N__35347\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__35347\,
            I => \N__35344\
        );

    \I__8392\ : Span4Mux_v
    port map (
            O => \N__35344\,
            I => \N__35341\
        );

    \I__8391\ : Odrv4
    port map (
            O => \N__35341\,
            I => \this_ppu.oam_cache.mem_12\
        );

    \I__8390\ : CascadeMux
    port map (
            O => \N__35338\,
            I => \N__35335\
        );

    \I__8389\ : InMux
    port map (
            O => \N__35335\,
            I => \N__35329\
        );

    \I__8388\ : InMux
    port map (
            O => \N__35334\,
            I => \N__35326\
        );

    \I__8387\ : InMux
    port map (
            O => \N__35333\,
            I => \N__35321\
        );

    \I__8386\ : InMux
    port map (
            O => \N__35332\,
            I => \N__35318\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__35329\,
            I => \N__35315\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__35326\,
            I => \N__35312\
        );

    \I__8383\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35309\
        );

    \I__8382\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35306\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__35321\,
            I => \N__35303\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__35318\,
            I => \N__35300\
        );

    \I__8379\ : Span4Mux_v
    port map (
            O => \N__35315\,
            I => \N__35297\
        );

    \I__8378\ : Span4Mux_h
    port map (
            O => \N__35312\,
            I => \N__35292\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__35309\,
            I => \N__35292\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__35306\,
            I => \N__35287\
        );

    \I__8375\ : Span4Mux_v
    port map (
            O => \N__35303\,
            I => \N__35287\
        );

    \I__8374\ : Span4Mux_h
    port map (
            O => \N__35300\,
            I => \N__35284\
        );

    \I__8373\ : Odrv4
    port map (
            O => \N__35297\,
            I => \this_ppu.M_hoffset_qZ0Z_2\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__35292\,
            I => \this_ppu.M_hoffset_qZ0Z_2\
        );

    \I__8371\ : Odrv4
    port map (
            O => \N__35287\,
            I => \this_ppu.M_hoffset_qZ0Z_2\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__35284\,
            I => \this_ppu.M_hoffset_qZ0Z_2\
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__35275\,
            I => \N__35272\
        );

    \I__8368\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35269\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__35269\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNOZ0\
        );

    \I__8366\ : InMux
    port map (
            O => \N__35266\,
            I => \N__35263\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__35263\,
            I => \N__35260\
        );

    \I__8364\ : Span4Mux_h
    port map (
            O => \N__35260\,
            I => \N__35257\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__35257\,
            I => \this_ppu.oam_cache.mem_9\
        );

    \I__8362\ : InMux
    port map (
            O => \N__35254\,
            I => \N__35251\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__35251\,
            I => \N__35248\
        );

    \I__8360\ : Span4Mux_h
    port map (
            O => \N__35248\,
            I => \N__35245\
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__35245\,
            I => \this_ppu.oam_cache.mem_8\
        );

    \I__8358\ : InMux
    port map (
            O => \N__35242\,
            I => \N__35239\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__35239\,
            I => \N__35236\
        );

    \I__8356\ : Span4Mux_h
    port map (
            O => \N__35236\,
            I => \N__35233\
        );

    \I__8355\ : Odrv4
    port map (
            O => \N__35233\,
            I => \this_ppu.oam_cache.mem_13\
        );

    \I__8354\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35221\
        );

    \I__8353\ : InMux
    port map (
            O => \N__35229\,
            I => \N__35221\
        );

    \I__8352\ : InMux
    port map (
            O => \N__35228\,
            I => \N__35216\
        );

    \I__8351\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35216\
        );

    \I__8350\ : InMux
    port map (
            O => \N__35226\,
            I => \N__35213\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__35221\,
            I => \this_ppu.un1_M_oam_cache_read_data_c4\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__35216\,
            I => \this_ppu.un1_M_oam_cache_read_data_c4\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__35213\,
            I => \this_ppu.un1_M_oam_cache_read_data_c4\
        );

    \I__8346\ : CascadeMux
    port map (
            O => \N__35206\,
            I => \N__35203\
        );

    \I__8345\ : CascadeBuf
    port map (
            O => \N__35203\,
            I => \N__35200\
        );

    \I__8344\ : CascadeMux
    port map (
            O => \N__35200\,
            I => \N__35196\
        );

    \I__8343\ : CascadeMux
    port map (
            O => \N__35199\,
            I => \N__35193\
        );

    \I__8342\ : InMux
    port map (
            O => \N__35196\,
            I => \N__35189\
        );

    \I__8341\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35186\
        );

    \I__8340\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35183\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__35189\,
            I => \N__35179\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__35186\,
            I => \N__35175\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__35183\,
            I => \N__35171\
        );

    \I__8336\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35168\
        );

    \I__8335\ : Span4Mux_h
    port map (
            O => \N__35179\,
            I => \N__35165\
        );

    \I__8334\ : InMux
    port map (
            O => \N__35178\,
            I => \N__35162\
        );

    \I__8333\ : Span4Mux_h
    port map (
            O => \N__35175\,
            I => \N__35159\
        );

    \I__8332\ : InMux
    port map (
            O => \N__35174\,
            I => \N__35156\
        );

    \I__8331\ : Span4Mux_v
    port map (
            O => \N__35171\,
            I => \N__35151\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__35168\,
            I => \N__35151\
        );

    \I__8329\ : Span4Mux_h
    port map (
            O => \N__35165\,
            I => \N__35148\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__35162\,
            I => \N__35141\
        );

    \I__8327\ : Span4Mux_h
    port map (
            O => \N__35159\,
            I => \N__35141\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__35156\,
            I => \N__35141\
        );

    \I__8325\ : Span4Mux_h
    port map (
            O => \N__35151\,
            I => \N__35136\
        );

    \I__8324\ : Span4Mux_h
    port map (
            O => \N__35148\,
            I => \N__35136\
        );

    \I__8323\ : Span4Mux_v
    port map (
            O => \N__35141\,
            I => \N__35133\
        );

    \I__8322\ : Span4Mux_v
    port map (
            O => \N__35136\,
            I => \N__35130\
        );

    \I__8321\ : Odrv4
    port map (
            O => \N__35133\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__35130\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__8319\ : InMux
    port map (
            O => \N__35125\,
            I => \N__35121\
        );

    \I__8318\ : InMux
    port map (
            O => \N__35124\,
            I => \N__35118\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__35112\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__35118\,
            I => \N__35112\
        );

    \I__8315\ : InMux
    port map (
            O => \N__35117\,
            I => \N__35109\
        );

    \I__8314\ : Span4Mux_h
    port map (
            O => \N__35112\,
            I => \N__35103\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__35109\,
            I => \N__35100\
        );

    \I__8312\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35097\
        );

    \I__8311\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35094\
        );

    \I__8310\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35091\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__35103\,
            I => \this_ppu.un1_M_hoffset_q_8\
        );

    \I__8308\ : Odrv4
    port map (
            O => \N__35100\,
            I => \this_ppu.un1_M_hoffset_q_8\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__35097\,
            I => \this_ppu.un1_M_hoffset_q_8\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__35094\,
            I => \this_ppu.un1_M_hoffset_q_8\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__35091\,
            I => \this_ppu.un1_M_hoffset_q_8\
        );

    \I__8304\ : CascadeMux
    port map (
            O => \N__35080\,
            I => \this_ppu.un1_M_oam_cache_read_data_c4_cascade_\
        );

    \I__8303\ : InMux
    port map (
            O => \N__35077\,
            I => \N__35074\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__35074\,
            I => \N__35069\
        );

    \I__8301\ : CascadeMux
    port map (
            O => \N__35073\,
            I => \N__35066\
        );

    \I__8300\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35058\
        );

    \I__8299\ : Span4Mux_h
    port map (
            O => \N__35069\,
            I => \N__35055\
        );

    \I__8298\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35050\
        );

    \I__8297\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35050\
        );

    \I__8296\ : InMux
    port map (
            O => \N__35064\,
            I => \N__35047\
        );

    \I__8295\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35042\
        );

    \I__8294\ : InMux
    port map (
            O => \N__35062\,
            I => \N__35042\
        );

    \I__8293\ : InMux
    port map (
            O => \N__35061\,
            I => \N__35039\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__35058\,
            I => \this_ppu.un1_M_hoffset_q_7\
        );

    \I__8291\ : Odrv4
    port map (
            O => \N__35055\,
            I => \this_ppu.un1_M_hoffset_q_7\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__35050\,
            I => \this_ppu.un1_M_hoffset_q_7\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__35047\,
            I => \this_ppu.un1_M_hoffset_q_7\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__35042\,
            I => \this_ppu.un1_M_hoffset_q_7\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__35039\,
            I => \this_ppu.un1_M_hoffset_q_7\
        );

    \I__8286\ : InMux
    port map (
            O => \N__35026\,
            I => \N__35023\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__35023\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNOZ0\
        );

    \I__8284\ : InMux
    port map (
            O => \N__35020\,
            I => \N__35017\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__35017\,
            I => \N__35014\
        );

    \I__8282\ : Span4Mux_h
    port map (
            O => \N__35014\,
            I => \N__35010\
        );

    \I__8281\ : InMux
    port map (
            O => \N__35013\,
            I => \N__35007\
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__35010\,
            I => \this_ppu.read_data_RNI80ET_11\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__35007\,
            I => \this_ppu.read_data_RNI80ET_11\
        );

    \I__8278\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34999\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__34999\,
            I => \N__34996\
        );

    \I__8276\ : Span4Mux_h
    port map (
            O => \N__34996\,
            I => \N__34993\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__34993\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__8274\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34987\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34984\
        );

    \I__8272\ : Odrv4
    port map (
            O => \N__34984\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_11\
        );

    \I__8271\ : InMux
    port map (
            O => \N__34981\,
            I => \N__34978\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__34978\,
            I => \N__34972\
        );

    \I__8269\ : InMux
    port map (
            O => \N__34977\,
            I => \N__34969\
        );

    \I__8268\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34963\
        );

    \I__8267\ : InMux
    port map (
            O => \N__34975\,
            I => \N__34959\
        );

    \I__8266\ : Span4Mux_v
    port map (
            O => \N__34972\,
            I => \N__34951\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34951\
        );

    \I__8264\ : InMux
    port map (
            O => \N__34968\,
            I => \N__34948\
        );

    \I__8263\ : InMux
    port map (
            O => \N__34967\,
            I => \N__34945\
        );

    \I__8262\ : InMux
    port map (
            O => \N__34966\,
            I => \N__34942\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34937\
        );

    \I__8260\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34934\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__34959\,
            I => \N__34931\
        );

    \I__8258\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34924\
        );

    \I__8257\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34924\
        );

    \I__8256\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34924\
        );

    \I__8255\ : Span4Mux_v
    port map (
            O => \N__34951\,
            I => \N__34918\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__34948\,
            I => \N__34918\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__34945\,
            I => \N__34913\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__34942\,
            I => \N__34913\
        );

    \I__8251\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34908\
        );

    \I__8250\ : InMux
    port map (
            O => \N__34940\,
            I => \N__34908\
        );

    \I__8249\ : Span4Mux_v
    port map (
            O => \N__34937\,
            I => \N__34903\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__34934\,
            I => \N__34903\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__34931\,
            I => \N__34898\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__34924\,
            I => \N__34898\
        );

    \I__8245\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34895\
        );

    \I__8244\ : Span4Mux_v
    port map (
            O => \N__34918\,
            I => \N__34892\
        );

    \I__8243\ : Span4Mux_h
    port map (
            O => \N__34913\,
            I => \N__34889\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34886\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__34903\,
            I => \N__34883\
        );

    \I__8240\ : Span4Mux_h
    port map (
            O => \N__34898\,
            I => \N__34880\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__34895\,
            I => \N__34877\
        );

    \I__8238\ : Span4Mux_h
    port map (
            O => \N__34892\,
            I => \N__34874\
        );

    \I__8237\ : Span4Mux_v
    port map (
            O => \N__34889\,
            I => \N__34869\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__34886\,
            I => \N__34869\
        );

    \I__8235\ : Odrv4
    port map (
            O => \N__34883\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__34880\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__8233\ : Odrv12
    port map (
            O => \N__34877\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__34874\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__34869\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__8230\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34854\
        );

    \I__8229\ : CascadeMux
    port map (
            O => \N__34857\,
            I => \N__34851\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__34854\,
            I => \N__34847\
        );

    \I__8227\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34844\
        );

    \I__8226\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34840\
        );

    \I__8225\ : Span4Mux_h
    port map (
            O => \N__34847\,
            I => \N__34834\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__34844\,
            I => \N__34834\
        );

    \I__8223\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34831\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__34840\,
            I => \N__34828\
        );

    \I__8221\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34825\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__34834\,
            I => \N__34822\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__34831\,
            I => \N__34817\
        );

    \I__8218\ : Span4Mux_v
    port map (
            O => \N__34828\,
            I => \N__34817\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__34825\,
            I => \this_ppu.vspr\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__34822\,
            I => \this_ppu.vspr\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__34817\,
            I => \this_ppu.vspr\
        );

    \I__8214\ : CascadeMux
    port map (
            O => \N__34810\,
            I => \N__34804\
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__34809\,
            I => \N__34801\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__34808\,
            I => \N__34789\
        );

    \I__8211\ : CascadeMux
    port map (
            O => \N__34807\,
            I => \N__34786\
        );

    \I__8210\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34782\
        );

    \I__8209\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34779\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__34800\,
            I => \N__34776\
        );

    \I__8207\ : CascadeMux
    port map (
            O => \N__34799\,
            I => \N__34773\
        );

    \I__8206\ : CascadeMux
    port map (
            O => \N__34798\,
            I => \N__34770\
        );

    \I__8205\ : CascadeMux
    port map (
            O => \N__34797\,
            I => \N__34767\
        );

    \I__8204\ : CascadeMux
    port map (
            O => \N__34796\,
            I => \N__34764\
        );

    \I__8203\ : CascadeMux
    port map (
            O => \N__34795\,
            I => \N__34761\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__34794\,
            I => \N__34757\
        );

    \I__8201\ : CascadeMux
    port map (
            O => \N__34793\,
            I => \N__34754\
        );

    \I__8200\ : CascadeMux
    port map (
            O => \N__34792\,
            I => \N__34751\
        );

    \I__8199\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34748\
        );

    \I__8198\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34745\
        );

    \I__8197\ : CascadeMux
    port map (
            O => \N__34785\,
            I => \N__34742\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__34782\,
            I => \N__34737\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__34779\,
            I => \N__34737\
        );

    \I__8194\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34734\
        );

    \I__8193\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34731\
        );

    \I__8192\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34728\
        );

    \I__8191\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34724\
        );

    \I__8190\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34721\
        );

    \I__8189\ : InMux
    port map (
            O => \N__34761\,
            I => \N__34718\
        );

    \I__8188\ : CascadeMux
    port map (
            O => \N__34760\,
            I => \N__34715\
        );

    \I__8187\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34712\
        );

    \I__8186\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34709\
        );

    \I__8185\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34706\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__34748\,
            I => \N__34703\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__34745\,
            I => \N__34700\
        );

    \I__8182\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34697\
        );

    \I__8181\ : Span4Mux_v
    port map (
            O => \N__34737\,
            I => \N__34690\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__34734\,
            I => \N__34690\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__34731\,
            I => \N__34690\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__34728\,
            I => \N__34687\
        );

    \I__8177\ : CascadeMux
    port map (
            O => \N__34727\,
            I => \N__34684\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__34724\,
            I => \N__34679\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34679\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__34718\,
            I => \N__34676\
        );

    \I__8173\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34673\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34670\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__34709\,
            I => \N__34665\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__34706\,
            I => \N__34665\
        );

    \I__8169\ : Span4Mux_v
    port map (
            O => \N__34703\,
            I => \N__34660\
        );

    \I__8168\ : Span4Mux_s1_v
    port map (
            O => \N__34700\,
            I => \N__34660\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__34697\,
            I => \N__34657\
        );

    \I__8166\ : Span4Mux_v
    port map (
            O => \N__34690\,
            I => \N__34652\
        );

    \I__8165\ : Span4Mux_v
    port map (
            O => \N__34687\,
            I => \N__34652\
        );

    \I__8164\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34649\
        );

    \I__8163\ : Span4Mux_v
    port map (
            O => \N__34679\,
            I => \N__34644\
        );

    \I__8162\ : Span4Mux_v
    port map (
            O => \N__34676\,
            I => \N__34644\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34641\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__34670\,
            I => \N__34634\
        );

    \I__8159\ : Span4Mux_v
    port map (
            O => \N__34665\,
            I => \N__34634\
        );

    \I__8158\ : Span4Mux_v
    port map (
            O => \N__34660\,
            I => \N__34634\
        );

    \I__8157\ : Span4Mux_v
    port map (
            O => \N__34657\,
            I => \N__34631\
        );

    \I__8156\ : Sp12to4
    port map (
            O => \N__34652\,
            I => \N__34628\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34625\
        );

    \I__8154\ : Span4Mux_h
    port map (
            O => \N__34644\,
            I => \N__34622\
        );

    \I__8153\ : Span4Mux_v
    port map (
            O => \N__34641\,
            I => \N__34619\
        );

    \I__8152\ : Sp12to4
    port map (
            O => \N__34634\,
            I => \N__34616\
        );

    \I__8151\ : Sp12to4
    port map (
            O => \N__34631\,
            I => \N__34613\
        );

    \I__8150\ : Span12Mux_h
    port map (
            O => \N__34628\,
            I => \N__34610\
        );

    \I__8149\ : Span4Mux_v
    port map (
            O => \N__34625\,
            I => \N__34603\
        );

    \I__8148\ : Span4Mux_v
    port map (
            O => \N__34622\,
            I => \N__34603\
        );

    \I__8147\ : Span4Mux_v
    port map (
            O => \N__34619\,
            I => \N__34603\
        );

    \I__8146\ : Span12Mux_s9_h
    port map (
            O => \N__34616\,
            I => \N__34600\
        );

    \I__8145\ : Span12Mux_h
    port map (
            O => \N__34613\,
            I => \N__34595\
        );

    \I__8144\ : Span12Mux_v
    port map (
            O => \N__34610\,
            I => \N__34595\
        );

    \I__8143\ : Odrv4
    port map (
            O => \N__34603\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__8142\ : Odrv12
    port map (
            O => \N__34600\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__8141\ : Odrv12
    port map (
            O => \N__34595\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__8140\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34585\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__34585\,
            I => \N__34582\
        );

    \I__8138\ : Span4Mux_h
    port map (
            O => \N__34582\,
            I => \N__34579\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__34579\,
            I => \this_ppu.oam_cache.mem_15\
        );

    \I__8136\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34573\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__8134\ : Span4Mux_h
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__8133\ : Odrv4
    port map (
            O => \N__34567\,
            I => \this_ppu.oam_cache.mem_14\
        );

    \I__8132\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34561\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__34561\,
            I => \N__34555\
        );

    \I__8130\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34547\
        );

    \I__8129\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34547\
        );

    \I__8128\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34547\
        );

    \I__8127\ : Span4Mux_v
    port map (
            O => \N__34555\,
            I => \N__34544\
        );

    \I__8126\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34541\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34538\
        );

    \I__8124\ : Span4Mux_v
    port map (
            O => \N__34544\,
            I => \N__34535\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34532\
        );

    \I__8122\ : Span4Mux_h
    port map (
            O => \N__34538\,
            I => \N__34529\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__34535\,
            I => \N__34526\
        );

    \I__8120\ : Span4Mux_h
    port map (
            O => \N__34532\,
            I => \N__34521\
        );

    \I__8119\ : Span4Mux_v
    port map (
            O => \N__34529\,
            I => \N__34521\
        );

    \I__8118\ : Odrv4
    port map (
            O => \N__34526\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__34521\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__8116\ : InMux
    port map (
            O => \N__34516\,
            I => \N__34513\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__34513\,
            I => \N__34510\
        );

    \I__8114\ : Span4Mux_v
    port map (
            O => \N__34510\,
            I => \N__34507\
        );

    \I__8113\ : Span4Mux_v
    port map (
            O => \N__34507\,
            I => \N__34504\
        );

    \I__8112\ : Odrv4
    port map (
            O => \N__34504\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_22\
        );

    \I__8111\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34496\
        );

    \I__8110\ : CascadeMux
    port map (
            O => \N__34500\,
            I => \N__34492\
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__34499\,
            I => \N__34489\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__34496\,
            I => \N__34485\
        );

    \I__8107\ : InMux
    port map (
            O => \N__34495\,
            I => \N__34475\
        );

    \I__8106\ : InMux
    port map (
            O => \N__34492\,
            I => \N__34475\
        );

    \I__8105\ : InMux
    port map (
            O => \N__34489\,
            I => \N__34475\
        );

    \I__8104\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34475\
        );

    \I__8103\ : Span4Mux_h
    port map (
            O => \N__34485\,
            I => \N__34472\
        );

    \I__8102\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34469\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__34475\,
            I => \N__34466\
        );

    \I__8100\ : Span4Mux_v
    port map (
            O => \N__34472\,
            I => \N__34463\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__34469\,
            I => \N__34460\
        );

    \I__8098\ : Span4Mux_h
    port map (
            O => \N__34466\,
            I => \N__34457\
        );

    \I__8097\ : Span4Mux_v
    port map (
            O => \N__34463\,
            I => \N__34454\
        );

    \I__8096\ : Span4Mux_h
    port map (
            O => \N__34460\,
            I => \N__34449\
        );

    \I__8095\ : Span4Mux_v
    port map (
            O => \N__34457\,
            I => \N__34449\
        );

    \I__8094\ : Odrv4
    port map (
            O => \N__34454\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__8093\ : Odrv4
    port map (
            O => \N__34449\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__8092\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34441\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__34441\,
            I => \N__34438\
        );

    \I__8090\ : Span4Mux_h
    port map (
            O => \N__34438\,
            I => \N__34435\
        );

    \I__8089\ : Span4Mux_v
    port map (
            O => \N__34435\,
            I => \N__34432\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__34432\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_21\
        );

    \I__8087\ : CascadeMux
    port map (
            O => \N__34429\,
            I => \N__34424\
        );

    \I__8086\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34420\
        );

    \I__8085\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34417\
        );

    \I__8084\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34414\
        );

    \I__8083\ : CascadeMux
    port map (
            O => \N__34423\,
            I => \N__34411\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34406\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__34417\,
            I => \N__34406\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__34414\,
            I => \N__34403\
        );

    \I__8079\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34400\
        );

    \I__8078\ : Odrv4
    port map (
            O => \N__34406\,
            I => \this_ppu.un1_M_hoffset_q_9\
        );

    \I__8077\ : Odrv4
    port map (
            O => \N__34403\,
            I => \this_ppu.un1_M_hoffset_q_9\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__34400\,
            I => \this_ppu.un1_M_hoffset_q_9\
        );

    \I__8075\ : InMux
    port map (
            O => \N__34393\,
            I => \N__34387\
        );

    \I__8074\ : InMux
    port map (
            O => \N__34392\,
            I => \N__34387\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34381\
        );

    \I__8072\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34374\
        );

    \I__8071\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34374\
        );

    \I__8070\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34374\
        );

    \I__8069\ : Odrv4
    port map (
            O => \N__34381\,
            I => \this_ppu.un1_M_oam_cache_read_data_c7\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__34374\,
            I => \this_ppu.un1_M_oam_cache_read_data_c7\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__34369\,
            I => \N__34363\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__34368\,
            I => \N__34360\
        );

    \I__8065\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34355\
        );

    \I__8064\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34355\
        );

    \I__8063\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34351\
        );

    \I__8062\ : InMux
    port map (
            O => \N__34360\,
            I => \N__34348\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__34355\,
            I => \N__34345\
        );

    \I__8060\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34339\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__34351\,
            I => \N__34336\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__34348\,
            I => \N__34333\
        );

    \I__8057\ : Span4Mux_h
    port map (
            O => \N__34345\,
            I => \N__34330\
        );

    \I__8056\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34325\
        );

    \I__8055\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34325\
        );

    \I__8054\ : InMux
    port map (
            O => \N__34342\,
            I => \N__34322\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__34339\,
            I => \this_ppu.un1_M_hoffset_q_10\
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__34336\,
            I => \this_ppu.un1_M_hoffset_q_10\
        );

    \I__8051\ : Odrv12
    port map (
            O => \N__34333\,
            I => \this_ppu.un1_M_hoffset_q_10\
        );

    \I__8050\ : Odrv4
    port map (
            O => \N__34330\,
            I => \this_ppu.un1_M_hoffset_q_10\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__34325\,
            I => \this_ppu.un1_M_hoffset_q_10\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__34322\,
            I => \this_ppu.un1_M_hoffset_q_10\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__34309\,
            I => \this_ppu.un1_M_oam_cache_read_data_c7_cascade_\
        );

    \I__8046\ : CascadeMux
    port map (
            O => \N__34306\,
            I => \N__34303\
        );

    \I__8045\ : CascadeBuf
    port map (
            O => \N__34303\,
            I => \N__34297\
        );

    \I__8044\ : CascadeMux
    port map (
            O => \N__34302\,
            I => \N__34293\
        );

    \I__8043\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34290\
        );

    \I__8042\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34287\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__34297\,
            I => \N__34283\
        );

    \I__8040\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34280\
        );

    \I__8039\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34277\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__34290\,
            I => \N__34272\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34272\
        );

    \I__8036\ : InMux
    port map (
            O => \N__34286\,
            I => \N__34269\
        );

    \I__8035\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34266\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34261\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34261\
        );

    \I__8032\ : Span4Mux_v
    port map (
            O => \N__34272\,
            I => \N__34256\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__34269\,
            I => \N__34256\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__34266\,
            I => \N__34253\
        );

    \I__8029\ : Span4Mux_h
    port map (
            O => \N__34261\,
            I => \N__34250\
        );

    \I__8028\ : Span4Mux_h
    port map (
            O => \N__34256\,
            I => \N__34247\
        );

    \I__8027\ : Span12Mux_v
    port map (
            O => \N__34253\,
            I => \N__34244\
        );

    \I__8026\ : Odrv4
    port map (
            O => \N__34250\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__8025\ : Odrv4
    port map (
            O => \N__34247\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__8024\ : Odrv12
    port map (
            O => \N__34244\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__8023\ : CascadeMux
    port map (
            O => \N__34237\,
            I => \N__34234\
        );

    \I__8022\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34231\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__34231\,
            I => \N__34228\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__34228\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNOZ0\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__34225\,
            I => \N__34222\
        );

    \I__8018\ : InMux
    port map (
            O => \N__34222\,
            I => \N__34219\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__34219\,
            I => \N__34216\
        );

    \I__8016\ : Odrv12
    port map (
            O => \N__34216\,
            I => \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNOZ0\
        );

    \I__8015\ : CEMux
    port map (
            O => \N__34213\,
            I => \N__34209\
        );

    \I__8014\ : CEMux
    port map (
            O => \N__34212\,
            I => \N__34206\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__34209\,
            I => \N__34203\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__34206\,
            I => \N__34200\
        );

    \I__8011\ : Span4Mux_h
    port map (
            O => \N__34203\,
            I => \N__34197\
        );

    \I__8010\ : Span12Mux_s10_v
    port map (
            O => \N__34200\,
            I => \N__34194\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__34197\,
            I => \N__34191\
        );

    \I__8008\ : Odrv12
    port map (
            O => \N__34194\,
            I => \this_spr_ram.mem_WE_0\
        );

    \I__8007\ : Odrv4
    port map (
            O => \N__34191\,
            I => \this_spr_ram.mem_WE_0\
        );

    \I__8006\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34183\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34180\
        );

    \I__8004\ : Span4Mux_h
    port map (
            O => \N__34180\,
            I => \N__34177\
        );

    \I__8003\ : Span4Mux_v
    port map (
            O => \N__34177\,
            I => \N__34174\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__34174\,
            I => \this_ppu.oam_cache.mem_7\
        );

    \I__8001\ : InMux
    port map (
            O => \N__34171\,
            I => \N__34168\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__34168\,
            I => \N__34165\
        );

    \I__7999\ : Span4Mux_h
    port map (
            O => \N__34165\,
            I => \N__34162\
        );

    \I__7998\ : Odrv4
    port map (
            O => \N__34162\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_7\
        );

    \I__7997\ : CascadeMux
    port map (
            O => \N__34159\,
            I => \N__34155\
        );

    \I__7996\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34151\
        );

    \I__7995\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34148\
        );

    \I__7994\ : CascadeMux
    port map (
            O => \N__34154\,
            I => \N__34145\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34139\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__34148\,
            I => \N__34139\
        );

    \I__7991\ : InMux
    port map (
            O => \N__34145\,
            I => \N__34136\
        );

    \I__7990\ : CascadeMux
    port map (
            O => \N__34144\,
            I => \N__34131\
        );

    \I__7989\ : Span4Mux_v
    port map (
            O => \N__34139\,
            I => \N__34128\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__34136\,
            I => \N__34125\
        );

    \I__7987\ : InMux
    port map (
            O => \N__34135\,
            I => \N__34121\
        );

    \I__7986\ : InMux
    port map (
            O => \N__34134\,
            I => \N__34118\
        );

    \I__7985\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34115\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__34128\,
            I => \N__34110\
        );

    \I__7983\ : Span4Mux_h
    port map (
            O => \N__34125\,
            I => \N__34110\
        );

    \I__7982\ : InMux
    port map (
            O => \N__34124\,
            I => \N__34107\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__34121\,
            I => \this_ppu.hspr\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__34118\,
            I => \this_ppu.hspr\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__34115\,
            I => \this_ppu.hspr\
        );

    \I__7978\ : Odrv4
    port map (
            O => \N__34110\,
            I => \this_ppu.hspr\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__34107\,
            I => \this_ppu.hspr\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__34096\,
            I => \N__34092\
        );

    \I__7975\ : CascadeMux
    port map (
            O => \N__34095\,
            I => \N__34089\
        );

    \I__7974\ : InMux
    port map (
            O => \N__34092\,
            I => \N__34082\
        );

    \I__7973\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34079\
        );

    \I__7972\ : CascadeMux
    port map (
            O => \N__34088\,
            I => \N__34076\
        );

    \I__7971\ : CascadeMux
    port map (
            O => \N__34087\,
            I => \N__34073\
        );

    \I__7970\ : CascadeMux
    port map (
            O => \N__34086\,
            I => \N__34069\
        );

    \I__7969\ : CascadeMux
    port map (
            O => \N__34085\,
            I => \N__34066\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__34082\,
            I => \N__34059\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__34079\,
            I => \N__34059\
        );

    \I__7966\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34056\
        );

    \I__7965\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34053\
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__34072\,
            I => \N__34050\
        );

    \I__7963\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34047\
        );

    \I__7962\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34044\
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__34065\,
            I => \N__34041\
        );

    \I__7960\ : CascadeMux
    port map (
            O => \N__34064\,
            I => \N__34038\
        );

    \I__7959\ : Span4Mux_v
    port map (
            O => \N__34059\,
            I => \N__34030\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__34056\,
            I => \N__34030\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__34053\,
            I => \N__34030\
        );

    \I__7956\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34027\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__34047\,
            I => \N__34022\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__34044\,
            I => \N__34022\
        );

    \I__7953\ : InMux
    port map (
            O => \N__34041\,
            I => \N__34019\
        );

    \I__7952\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34016\
        );

    \I__7951\ : CascadeMux
    port map (
            O => \N__34037\,
            I => \N__34013\
        );

    \I__7950\ : Span4Mux_v
    port map (
            O => \N__34030\,
            I => \N__34006\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__34006\
        );

    \I__7948\ : Span4Mux_s2_v
    port map (
            O => \N__34022\,
            I => \N__34001\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__34019\,
            I => \N__34001\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__34016\,
            I => \N__33998\
        );

    \I__7945\ : InMux
    port map (
            O => \N__34013\,
            I => \N__33995\
        );

    \I__7944\ : CascadeMux
    port map (
            O => \N__34012\,
            I => \N__33990\
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \N__33985\
        );

    \I__7942\ : Span4Mux_v
    port map (
            O => \N__34006\,
            I => \N__33982\
        );

    \I__7941\ : Span4Mux_v
    port map (
            O => \N__34001\,
            I => \N__33975\
        );

    \I__7940\ : Span4Mux_h
    port map (
            O => \N__33998\,
            I => \N__33975\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__33995\,
            I => \N__33975\
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__33994\,
            I => \N__33972\
        );

    \I__7937\ : CascadeMux
    port map (
            O => \N__33993\,
            I => \N__33969\
        );

    \I__7936\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33966\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__33989\,
            I => \N__33963\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__33988\,
            I => \N__33960\
        );

    \I__7933\ : InMux
    port map (
            O => \N__33985\,
            I => \N__33957\
        );

    \I__7932\ : Span4Mux_h
    port map (
            O => \N__33982\,
            I => \N__33954\
        );

    \I__7931\ : Span4Mux_v
    port map (
            O => \N__33975\,
            I => \N__33951\
        );

    \I__7930\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33948\
        );

    \I__7929\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33945\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__33966\,
            I => \N__33942\
        );

    \I__7927\ : InMux
    port map (
            O => \N__33963\,
            I => \N__33939\
        );

    \I__7926\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33936\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__33957\,
            I => \N__33933\
        );

    \I__7924\ : Span4Mux_h
    port map (
            O => \N__33954\,
            I => \N__33930\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__33951\,
            I => \N__33923\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__33948\,
            I => \N__33923\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__33945\,
            I => \N__33923\
        );

    \I__7920\ : Span4Mux_h
    port map (
            O => \N__33942\,
            I => \N__33918\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__33939\,
            I => \N__33918\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__33936\,
            I => \N__33915\
        );

    \I__7917\ : Span12Mux_h
    port map (
            O => \N__33933\,
            I => \N__33912\
        );

    \I__7916\ : Span4Mux_h
    port map (
            O => \N__33930\,
            I => \N__33903\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__33923\,
            I => \N__33903\
        );

    \I__7914\ : Span4Mux_v
    port map (
            O => \N__33918\,
            I => \N__33903\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__33915\,
            I => \N__33903\
        );

    \I__7912\ : Odrv12
    port map (
            O => \N__33912\,
            I => \M_this_ppu_spr_addr_0\
        );

    \I__7911\ : Odrv4
    port map (
            O => \N__33903\,
            I => \M_this_ppu_spr_addr_0\
        );

    \I__7910\ : InMux
    port map (
            O => \N__33898\,
            I => \N__33895\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__33895\,
            I => \N__33891\
        );

    \I__7908\ : InMux
    port map (
            O => \N__33894\,
            I => \N__33888\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__33891\,
            I => \N__33884\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__33888\,
            I => \N__33881\
        );

    \I__7905\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33878\
        );

    \I__7904\ : Span4Mux_v
    port map (
            O => \N__33884\,
            I => \N__33871\
        );

    \I__7903\ : Span4Mux_h
    port map (
            O => \N__33881\,
            I => \N__33871\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__33878\,
            I => \N__33868\
        );

    \I__7901\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33865\
        );

    \I__7900\ : InMux
    port map (
            O => \N__33876\,
            I => \N__33860\
        );

    \I__7899\ : Span4Mux_h
    port map (
            O => \N__33871\,
            I => \N__33857\
        );

    \I__7898\ : Span4Mux_h
    port map (
            O => \N__33868\,
            I => \N__33854\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__33865\,
            I => \N__33851\
        );

    \I__7896\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33848\
        );

    \I__7895\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33845\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__33860\,
            I => \N__33841\
        );

    \I__7893\ : Span4Mux_h
    port map (
            O => \N__33857\,
            I => \N__33838\
        );

    \I__7892\ : Span4Mux_v
    port map (
            O => \N__33854\,
            I => \N__33833\
        );

    \I__7891\ : Span4Mux_h
    port map (
            O => \N__33851\,
            I => \N__33833\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33830\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__33845\,
            I => \N__33827\
        );

    \I__7888\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33824\
        );

    \I__7887\ : Span12Mux_h
    port map (
            O => \N__33841\,
            I => \N__33821\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__33838\,
            I => \N__33814\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__33833\,
            I => \N__33814\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__33830\,
            I => \N__33814\
        );

    \I__7883\ : Span4Mux_v
    port map (
            O => \N__33827\,
            I => \N__33809\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__33824\,
            I => \N__33809\
        );

    \I__7881\ : Odrv12
    port map (
            O => \N__33821\,
            I => \M_this_spr_ram_write_data_0\
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__33814\,
            I => \M_this_spr_ram_write_data_0\
        );

    \I__7879\ : Odrv4
    port map (
            O => \N__33809\,
            I => \M_this_spr_ram_write_data_0\
        );

    \I__7878\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33799\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__33799\,
            I => \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_2\
        );

    \I__7876\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33793\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__33793\,
            I => \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_3\
        );

    \I__7874\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33786\
        );

    \I__7873\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33783\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__33786\,
            I => \N__33780\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__33783\,
            I => \N__33775\
        );

    \I__7870\ : Span4Mux_v
    port map (
            O => \N__33780\,
            I => \N__33771\
        );

    \I__7869\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33766\
        );

    \I__7868\ : InMux
    port map (
            O => \N__33778\,
            I => \N__33766\
        );

    \I__7867\ : Span4Mux_h
    port map (
            O => \N__33775\,
            I => \N__33763\
        );

    \I__7866\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33760\
        );

    \I__7865\ : Odrv4
    port map (
            O => \N__33771\,
            I => \this_ppu.N_510\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__33766\,
            I => \this_ppu.N_510\
        );

    \I__7863\ : Odrv4
    port map (
            O => \N__33763\,
            I => \this_ppu.N_510\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__33760\,
            I => \this_ppu.N_510\
        );

    \I__7861\ : InMux
    port map (
            O => \N__33751\,
            I => \N__33748\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__33748\,
            I => \N__33742\
        );

    \I__7859\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33739\
        );

    \I__7858\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33734\
        );

    \I__7857\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33734\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__33742\,
            I => \N__33731\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__33739\,
            I => \N__33726\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__33734\,
            I => \N__33726\
        );

    \I__7853\ : Sp12to4
    port map (
            O => \N__33731\,
            I => \N__33721\
        );

    \I__7852\ : Span12Mux_h
    port map (
            O => \N__33726\,
            I => \N__33721\
        );

    \I__7851\ : Span12Mux_v
    port map (
            O => \N__33721\,
            I => \N__33718\
        );

    \I__7850\ : Odrv12
    port map (
            O => \N__33718\,
            I => port_address_in_1
        );

    \I__7849\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33710\
        );

    \I__7848\ : InMux
    port map (
            O => \N__33714\,
            I => \N__33705\
        );

    \I__7847\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33705\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__33710\,
            I => \this_ppu.N_916\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__33705\,
            I => \this_ppu.N_916\
        );

    \I__7844\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33697\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__33697\,
            I => \N__33694\
        );

    \I__7842\ : Span4Mux_v
    port map (
            O => \N__33694\,
            I => \N__33691\
        );

    \I__7841\ : Odrv4
    port map (
            O => \N__33691\,
            I => \N_433\
        );

    \I__7840\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33685\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__33685\,
            I => \N__33682\
        );

    \I__7838\ : Span4Mux_v
    port map (
            O => \N__33682\,
            I => \N__33679\
        );

    \I__7837\ : Span4Mux_h
    port map (
            O => \N__33679\,
            I => \N__33676\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__33676\,
            I => \N_438\
        );

    \I__7835\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33670\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__33670\,
            I => \N__33667\
        );

    \I__7833\ : Odrv12
    port map (
            O => \N__33667\,
            I => \M_this_data_tmp_qZ0Z_12\
        );

    \I__7832\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33661\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__33661\,
            I => \N__33658\
        );

    \I__7830\ : Odrv12
    port map (
            O => \N__33658\,
            I => \M_this_oam_ram_write_data_12\
        );

    \I__7829\ : CascadeMux
    port map (
            O => \N__33655\,
            I => \N__33652\
        );

    \I__7828\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33649\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__33649\,
            I => \N__33646\
        );

    \I__7826\ : Span4Mux_h
    port map (
            O => \N__33646\,
            I => \N__33643\
        );

    \I__7825\ : Odrv4
    port map (
            O => \N__33643\,
            I => \M_this_scroll_qZ0Z_2\
        );

    \I__7824\ : CEMux
    port map (
            O => \N__33640\,
            I => \N__33637\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__33637\,
            I => \N__33634\
        );

    \I__7822\ : Span4Mux_v
    port map (
            O => \N__33634\,
            I => \N__33630\
        );

    \I__7821\ : CEMux
    port map (
            O => \N__33633\,
            I => \N__33627\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__33630\,
            I => \N__33622\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33622\
        );

    \I__7818\ : Sp12to4
    port map (
            O => \N__33622\,
            I => \N__33619\
        );

    \I__7817\ : Odrv12
    port map (
            O => \N__33619\,
            I => \N_1318_0\
        );

    \I__7816\ : InMux
    port map (
            O => \N__33616\,
            I => \N__33613\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__33613\,
            I => \M_this_data_tmp_qZ0Z_0\
        );

    \I__7814\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33604\
        );

    \I__7812\ : Span4Mux_h
    port map (
            O => \N__33604\,
            I => \N__33601\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__33601\,
            I => \M_this_oam_ram_write_data_0\
        );

    \I__7810\ : InMux
    port map (
            O => \N__33598\,
            I => \N__33595\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__33595\,
            I => \M_this_data_tmp_qZ0Z_1\
        );

    \I__7808\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33589\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33586\
        );

    \I__7806\ : Span4Mux_h
    port map (
            O => \N__33586\,
            I => \N__33583\
        );

    \I__7805\ : Odrv4
    port map (
            O => \N__33583\,
            I => \M_this_oam_ram_write_data_1\
        );

    \I__7804\ : InMux
    port map (
            O => \N__33580\,
            I => \N__33577\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__7802\ : Odrv12
    port map (
            O => \N__33574\,
            I => \N_434\
        );

    \I__7801\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33568\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__33568\,
            I => \N__33565\
        );

    \I__7799\ : Odrv4
    port map (
            O => \N__33565\,
            I => \this_spr_ram.mem_out_bus5_3\
        );

    \I__7798\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33559\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__33559\,
            I => \N__33556\
        );

    \I__7796\ : Span4Mux_h
    port map (
            O => \N__33556\,
            I => \N__33553\
        );

    \I__7795\ : Odrv4
    port map (
            O => \N__33553\,
            I => \this_spr_ram.mem_out_bus1_3\
        );

    \I__7794\ : InMux
    port map (
            O => \N__33550\,
            I => \N__33547\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__33547\,
            I => \N__33544\
        );

    \I__7792\ : Span4Mux_h
    port map (
            O => \N__33544\,
            I => \N__33541\
        );

    \I__7791\ : Odrv4
    port map (
            O => \N__33541\,
            I => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__33538\,
            I => \N__33534\
        );

    \I__7789\ : CascadeMux
    port map (
            O => \N__33537\,
            I => \N__33531\
        );

    \I__7788\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33528\
        );

    \I__7787\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33524\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__33528\,
            I => \N__33521\
        );

    \I__7785\ : InMux
    port map (
            O => \N__33527\,
            I => \N__33518\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__33524\,
            I => \this_ppu.M_voffset_qZ0Z_2\
        );

    \I__7783\ : Odrv12
    port map (
            O => \N__33521\,
            I => \this_ppu.M_voffset_qZ0Z_2\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__33518\,
            I => \this_ppu.M_voffset_qZ0Z_2\
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__33511\,
            I => \N__33508\
        );

    \I__7780\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33505\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__33505\,
            I => \this_ppu.M_voffset_q_i_2\
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__33502\,
            I => \N__33499\
        );

    \I__7777\ : CascadeBuf
    port map (
            O => \N__33499\,
            I => \N__33496\
        );

    \I__7776\ : CascadeMux
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__7775\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33490\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__33490\,
            I => \N__33486\
        );

    \I__7773\ : CascadeMux
    port map (
            O => \N__33489\,
            I => \N__33483\
        );

    \I__7772\ : Span4Mux_h
    port map (
            O => \N__33486\,
            I => \N__33480\
        );

    \I__7771\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33477\
        );

    \I__7770\ : Span4Mux_h
    port map (
            O => \N__33480\,
            I => \N__33473\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__33477\,
            I => \N__33470\
        );

    \I__7768\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33467\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__33473\,
            I => \N__33464\
        );

    \I__7766\ : Odrv4
    port map (
            O => \N__33470\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__33467\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__7764\ : Odrv4
    port map (
            O => \N__33464\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__7763\ : CascadeMux
    port map (
            O => \N__33457\,
            I => \N__33454\
        );

    \I__7762\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33451\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__33451\,
            I => \this_ppu.M_this_ppu_map_addr_i_5\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__33448\,
            I => \N__33445\
        );

    \I__7759\ : CascadeBuf
    port map (
            O => \N__33445\,
            I => \N__33442\
        );

    \I__7758\ : CascadeMux
    port map (
            O => \N__33442\,
            I => \N__33439\
        );

    \I__7757\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33435\
        );

    \I__7756\ : CascadeMux
    port map (
            O => \N__33438\,
            I => \N__33432\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__33435\,
            I => \N__33429\
        );

    \I__7754\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33426\
        );

    \I__7753\ : Span12Mux_s8_h
    port map (
            O => \N__33429\,
            I => \N__33422\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33419\
        );

    \I__7751\ : InMux
    port map (
            O => \N__33425\,
            I => \N__33416\
        );

    \I__7750\ : Span12Mux_h
    port map (
            O => \N__33422\,
            I => \N__33413\
        );

    \I__7749\ : Odrv12
    port map (
            O => \N__33419\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__33416\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__7747\ : Odrv12
    port map (
            O => \N__33413\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__7746\ : CascadeMux
    port map (
            O => \N__33406\,
            I => \N__33403\
        );

    \I__7745\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33400\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__33400\,
            I => \this_ppu.M_this_ppu_map_addr_i_6\
        );

    \I__7743\ : CascadeMux
    port map (
            O => \N__33397\,
            I => \N__33394\
        );

    \I__7742\ : CascadeBuf
    port map (
            O => \N__33394\,
            I => \N__33391\
        );

    \I__7741\ : CascadeMux
    port map (
            O => \N__33391\,
            I => \N__33387\
        );

    \I__7740\ : CascadeMux
    port map (
            O => \N__33390\,
            I => \N__33384\
        );

    \I__7739\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33381\
        );

    \I__7738\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33378\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__33381\,
            I => \N__33374\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__33378\,
            I => \N__33371\
        );

    \I__7735\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33368\
        );

    \I__7734\ : Span12Mux_h
    port map (
            O => \N__33374\,
            I => \N__33365\
        );

    \I__7733\ : Odrv4
    port map (
            O => \N__33371\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__33368\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__7731\ : Odrv12
    port map (
            O => \N__33365\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__33358\,
            I => \N__33355\
        );

    \I__7729\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33352\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__33352\,
            I => \this_ppu.M_this_ppu_map_addr_i_7\
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__33349\,
            I => \N__33346\
        );

    \I__7726\ : CascadeBuf
    port map (
            O => \N__33346\,
            I => \N__33342\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__33345\,
            I => \N__33339\
        );

    \I__7724\ : CascadeMux
    port map (
            O => \N__33342\,
            I => \N__33336\
        );

    \I__7723\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33333\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33336\,
            I => \N__33330\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33327\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__33330\,
            I => \N__33323\
        );

    \I__7719\ : Span4Mux_h
    port map (
            O => \N__33327\,
            I => \N__33320\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33317\
        );

    \I__7717\ : Span12Mux_s10_h
    port map (
            O => \N__33323\,
            I => \N__33314\
        );

    \I__7716\ : Odrv4
    port map (
            O => \N__33320\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__33317\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__7714\ : Odrv12
    port map (
            O => \N__33314\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__7713\ : CascadeMux
    port map (
            O => \N__33307\,
            I => \N__33304\
        );

    \I__7712\ : InMux
    port map (
            O => \N__33304\,
            I => \N__33301\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__33301\,
            I => \this_ppu.M_this_ppu_map_addr_i_8\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__33298\,
            I => \N__33295\
        );

    \I__7709\ : CascadeBuf
    port map (
            O => \N__33295\,
            I => \N__33292\
        );

    \I__7708\ : CascadeMux
    port map (
            O => \N__33292\,
            I => \N__33288\
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__33291\,
            I => \N__33285\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33282\
        );

    \I__7705\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33279\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33275\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__33279\,
            I => \N__33272\
        );

    \I__7702\ : InMux
    port map (
            O => \N__33278\,
            I => \N__33269\
        );

    \I__7701\ : Span12Mux_s9_h
    port map (
            O => \N__33275\,
            I => \N__33266\
        );

    \I__7700\ : Odrv12
    port map (
            O => \N__33272\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__33269\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__7698\ : Odrv12
    port map (
            O => \N__33266\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__7697\ : CascadeMux
    port map (
            O => \N__33259\,
            I => \N__33256\
        );

    \I__7696\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33253\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__33253\,
            I => \this_ppu.M_this_ppu_map_addr_i_9\
        );

    \I__7694\ : CascadeMux
    port map (
            O => \N__33250\,
            I => \N__33247\
        );

    \I__7693\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33244\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__33244\,
            I => \N__33240\
        );

    \I__7691\ : InMux
    port map (
            O => \N__33243\,
            I => \N__33237\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__33240\,
            I => \this_ppu.M_voffset_qZ0Z_8\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__33237\,
            I => \this_ppu.M_voffset_qZ0Z_8\
        );

    \I__7688\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33229\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__33229\,
            I => \this_ppu.M_voffset_q_i_8\
        );

    \I__7686\ : InMux
    port map (
            O => \N__33226\,
            I => \this_ppu.un1_M_voffset_q_cry_8\
        );

    \I__7685\ : InMux
    port map (
            O => \N__33223\,
            I => \N__33220\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__33220\,
            I => \N__33217\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__33217\,
            I => \N__33212\
        );

    \I__7682\ : InMux
    port map (
            O => \N__33216\,
            I => \N__33209\
        );

    \I__7681\ : InMux
    port map (
            O => \N__33215\,
            I => \N__33206\
        );

    \I__7680\ : Span4Mux_v
    port map (
            O => \N__33212\,
            I => \N__33203\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__33209\,
            I => \N__33198\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33198\
        );

    \I__7677\ : Span4Mux_v
    port map (
            O => \N__33203\,
            I => \N__33195\
        );

    \I__7676\ : Span4Mux_h
    port map (
            O => \N__33198\,
            I => \N__33192\
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__33195\,
            I => \this_ppu.M_state_d14_1\
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__33192\,
            I => \this_ppu.M_state_d14_1\
        );

    \I__7673\ : CascadeMux
    port map (
            O => \N__33187\,
            I => \N__33184\
        );

    \I__7672\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33181\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__33181\,
            I => \N__33177\
        );

    \I__7670\ : CascadeMux
    port map (
            O => \N__33180\,
            I => \N__33174\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__33177\,
            I => \N__33171\
        );

    \I__7668\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33168\
        );

    \I__7667\ : Odrv4
    port map (
            O => \N__33171\,
            I => \M_this_scroll_qZ0Z_0\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__33168\,
            I => \M_this_scroll_qZ0Z_0\
        );

    \I__7665\ : CascadeMux
    port map (
            O => \N__33163\,
            I => \N__33160\
        );

    \I__7664\ : InMux
    port map (
            O => \N__33160\,
            I => \N__33157\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__33157\,
            I => \M_this_scroll_qZ0Z_1\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__33154\,
            I => \N__33151\
        );

    \I__7661\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33148\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__33148\,
            I => \M_this_scroll_qZ0Z_5\
        );

    \I__7659\ : CascadeMux
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__7658\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33139\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__33139\,
            I => \M_this_scroll_qZ0Z_3\
        );

    \I__7656\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33133\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__33133\,
            I => \M_this_scroll_qZ0Z_4\
        );

    \I__7654\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33127\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__33127\,
            I => \M_this_scroll_qZ0Z_6\
        );

    \I__7652\ : CascadeMux
    port map (
            O => \N__33124\,
            I => \N__33121\
        );

    \I__7651\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33118\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__33118\,
            I => \M_this_scroll_qZ0Z_7\
        );

    \I__7649\ : CascadeMux
    port map (
            O => \N__33115\,
            I => \N__33112\
        );

    \I__7648\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33109\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__33109\,
            I => \this_ppu.M_voffset_q_i_0\
        );

    \I__7646\ : CascadeMux
    port map (
            O => \N__33106\,
            I => \N__33103\
        );

    \I__7645\ : InMux
    port map (
            O => \N__33103\,
            I => \N__33099\
        );

    \I__7644\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33095\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33092\
        );

    \I__7642\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33089\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__33095\,
            I => \this_ppu.M_voffset_qZ0Z_1\
        );

    \I__7640\ : Odrv12
    port map (
            O => \N__33092\,
            I => \this_ppu.M_voffset_qZ0Z_1\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__33089\,
            I => \this_ppu.M_voffset_qZ0Z_1\
        );

    \I__7638\ : CascadeMux
    port map (
            O => \N__33082\,
            I => \N__33079\
        );

    \I__7637\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33076\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__33076\,
            I => \this_ppu.M_voffset_q_i_1\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__33073\,
            I => \N__33070\
        );

    \I__7634\ : CascadeBuf
    port map (
            O => \N__33070\,
            I => \N__33067\
        );

    \I__7633\ : CascadeMux
    port map (
            O => \N__33067\,
            I => \N__33064\
        );

    \I__7632\ : InMux
    port map (
            O => \N__33064\,
            I => \N__33060\
        );

    \I__7631\ : CascadeMux
    port map (
            O => \N__33063\,
            I => \N__33057\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__33060\,
            I => \N__33054\
        );

    \I__7629\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33051\
        );

    \I__7628\ : Span4Mux_v
    port map (
            O => \N__33054\,
            I => \N__33046\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33043\
        );

    \I__7626\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33040\
        );

    \I__7625\ : CascadeMux
    port map (
            O => \N__33049\,
            I => \N__33037\
        );

    \I__7624\ : Span4Mux_h
    port map (
            O => \N__33046\,
            I => \N__33034\
        );

    \I__7623\ : Span4Mux_v
    port map (
            O => \N__33043\,
            I => \N__33029\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__33040\,
            I => \N__33029\
        );

    \I__7621\ : InMux
    port map (
            O => \N__33037\,
            I => \N__33026\
        );

    \I__7620\ : Span4Mux_h
    port map (
            O => \N__33034\,
            I => \N__33023\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__33029\,
            I => \N__33020\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__33026\,
            I => \N__33015\
        );

    \I__7617\ : Span4Mux_h
    port map (
            O => \N__33023\,
            I => \N__33015\
        );

    \I__7616\ : Odrv4
    port map (
            O => \N__33020\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__33015\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__7614\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33007\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__33007\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNOZ0\
        );

    \I__7612\ : CascadeMux
    port map (
            O => \N__33004\,
            I => \N__33001\
        );

    \I__7611\ : CascadeBuf
    port map (
            O => \N__33001\,
            I => \N__32998\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__32998\,
            I => \N__32995\
        );

    \I__7609\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32991\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__32994\,
            I => \N__32986\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32982\
        );

    \I__7606\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32979\
        );

    \I__7605\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32975\
        );

    \I__7604\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32972\
        );

    \I__7603\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32969\
        );

    \I__7602\ : Span4Mux_h
    port map (
            O => \N__32982\,
            I => \N__32966\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__32979\,
            I => \N__32963\
        );

    \I__7600\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32960\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32955\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__32972\,
            I => \N__32955\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__32969\,
            I => \N__32952\
        );

    \I__7596\ : Sp12to4
    port map (
            O => \N__32966\,
            I => \N__32949\
        );

    \I__7595\ : Span4Mux_h
    port map (
            O => \N__32963\,
            I => \N__32946\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32943\
        );

    \I__7593\ : Span4Mux_v
    port map (
            O => \N__32955\,
            I => \N__32940\
        );

    \I__7592\ : Span4Mux_v
    port map (
            O => \N__32952\,
            I => \N__32937\
        );

    \I__7591\ : Span12Mux_v
    port map (
            O => \N__32949\,
            I => \N__32934\
        );

    \I__7590\ : Odrv4
    port map (
            O => \N__32946\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__7589\ : Odrv4
    port map (
            O => \N__32943\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__7588\ : Odrv4
    port map (
            O => \N__32940\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__7587\ : Odrv4
    port map (
            O => \N__32937\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__7586\ : Odrv12
    port map (
            O => \N__32934\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__7584\ : CascadeBuf
    port map (
            O => \N__32920\,
            I => \N__32916\
        );

    \I__7583\ : InMux
    port map (
            O => \N__32919\,
            I => \N__32912\
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__32916\,
            I => \N__32909\
        );

    \I__7581\ : CascadeMux
    port map (
            O => \N__32915\,
            I => \N__32906\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__32912\,
            I => \N__32903\
        );

    \I__7579\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32899\
        );

    \I__7578\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32896\
        );

    \I__7577\ : Span4Mux_v
    port map (
            O => \N__32903\,
            I => \N__32893\
        );

    \I__7576\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32890\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__32899\,
            I => \N__32887\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__32896\,
            I => \N__32884\
        );

    \I__7573\ : Span4Mux_h
    port map (
            O => \N__32893\,
            I => \N__32879\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__32890\,
            I => \N__32879\
        );

    \I__7571\ : Sp12to4
    port map (
            O => \N__32887\,
            I => \N__32876\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__32884\,
            I => \N__32873\
        );

    \I__7569\ : Span4Mux_h
    port map (
            O => \N__32879\,
            I => \N__32870\
        );

    \I__7568\ : Span12Mux_h
    port map (
            O => \N__32876\,
            I => \N__32867\
        );

    \I__7567\ : Odrv4
    port map (
            O => \N__32873\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__7566\ : Odrv4
    port map (
            O => \N__32870\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__7565\ : Odrv12
    port map (
            O => \N__32867\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__7564\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32857\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32853\
        );

    \I__7562\ : CascadeMux
    port map (
            O => \N__32856\,
            I => \N__32850\
        );

    \I__7561\ : Span4Mux_h
    port map (
            O => \N__32853\,
            I => \N__32847\
        );

    \I__7560\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32844\
        );

    \I__7559\ : Odrv4
    port map (
            O => \N__32847\,
            I => \this_ppu.read_data_RNI3DGK1_14\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__32844\,
            I => \this_ppu.read_data_RNI3DGK1_14\
        );

    \I__7557\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32836\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__32836\,
            I => \N__32833\
        );

    \I__7555\ : Odrv4
    port map (
            O => \N__32833\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNOZ0\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__32830\,
            I => \N__32827\
        );

    \I__7553\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32823\
        );

    \I__7552\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32819\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__32823\,
            I => \N__32816\
        );

    \I__7550\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32813\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__32819\,
            I => \N__32806\
        );

    \I__7548\ : Span4Mux_v
    port map (
            O => \N__32816\,
            I => \N__32806\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__32813\,
            I => \N__32806\
        );

    \I__7546\ : Span4Mux_h
    port map (
            O => \N__32806\,
            I => \N__32803\
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__32803\,
            I => \this_ppu.M_hoffset_qZ0Z_8\
        );

    \I__7544\ : InMux
    port map (
            O => \N__32800\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_8\
        );

    \I__7543\ : CascadeMux
    port map (
            O => \N__32797\,
            I => \N__32794\
        );

    \I__7542\ : InMux
    port map (
            O => \N__32794\,
            I => \N__32791\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__32791\,
            I => \N__32788\
        );

    \I__7540\ : Span4Mux_h
    port map (
            O => \N__32788\,
            I => \N__32785\
        );

    \I__7539\ : Odrv4
    port map (
            O => \N__32785\,
            I => \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_CO\
        );

    \I__7538\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32779\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__32779\,
            I => \N__32776\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__32776\,
            I => \N__32773\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__32773\,
            I => \this_ppu.oam_cache.mem_18\
        );

    \I__7534\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32767\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__32767\,
            I => \this_ppu.M_oam_cache_read_data_18\
        );

    \I__7532\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32761\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__32761\,
            I => \this_ppu.un1_oam_data_1_6\
        );

    \I__7530\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32755\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__32755\,
            I => \this_ppu.un1_oam_data_1_8\
        );

    \I__7528\ : InMux
    port map (
            O => \N__32752\,
            I => \N__32749\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__32749\,
            I => \this_ppu.un1_oam_data_1_7\
        );

    \I__7526\ : InMux
    port map (
            O => \N__32746\,
            I => \N__32743\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__32743\,
            I => \this_ppu.un1_oam_data_1_5\
        );

    \I__7524\ : CascadeMux
    port map (
            O => \N__32740\,
            I => \N__32736\
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__32739\,
            I => \N__32733\
        );

    \I__7522\ : InMux
    port map (
            O => \N__32736\,
            I => \N__32730\
        );

    \I__7521\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32727\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__32730\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__32727\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__7518\ : CascadeMux
    port map (
            O => \N__32722\,
            I => \N__32718\
        );

    \I__7517\ : CascadeMux
    port map (
            O => \N__32721\,
            I => \N__32715\
        );

    \I__7516\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32712\
        );

    \I__7515\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32709\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__32712\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__32709\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__7512\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32700\
        );

    \I__7511\ : InMux
    port map (
            O => \N__32703\,
            I => \N__32697\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__32700\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__32697\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__7508\ : InMux
    port map (
            O => \N__32692\,
            I => \bfn_22_19_0_\
        );

    \I__7507\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32686\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__32686\,
            I => \N__32683\
        );

    \I__7505\ : Span4Mux_h
    port map (
            O => \N__32683\,
            I => \N__32680\
        );

    \I__7504\ : Odrv4
    port map (
            O => \N__32680\,
            I => \this_ppu.vspr16_0\
        );

    \I__7503\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32674\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__32674\,
            I => \N__32671\
        );

    \I__7501\ : Span4Mux_h
    port map (
            O => \N__32671\,
            I => \N__32668\
        );

    \I__7500\ : Odrv4
    port map (
            O => \N__32668\,
            I => \this_ppu.un1_M_oam_cache_read_data_ac0_13_i\
        );

    \I__7499\ : CascadeMux
    port map (
            O => \N__32665\,
            I => \N__32662\
        );

    \I__7498\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32659\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__32659\,
            I => \N__32656\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__32656\,
            I => \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNOZ0\
        );

    \I__7495\ : CascadeMux
    port map (
            O => \N__32653\,
            I => \N__32650\
        );

    \I__7494\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32647\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32644\
        );

    \I__7492\ : Odrv12
    port map (
            O => \N__32644\,
            I => \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNOZ0\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__32641\,
            I => \N__32638\
        );

    \I__7490\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32635\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32632\
        );

    \I__7488\ : Odrv4
    port map (
            O => \N__32632\,
            I => \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNOZ0\
        );

    \I__7487\ : CascadeMux
    port map (
            O => \N__32629\,
            I => \N__32622\
        );

    \I__7486\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32617\
        );

    \I__7485\ : InMux
    port map (
            O => \N__32627\,
            I => \N__32617\
        );

    \I__7484\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32614\
        );

    \I__7483\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32609\
        );

    \I__7482\ : InMux
    port map (
            O => \N__32622\,
            I => \N__32609\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__32617\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__32614\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__32609\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__7478\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32598\
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__32601\,
            I => \N__32594\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__32598\,
            I => \N__32591\
        );

    \I__7475\ : CascadeMux
    port map (
            O => \N__32597\,
            I => \N__32587\
        );

    \I__7474\ : InMux
    port map (
            O => \N__32594\,
            I => \N__32583\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__32591\,
            I => \N__32580\
        );

    \I__7472\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32575\
        );

    \I__7471\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32575\
        );

    \I__7470\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32572\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__32583\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__7468\ : Odrv4
    port map (
            O => \N__32580\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__32575\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__32572\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__7465\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32560\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__32560\,
            I => \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0\
        );

    \I__7463\ : CascadeMux
    port map (
            O => \N__32557\,
            I => \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0_cascade_\
        );

    \I__7462\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32551\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__32551\,
            I => \this_ppu.M_this_state_q_srsts_0_i_i_1_0Z0Z_0\
        );

    \I__7460\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32545\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32542\
        );

    \I__7458\ : Odrv4
    port map (
            O => \N__32542\,
            I => \this_ppu.N_416\
        );

    \I__7457\ : CascadeMux
    port map (
            O => \N__32539\,
            I => \N__32535\
        );

    \I__7456\ : CascadeMux
    port map (
            O => \N__32538\,
            I => \N__32532\
        );

    \I__7455\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32529\
        );

    \I__7454\ : InMux
    port map (
            O => \N__32532\,
            I => \N__32526\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__32529\,
            I => \this_ppu.M_hoffset_q_i_0\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__32526\,
            I => \this_ppu.M_hoffset_q_i_0\
        );

    \I__7451\ : CascadeMux
    port map (
            O => \N__32521\,
            I => \N__32517\
        );

    \I__7450\ : CascadeMux
    port map (
            O => \N__32520\,
            I => \N__32514\
        );

    \I__7449\ : InMux
    port map (
            O => \N__32517\,
            I => \N__32511\
        );

    \I__7448\ : InMux
    port map (
            O => \N__32514\,
            I => \N__32508\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__32511\,
            I => \this_ppu.M_hoffset_q_i_1\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__32508\,
            I => \this_ppu.M_hoffset_q_i_1\
        );

    \I__7445\ : CascadeMux
    port map (
            O => \N__32503\,
            I => \N__32499\
        );

    \I__7444\ : CascadeMux
    port map (
            O => \N__32502\,
            I => \N__32496\
        );

    \I__7443\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32493\
        );

    \I__7442\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32490\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__32493\,
            I => \this_ppu.M_hoffset_q_i_2\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__32490\,
            I => \this_ppu.M_hoffset_q_i_2\
        );

    \I__7439\ : CascadeMux
    port map (
            O => \N__32485\,
            I => \N__32482\
        );

    \I__7438\ : InMux
    port map (
            O => \N__32482\,
            I => \N__32478\
        );

    \I__7437\ : CascadeMux
    port map (
            O => \N__32481\,
            I => \N__32475\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__32478\,
            I => \N__32472\
        );

    \I__7435\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32469\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__32472\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__32469\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__7432\ : CascadeMux
    port map (
            O => \N__32464\,
            I => \N__32460\
        );

    \I__7431\ : CascadeMux
    port map (
            O => \N__32463\,
            I => \N__32457\
        );

    \I__7430\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32454\
        );

    \I__7429\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32451\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__32454\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__32451\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__7426\ : CEMux
    port map (
            O => \N__32446\,
            I => \N__32443\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__32443\,
            I => \N__32439\
        );

    \I__7424\ : CEMux
    port map (
            O => \N__32442\,
            I => \N__32434\
        );

    \I__7423\ : Span4Mux_v
    port map (
            O => \N__32439\,
            I => \N__32431\
        );

    \I__7422\ : CEMux
    port map (
            O => \N__32438\,
            I => \N__32428\
        );

    \I__7421\ : CEMux
    port map (
            O => \N__32437\,
            I => \N__32424\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__32434\,
            I => \N__32419\
        );

    \I__7419\ : Span4Mux_h
    port map (
            O => \N__32431\,
            I => \N__32414\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__32428\,
            I => \N__32414\
        );

    \I__7417\ : CEMux
    port map (
            O => \N__32427\,
            I => \N__32411\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__32424\,
            I => \N__32408\
        );

    \I__7415\ : CEMux
    port map (
            O => \N__32423\,
            I => \N__32405\
        );

    \I__7414\ : CEMux
    port map (
            O => \N__32422\,
            I => \N__32402\
        );

    \I__7413\ : Span4Mux_h
    port map (
            O => \N__32419\,
            I => \N__32395\
        );

    \I__7412\ : Span4Mux_v
    port map (
            O => \N__32414\,
            I => \N__32395\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__32411\,
            I => \N__32395\
        );

    \I__7410\ : Span4Mux_v
    port map (
            O => \N__32408\,
            I => \N__32390\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__32405\,
            I => \N__32390\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__32402\,
            I => \N__32387\
        );

    \I__7407\ : Span4Mux_h
    port map (
            O => \N__32395\,
            I => \N__32384\
        );

    \I__7406\ : Span4Mux_h
    port map (
            O => \N__32390\,
            I => \N__32381\
        );

    \I__7405\ : Span4Mux_v
    port map (
            O => \N__32387\,
            I => \N__32378\
        );

    \I__7404\ : Span4Mux_v
    port map (
            O => \N__32384\,
            I => \N__32375\
        );

    \I__7403\ : Span4Mux_v
    port map (
            O => \N__32381\,
            I => \N__32370\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__32378\,
            I => \N__32370\
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__32375\,
            I => \N_1286_0\
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__32370\,
            I => \N_1286_0\
        );

    \I__7399\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32362\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__32362\,
            I => \N__32359\
        );

    \I__7397\ : Span12Mux_h
    port map (
            O => \N__32359\,
            I => \N__32356\
        );

    \I__7396\ : Span12Mux_v
    port map (
            O => \N__32356\,
            I => \N__32353\
        );

    \I__7395\ : Odrv12
    port map (
            O => \N__32353\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__32350\,
            I => \N__32347\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32343\
        );

    \I__7392\ : CascadeMux
    port map (
            O => \N__32346\,
            I => \N__32340\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32337\
        );

    \I__7390\ : InMux
    port map (
            O => \N__32340\,
            I => \N__32334\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__32337\,
            I => \N__32331\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__32334\,
            I => \N__32328\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__32331\,
            I => \N__32325\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__32328\,
            I => \N__32322\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__32325\,
            I => \this_ppu.N_511\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__32322\,
            I => \this_ppu.N_511\
        );

    \I__7383\ : CascadeMux
    port map (
            O => \N__32317\,
            I => \this_ppu.M_this_state_q_srsts_0_i_0_i_1Z0Z_6_cascade_\
        );

    \I__7382\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32311\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__32311\,
            I => \N__32306\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32310\,
            I => \N__32303\
        );

    \I__7379\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32298\
        );

    \I__7378\ : Span4Mux_h
    port map (
            O => \N__32306\,
            I => \N__32295\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__32303\,
            I => \N__32292\
        );

    \I__7376\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32289\
        );

    \I__7375\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32286\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__32298\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7373\ : Odrv4
    port map (
            O => \N__32295\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7372\ : Odrv12
    port map (
            O => \N__32292\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__32289\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__32286\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__7369\ : CascadeMux
    port map (
            O => \N__32275\,
            I => \N__32272\
        );

    \I__7368\ : InMux
    port map (
            O => \N__32272\,
            I => \N__32269\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__32269\,
            I => \N__32263\
        );

    \I__7366\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32257\
        );

    \I__7365\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32252\
        );

    \I__7364\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32252\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__32263\,
            I => \N__32249\
        );

    \I__7362\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32246\
        );

    \I__7361\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32241\
        );

    \I__7360\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32241\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__32257\,
            I => \N__32238\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__32252\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__7357\ : Odrv4
    port map (
            O => \N__32249\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__32246\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__32241\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__7354\ : Odrv4
    port map (
            O => \N__32238\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__7353\ : InMux
    port map (
            O => \N__32227\,
            I => \N__32224\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__32224\,
            I => this_ppu_un20_i_a4_0_a3_0_a2_1_1
        );

    \I__7351\ : InMux
    port map (
            O => \N__32221\,
            I => \N__32218\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__32218\,
            I => \N__32214\
        );

    \I__7349\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32211\
        );

    \I__7348\ : Span12Mux_v
    port map (
            O => \N__32214\,
            I => \N__32208\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__32211\,
            I => \N__32205\
        );

    \I__7346\ : Span12Mux_h
    port map (
            O => \N__32208\,
            I => \N__32202\
        );

    \I__7345\ : Span4Mux_v
    port map (
            O => \N__32205\,
            I => \N__32199\
        );

    \I__7344\ : Odrv12
    port map (
            O => \N__32202\,
            I => port_rw_in
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__32199\,
            I => port_rw_in
        );

    \I__7342\ : CascadeMux
    port map (
            O => \N__32194\,
            I => \N__32190\
        );

    \I__7341\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32186\
        );

    \I__7340\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32180\
        );

    \I__7339\ : CascadeMux
    port map (
            O => \N__32189\,
            I => \N__32177\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__32186\,
            I => \N__32174\
        );

    \I__7337\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32171\
        );

    \I__7336\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32168\
        );

    \I__7335\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32165\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__32180\,
            I => \N__32162\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32159\
        );

    \I__7332\ : Span4Mux_v
    port map (
            O => \N__32174\,
            I => \N__32152\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__32171\,
            I => \N__32152\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32152\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__32165\,
            I => \N__32149\
        );

    \I__7328\ : Span4Mux_v
    port map (
            O => \N__32162\,
            I => \N__32142\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__32159\,
            I => \N__32142\
        );

    \I__7326\ : Span4Mux_h
    port map (
            O => \N__32152\,
            I => \N__32142\
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__32149\,
            I => \this_ppu.N_321_0\
        );

    \I__7324\ : Odrv4
    port map (
            O => \N__32142\,
            I => \this_ppu.N_321_0\
        );

    \I__7323\ : CascadeMux
    port map (
            O => \N__32137\,
            I => \N__32133\
        );

    \I__7322\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32129\
        );

    \I__7321\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32124\
        );

    \I__7320\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32124\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__32129\,
            I => \N__32118\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__32124\,
            I => \N__32115\
        );

    \I__7317\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32112\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__32122\,
            I => \N__32108\
        );

    \I__7315\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32104\
        );

    \I__7314\ : Span4Mux_h
    port map (
            O => \N__32118\,
            I => \N__32097\
        );

    \I__7313\ : Span4Mux_v
    port map (
            O => \N__32115\,
            I => \N__32097\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__32112\,
            I => \N__32097\
        );

    \I__7311\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32094\
        );

    \I__7310\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32089\
        );

    \I__7309\ : InMux
    port map (
            O => \N__32107\,
            I => \N__32089\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__32104\,
            I => \this_ppu.N_328_0\
        );

    \I__7307\ : Odrv4
    port map (
            O => \N__32097\,
            I => \this_ppu.N_328_0\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__32094\,
            I => \this_ppu.N_328_0\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__32089\,
            I => \this_ppu.N_328_0\
        );

    \I__7304\ : InMux
    port map (
            O => \N__32080\,
            I => \this_ppu.un1_M_voffset_d_cry_5\
        );

    \I__7303\ : InMux
    port map (
            O => \N__32077\,
            I => \N__32073\
        );

    \I__7302\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32070\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__32073\,
            I => \this_ppu.M_vaddress_qZ0Z_7\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__32070\,
            I => \this_ppu.M_vaddress_qZ0Z_7\
        );

    \I__7299\ : InMux
    port map (
            O => \N__32065\,
            I => \this_ppu.un1_M_voffset_d_cry_6\
        );

    \I__7298\ : InMux
    port map (
            O => \N__32062\,
            I => \bfn_21_24_0_\
        );

    \I__7297\ : CEMux
    port map (
            O => \N__32059\,
            I => \N__32054\
        );

    \I__7296\ : CEMux
    port map (
            O => \N__32058\,
            I => \N__32051\
        );

    \I__7295\ : CEMux
    port map (
            O => \N__32057\,
            I => \N__32047\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__32054\,
            I => \N__32044\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__32051\,
            I => \N__32041\
        );

    \I__7292\ : CEMux
    port map (
            O => \N__32050\,
            I => \N__32038\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32035\
        );

    \I__7290\ : Span4Mux_h
    port map (
            O => \N__32044\,
            I => \N__32032\
        );

    \I__7289\ : Span4Mux_v
    port map (
            O => \N__32041\,
            I => \N__32029\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__32038\,
            I => \N__32026\
        );

    \I__7287\ : Span4Mux_h
    port map (
            O => \N__32035\,
            I => \N__32023\
        );

    \I__7286\ : Span4Mux_v
    port map (
            O => \N__32032\,
            I => \N__32016\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__32029\,
            I => \N__32016\
        );

    \I__7284\ : Span4Mux_v
    port map (
            O => \N__32026\,
            I => \N__32016\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__32023\,
            I => \this_ppu.N_756_0_0\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__32016\,
            I => \this_ppu.N_756_0_0\
        );

    \I__7281\ : InMux
    port map (
            O => \N__32011\,
            I => \N__32008\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__32008\,
            I => \M_this_data_tmp_qZ0Z_2\
        );

    \I__7279\ : InMux
    port map (
            O => \N__32005\,
            I => \N__32002\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__32002\,
            I => \N__31999\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__31999\,
            I => \N__31996\
        );

    \I__7276\ : Odrv4
    port map (
            O => \N__31996\,
            I => \M_this_oam_ram_write_data_2\
        );

    \I__7275\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31990\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__31990\,
            I => \N__31987\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__31987\,
            I => \N__31984\
        );

    \I__7272\ : Span4Mux_h
    port map (
            O => \N__31984\,
            I => \N__31981\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__31981\,
            I => \M_this_data_tmp_qZ0Z_16\
        );

    \I__7270\ : InMux
    port map (
            O => \N__31978\,
            I => \N__31975\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__31975\,
            I => \N__31972\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__31972\,
            I => \N__31969\
        );

    \I__7267\ : Odrv4
    port map (
            O => \N__31969\,
            I => \M_this_oam_ram_write_data_16\
        );

    \I__7266\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31963\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__31963\,
            I => \M_this_data_tmp_qZ0Z_5\
        );

    \I__7264\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31957\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__31957\,
            I => \N__31954\
        );

    \I__7262\ : Span4Mux_v
    port map (
            O => \N__31954\,
            I => \N__31951\
        );

    \I__7261\ : Odrv4
    port map (
            O => \N__31951\,
            I => \M_this_oam_ram_write_data_5\
        );

    \I__7260\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31945\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__31945\,
            I => \N__31942\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__31942\,
            I => \M_this_data_tmp_qZ0Z_15\
        );

    \I__7257\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31936\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__31936\,
            I => \N__31933\
        );

    \I__7255\ : Odrv12
    port map (
            O => \N__31933\,
            I => \M_this_oam_ram_write_data_15\
        );

    \I__7254\ : InMux
    port map (
            O => \N__31930\,
            I => \N__31927\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__31927\,
            I => \M_this_data_tmp_qZ0Z_19\
        );

    \I__7252\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31921\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__31921\,
            I => \N__31918\
        );

    \I__7250\ : Span4Mux_h
    port map (
            O => \N__31918\,
            I => \N__31915\
        );

    \I__7249\ : Odrv4
    port map (
            O => \N__31915\,
            I => \M_this_oam_ram_write_data_19\
        );

    \I__7248\ : CascadeMux
    port map (
            O => \N__31912\,
            I => \N__31909\
        );

    \I__7247\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31906\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__31906\,
            I => \this_ppu.M_oam_cache_read_data_i_17\
        );

    \I__7245\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31900\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__31900\,
            I => \N__31897\
        );

    \I__7243\ : Span4Mux_h
    port map (
            O => \N__31897\,
            I => \N__31894\
        );

    \I__7242\ : Odrv4
    port map (
            O => \N__31894\,
            I => \this_ppu.oam_cache.mem_17\
        );

    \I__7241\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31888\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__31888\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_17\
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__31885\,
            I => \N__31881\
        );

    \I__7238\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31877\
        );

    \I__7237\ : InMux
    port map (
            O => \N__31881\,
            I => \N__31873\
        );

    \I__7236\ : InMux
    port map (
            O => \N__31880\,
            I => \N__31870\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__31877\,
            I => \N__31867\
        );

    \I__7234\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31864\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__31873\,
            I => \N__31853\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__31870\,
            I => \N__31853\
        );

    \I__7231\ : Span4Mux_h
    port map (
            O => \N__31867\,
            I => \N__31853\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__31864\,
            I => \N__31853\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__31863\,
            I => \N__31850\
        );

    \I__7228\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31847\
        );

    \I__7227\ : Span4Mux_v
    port map (
            O => \N__31853\,
            I => \N__31844\
        );

    \I__7226\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31840\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__31847\,
            I => \N__31837\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__31844\,
            I => \N__31834\
        );

    \I__7223\ : CascadeMux
    port map (
            O => \N__31843\,
            I => \N__31831\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31828\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__31837\,
            I => \N__31823\
        );

    \I__7220\ : Span4Mux_h
    port map (
            O => \N__31834\,
            I => \N__31823\
        );

    \I__7219\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31820\
        );

    \I__7218\ : Span12Mux_s11_h
    port map (
            O => \N__31828\,
            I => \N__31817\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__31823\,
            I => \N__31814\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__31820\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7215\ : Odrv12
    port map (
            O => \N__31817\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7214\ : Odrv4
    port map (
            O => \N__31814\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7213\ : InMux
    port map (
            O => \N__31807\,
            I => \N__31803\
        );

    \I__7212\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31800\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__31803\,
            I => \N__31794\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__31800\,
            I => \N__31794\
        );

    \I__7209\ : InMux
    port map (
            O => \N__31799\,
            I => \N__31791\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__31794\,
            I => \N__31787\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__31791\,
            I => \N__31784\
        );

    \I__7206\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31781\
        );

    \I__7205\ : Sp12to4
    port map (
            O => \N__31787\,
            I => \N__31776\
        );

    \I__7204\ : Span12Mux_s10_v
    port map (
            O => \N__31784\,
            I => \N__31776\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__31781\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7202\ : Odrv12
    port map (
            O => \N__31776\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7201\ : InMux
    port map (
            O => \N__31771\,
            I => \this_ppu.un1_M_voffset_d_cry_0\
        );

    \I__7200\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31759\
        );

    \I__7199\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31759\
        );

    \I__7198\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31759\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__31759\,
            I => \N__31754\
        );

    \I__7196\ : InMux
    port map (
            O => \N__31758\,
            I => \N__31751\
        );

    \I__7195\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31748\
        );

    \I__7194\ : Odrv4
    port map (
            O => \N__31754\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__31751\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__31748\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7191\ : InMux
    port map (
            O => \N__31741\,
            I => \this_ppu.un1_M_voffset_d_cry_1\
        );

    \I__7190\ : CascadeMux
    port map (
            O => \N__31738\,
            I => \N__31735\
        );

    \I__7189\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31731\
        );

    \I__7188\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31728\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31722\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__31728\,
            I => \N__31722\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__31727\,
            I => \N__31719\
        );

    \I__7184\ : Span12Mux_s10_v
    port map (
            O => \N__31722\,
            I => \N__31713\
        );

    \I__7183\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31708\
        );

    \I__7182\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31708\
        );

    \I__7181\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31705\
        );

    \I__7180\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31702\
        );

    \I__7179\ : Span12Mux_v
    port map (
            O => \N__31713\,
            I => \N__31699\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__31708\,
            I => \this_ppu.M_vaddress_qZ0Z_3\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__31705\,
            I => \this_ppu.M_vaddress_qZ0Z_3\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__31702\,
            I => \this_ppu.M_vaddress_qZ0Z_3\
        );

    \I__7175\ : Odrv12
    port map (
            O => \N__31699\,
            I => \this_ppu.M_vaddress_qZ0Z_3\
        );

    \I__7174\ : InMux
    port map (
            O => \N__31690\,
            I => \this_ppu.un1_M_voffset_d_cry_2\
        );

    \I__7173\ : CascadeMux
    port map (
            O => \N__31687\,
            I => \N__31684\
        );

    \I__7172\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31681\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__31681\,
            I => \N__31678\
        );

    \I__7170\ : Span4Mux_h
    port map (
            O => \N__31678\,
            I => \N__31674\
        );

    \I__7169\ : CascadeMux
    port map (
            O => \N__31677\,
            I => \N__31670\
        );

    \I__7168\ : Sp12to4
    port map (
            O => \N__31674\,
            I => \N__31666\
        );

    \I__7167\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31663\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31660\
        );

    \I__7165\ : InMux
    port map (
            O => \N__31669\,
            I => \N__31657\
        );

    \I__7164\ : Span12Mux_v
    port map (
            O => \N__31666\,
            I => \N__31654\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__31663\,
            I => \this_ppu.M_vaddress_qZ0Z_4\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__31660\,
            I => \this_ppu.M_vaddress_qZ0Z_4\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__31657\,
            I => \this_ppu.M_vaddress_qZ0Z_4\
        );

    \I__7160\ : Odrv12
    port map (
            O => \N__31654\,
            I => \this_ppu.M_vaddress_qZ0Z_4\
        );

    \I__7159\ : InMux
    port map (
            O => \N__31645\,
            I => \this_ppu.un1_M_voffset_d_cry_3\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__31642\,
            I => \N__31639\
        );

    \I__7157\ : InMux
    port map (
            O => \N__31639\,
            I => \N__31636\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__31636\,
            I => \N__31633\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__31633\,
            I => \N__31628\
        );

    \I__7154\ : CascadeMux
    port map (
            O => \N__31632\,
            I => \N__31625\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__31631\,
            I => \N__31622\
        );

    \I__7152\ : Sp12to4
    port map (
            O => \N__31628\,
            I => \N__31618\
        );

    \I__7151\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31610\
        );

    \I__7150\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31610\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31610\
        );

    \I__7148\ : Span12Mux_v
    port map (
            O => \N__31618\,
            I => \N__31607\
        );

    \I__7147\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31604\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__31610\,
            I => \this_ppu.M_vaddress_qZ0Z_5\
        );

    \I__7145\ : Odrv12
    port map (
            O => \N__31607\,
            I => \this_ppu.M_vaddress_qZ0Z_5\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__31604\,
            I => \this_ppu.M_vaddress_qZ0Z_5\
        );

    \I__7143\ : InMux
    port map (
            O => \N__31597\,
            I => \this_ppu.un1_M_voffset_d_cry_4\
        );

    \I__7142\ : CascadeMux
    port map (
            O => \N__31594\,
            I => \N__31591\
        );

    \I__7141\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31588\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__31588\,
            I => \N__31585\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__31585\,
            I => \N__31582\
        );

    \I__7138\ : Span4Mux_h
    port map (
            O => \N__31582\,
            I => \N__31578\
        );

    \I__7137\ : CascadeMux
    port map (
            O => \N__31581\,
            I => \N__31573\
        );

    \I__7136\ : Sp12to4
    port map (
            O => \N__31578\,
            I => \N__31570\
        );

    \I__7135\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31565\
        );

    \I__7134\ : InMux
    port map (
            O => \N__31576\,
            I => \N__31565\
        );

    \I__7133\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31562\
        );

    \I__7132\ : Span12Mux_v
    port map (
            O => \N__31570\,
            I => \N__31559\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__31565\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__31562\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__7129\ : Odrv12
    port map (
            O => \N__31559\,
            I => \this_ppu.M_vaddress_qZ0Z_6\
        );

    \I__7128\ : InMux
    port map (
            O => \N__31552\,
            I => \this_ppu.un1_oam_data_1_cry_8\
        );

    \I__7127\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31545\
        );

    \I__7126\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31542\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__31545\,
            I => \N__31539\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__31542\,
            I => \N__31535\
        );

    \I__7123\ : Span4Mux_v
    port map (
            O => \N__31539\,
            I => \N__31532\
        );

    \I__7122\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31529\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__31535\,
            I => \this_ppu.un1_oam_data_1_cry_8_THRU_CO\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__31532\,
            I => \this_ppu.un1_oam_data_1_cry_8_THRU_CO\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__31529\,
            I => \this_ppu.un1_oam_data_1_cry_8_THRU_CO\
        );

    \I__7118\ : CascadeMux
    port map (
            O => \N__31522\,
            I => \N__31519\
        );

    \I__7117\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31516\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__31516\,
            I => \this_ppu.vspr_cry_0_c_inv_RNIFK43\
        );

    \I__7115\ : CascadeMux
    port map (
            O => \N__31513\,
            I => \N__31509\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__31512\,
            I => \N__31506\
        );

    \I__7113\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31500\
        );

    \I__7112\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31497\
        );

    \I__7111\ : CascadeMux
    port map (
            O => \N__31505\,
            I => \N__31494\
        );

    \I__7110\ : CascadeMux
    port map (
            O => \N__31504\,
            I => \N__31490\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__31503\,
            I => \N__31487\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__31500\,
            I => \N__31480\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__31497\,
            I => \N__31480\
        );

    \I__7106\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31477\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__31493\,
            I => \N__31474\
        );

    \I__7104\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31470\
        );

    \I__7103\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31467\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__31486\,
            I => \N__31464\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__31485\,
            I => \N__31461\
        );

    \I__7100\ : Span4Mux_s2_v
    port map (
            O => \N__31480\,
            I => \N__31454\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__31477\,
            I => \N__31454\
        );

    \I__7098\ : InMux
    port map (
            O => \N__31474\,
            I => \N__31451\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__31473\,
            I => \N__31448\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__31470\,
            I => \N__31442\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31442\
        );

    \I__7094\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31439\
        );

    \I__7093\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31436\
        );

    \I__7092\ : CascadeMux
    port map (
            O => \N__31460\,
            I => \N__31433\
        );

    \I__7091\ : CascadeMux
    port map (
            O => \N__31459\,
            I => \N__31430\
        );

    \I__7090\ : Span4Mux_v
    port map (
            O => \N__31454\,
            I => \N__31424\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__31451\,
            I => \N__31424\
        );

    \I__7088\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31421\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__31447\,
            I => \N__31418\
        );

    \I__7086\ : Span4Mux_v
    port map (
            O => \N__31442\,
            I => \N__31410\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31410\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__31436\,
            I => \N__31410\
        );

    \I__7083\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31407\
        );

    \I__7082\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31404\
        );

    \I__7081\ : CascadeMux
    port map (
            O => \N__31429\,
            I => \N__31401\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__31424\,
            I => \N__31395\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__31421\,
            I => \N__31395\
        );

    \I__7078\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31392\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__31417\,
            I => \N__31389\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__31410\,
            I => \N__31381\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__31407\,
            I => \N__31381\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31381\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31378\
        );

    \I__7072\ : CascadeMux
    port map (
            O => \N__31400\,
            I => \N__31375\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__31395\,
            I => \N__31370\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__31392\,
            I => \N__31370\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31367\
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__31388\,
            I => \N__31364\
        );

    \I__7067\ : Sp12to4
    port map (
            O => \N__31381\,
            I => \N__31361\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__31378\,
            I => \N__31358\
        );

    \I__7065\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31355\
        );

    \I__7064\ : Span4Mux_h
    port map (
            O => \N__31370\,
            I => \N__31350\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__31367\,
            I => \N__31350\
        );

    \I__7062\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31347\
        );

    \I__7061\ : Span12Mux_v
    port map (
            O => \N__31361\,
            I => \N__31344\
        );

    \I__7060\ : Span12Mux_s11_h
    port map (
            O => \N__31358\,
            I => \N__31341\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__31355\,
            I => \N__31338\
        );

    \I__7058\ : Span4Mux_v
    port map (
            O => \N__31350\,
            I => \N__31333\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__31347\,
            I => \N__31333\
        );

    \I__7056\ : Span12Mux_h
    port map (
            O => \N__31344\,
            I => \N__31328\
        );

    \I__7055\ : Span12Mux_v
    port map (
            O => \N__31341\,
            I => \N__31328\
        );

    \I__7054\ : Span12Mux_s11_h
    port map (
            O => \N__31338\,
            I => \N__31325\
        );

    \I__7053\ : Span4Mux_h
    port map (
            O => \N__31333\,
            I => \N__31322\
        );

    \I__7052\ : Odrv12
    port map (
            O => \N__31328\,
            I => \M_this_ppu_spr_addr_4\
        );

    \I__7051\ : Odrv12
    port map (
            O => \N__31325\,
            I => \M_this_ppu_spr_addr_4\
        );

    \I__7050\ : Odrv4
    port map (
            O => \N__31322\,
            I => \M_this_ppu_spr_addr_4\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31315\,
            I => \this_ppu.vspr_cry_0\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31312\,
            I => \this_ppu.vspr_cry_1\
        );

    \I__7047\ : CascadeMux
    port map (
            O => \N__31309\,
            I => \N__31305\
        );

    \I__7046\ : CascadeMux
    port map (
            O => \N__31308\,
            I => \N__31302\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31298\
        );

    \I__7044\ : InMux
    port map (
            O => \N__31302\,
            I => \N__31295\
        );

    \I__7043\ : CascadeMux
    port map (
            O => \N__31301\,
            I => \N__31292\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__31298\,
            I => \N__31286\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__31295\,
            I => \N__31286\
        );

    \I__7040\ : InMux
    port map (
            O => \N__31292\,
            I => \N__31283\
        );

    \I__7039\ : CascadeMux
    port map (
            O => \N__31291\,
            I => \N__31280\
        );

    \I__7038\ : Span4Mux_s2_v
    port map (
            O => \N__31286\,
            I => \N__31272\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__31283\,
            I => \N__31272\
        );

    \I__7036\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31269\
        );

    \I__7035\ : CascadeMux
    port map (
            O => \N__31279\,
            I => \N__31266\
        );

    \I__7034\ : CascadeMux
    port map (
            O => \N__31278\,
            I => \N__31262\
        );

    \I__7033\ : CascadeMux
    port map (
            O => \N__31277\,
            I => \N__31259\
        );

    \I__7032\ : Span4Mux_v
    port map (
            O => \N__31272\,
            I => \N__31252\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31252\
        );

    \I__7030\ : InMux
    port map (
            O => \N__31266\,
            I => \N__31249\
        );

    \I__7029\ : CascadeMux
    port map (
            O => \N__31265\,
            I => \N__31246\
        );

    \I__7028\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31242\
        );

    \I__7027\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31239\
        );

    \I__7026\ : CascadeMux
    port map (
            O => \N__31258\,
            I => \N__31236\
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__31257\,
            I => \N__31233\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__31252\,
            I => \N__31226\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31226\
        );

    \I__7022\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31223\
        );

    \I__7021\ : CascadeMux
    port map (
            O => \N__31245\,
            I => \N__31220\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__31242\,
            I => \N__31214\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__31239\,
            I => \N__31214\
        );

    \I__7018\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31211\
        );

    \I__7017\ : InMux
    port map (
            O => \N__31233\,
            I => \N__31208\
        );

    \I__7016\ : CascadeMux
    port map (
            O => \N__31232\,
            I => \N__31205\
        );

    \I__7015\ : CascadeMux
    port map (
            O => \N__31231\,
            I => \N__31202\
        );

    \I__7014\ : Span4Mux_v
    port map (
            O => \N__31226\,
            I => \N__31197\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__31223\,
            I => \N__31197\
        );

    \I__7012\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31194\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__31219\,
            I => \N__31191\
        );

    \I__7010\ : Span4Mux_v
    port map (
            O => \N__31214\,
            I => \N__31183\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__31211\,
            I => \N__31183\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31183\
        );

    \I__7007\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31180\
        );

    \I__7006\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31177\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__31197\,
            I => \N__31172\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31172\
        );

    \I__7003\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31169\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__31190\,
            I => \N__31166\
        );

    \I__7001\ : Span4Mux_v
    port map (
            O => \N__31183\,
            I => \N__31158\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__31180\,
            I => \N__31158\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__31177\,
            I => \N__31158\
        );

    \I__6998\ : Span4Mux_v
    port map (
            O => \N__31172\,
            I => \N__31153\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__31169\,
            I => \N__31153\
        );

    \I__6996\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31150\
        );

    \I__6995\ : CascadeMux
    port map (
            O => \N__31165\,
            I => \N__31147\
        );

    \I__6994\ : Sp12to4
    port map (
            O => \N__31158\,
            I => \N__31144\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__31153\,
            I => \N__31139\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__31150\,
            I => \N__31139\
        );

    \I__6991\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31136\
        );

    \I__6990\ : Span12Mux_v
    port map (
            O => \N__31144\,
            I => \N__31133\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__31139\,
            I => \N__31128\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__31136\,
            I => \N__31128\
        );

    \I__6987\ : Span12Mux_h
    port map (
            O => \N__31133\,
            I => \N__31125\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__31128\,
            I => \N__31122\
        );

    \I__6985\ : Odrv12
    port map (
            O => \N__31125\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__31122\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__6983\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31114\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__31114\,
            I => \this_ppu.M_hoffset_q_i_8\
        );

    \I__6981\ : InMux
    port map (
            O => \N__31111\,
            I => \this_ppu.un1_M_hoffset_q_2_cry_8\
        );

    \I__6980\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31105\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__31105\,
            I => \this_ppu.vspr12_0\
        );

    \I__6978\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31099\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__31099\,
            I => \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNOZ0\
        );

    \I__6976\ : CascadeMux
    port map (
            O => \N__31096\,
            I => \N__31092\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__31095\,
            I => \N__31089\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31083\
        );

    \I__6973\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31080\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__31088\,
            I => \N__31077\
        );

    \I__6971\ : CascadeMux
    port map (
            O => \N__31087\,
            I => \N__31073\
        );

    \I__6970\ : CascadeMux
    port map (
            O => \N__31086\,
            I => \N__31070\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__31083\,
            I => \N__31064\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__31080\,
            I => \N__31064\
        );

    \I__6967\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31061\
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__31076\,
            I => \N__31058\
        );

    \I__6965\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31054\
        );

    \I__6964\ : InMux
    port map (
            O => \N__31070\,
            I => \N__31051\
        );

    \I__6963\ : CascadeMux
    port map (
            O => \N__31069\,
            I => \N__31048\
        );

    \I__6962\ : Span4Mux_s2_v
    port map (
            O => \N__31064\,
            I => \N__31042\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__31061\,
            I => \N__31042\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31058\,
            I => \N__31039\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__31057\,
            I => \N__31036\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__31032\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__31051\,
            I => \N__31029\
        );

    \I__6956\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31026\
        );

    \I__6955\ : CascadeMux
    port map (
            O => \N__31047\,
            I => \N__31023\
        );

    \I__6954\ : Span4Mux_v
    port map (
            O => \N__31042\,
            I => \N__31017\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__31039\,
            I => \N__31017\
        );

    \I__6952\ : InMux
    port map (
            O => \N__31036\,
            I => \N__31014\
        );

    \I__6951\ : CascadeMux
    port map (
            O => \N__31035\,
            I => \N__31011\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__31032\,
            I => \N__31002\
        );

    \I__6949\ : Span4Mux_h
    port map (
            O => \N__31029\,
            I => \N__31002\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__31026\,
            I => \N__31002\
        );

    \I__6947\ : InMux
    port map (
            O => \N__31023\,
            I => \N__30999\
        );

    \I__6946\ : CascadeMux
    port map (
            O => \N__31022\,
            I => \N__30996\
        );

    \I__6945\ : Span4Mux_h
    port map (
            O => \N__31017\,
            I => \N__30990\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__31014\,
            I => \N__30990\
        );

    \I__6943\ : InMux
    port map (
            O => \N__31011\,
            I => \N__30987\
        );

    \I__6942\ : CascadeMux
    port map (
            O => \N__31010\,
            I => \N__30984\
        );

    \I__6941\ : CascadeMux
    port map (
            O => \N__31009\,
            I => \N__30980\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__31002\,
            I => \N__30975\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30975\
        );

    \I__6938\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30972\
        );

    \I__6937\ : CascadeMux
    port map (
            O => \N__30995\,
            I => \N__30969\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__30990\,
            I => \N__30964\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__30987\,
            I => \N__30964\
        );

    \I__6934\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30961\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__30983\,
            I => \N__30958\
        );

    \I__6932\ : InMux
    port map (
            O => \N__30980\,
            I => \N__30955\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__30975\,
            I => \N__30950\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30950\
        );

    \I__6929\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30946\
        );

    \I__6928\ : Span4Mux_h
    port map (
            O => \N__30964\,
            I => \N__30941\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30941\
        );

    \I__6926\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30938\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__30955\,
            I => \N__30935\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__30950\,
            I => \N__30932\
        );

    \I__6923\ : CascadeMux
    port map (
            O => \N__30949\,
            I => \N__30929\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__30946\,
            I => \N__30926\
        );

    \I__6921\ : Span4Mux_v
    port map (
            O => \N__30941\,
            I => \N__30921\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__30938\,
            I => \N__30921\
        );

    \I__6919\ : Span12Mux_h
    port map (
            O => \N__30935\,
            I => \N__30918\
        );

    \I__6918\ : Sp12to4
    port map (
            O => \N__30932\,
            I => \N__30915\
        );

    \I__6917\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30912\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__30926\,
            I => \N__30907\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__30921\,
            I => \N__30907\
        );

    \I__6914\ : Span12Mux_v
    port map (
            O => \N__30918\,
            I => \N__30900\
        );

    \I__6913\ : Span12Mux_h
    port map (
            O => \N__30915\,
            I => \N__30900\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30900\
        );

    \I__6911\ : Odrv4
    port map (
            O => \N__30907\,
            I => \M_this_ppu_spr_addr_1\
        );

    \I__6910\ : Odrv12
    port map (
            O => \N__30900\,
            I => \M_this_ppu_spr_addr_1\
        );

    \I__6909\ : InMux
    port map (
            O => \N__30895\,
            I => \this_ppu.hspr_cry_0\
        );

    \I__6908\ : InMux
    port map (
            O => \N__30892\,
            I => \this_ppu.hspr_cry_1\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__30889\,
            I => \N__30885\
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__30888\,
            I => \N__30882\
        );

    \I__6905\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30876\
        );

    \I__6904\ : InMux
    port map (
            O => \N__30882\,
            I => \N__30873\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__30881\,
            I => \N__30870\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__30880\,
            I => \N__30867\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__30879\,
            I => \N__30863\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__30876\,
            I => \N__30859\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__30873\,
            I => \N__30856\
        );

    \I__6898\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30853\
        );

    \I__6897\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30850\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__30866\,
            I => \N__30847\
        );

    \I__6895\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30844\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__30862\,
            I => \N__30841\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__30859\,
            I => \N__30832\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__30856\,
            I => \N__30832\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__30853\,
            I => \N__30832\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__30850\,
            I => \N__30829\
        );

    \I__6889\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30826\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__30844\,
            I => \N__30823\
        );

    \I__6887\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30820\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__30840\,
            I => \N__30817\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__30839\,
            I => \N__30812\
        );

    \I__6884\ : Span4Mux_v
    port map (
            O => \N__30832\,
            I => \N__30803\
        );

    \I__6883\ : Span4Mux_h
    port map (
            O => \N__30829\,
            I => \N__30803\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__30826\,
            I => \N__30803\
        );

    \I__6881\ : Span4Mux_s0_v
    port map (
            O => \N__30823\,
            I => \N__30797\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30797\
        );

    \I__6879\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30794\
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__30816\,
            I => \N__30791\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__30815\,
            I => \N__30788\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30812\,
            I => \N__30784\
        );

    \I__6875\ : CascadeMux
    port map (
            O => \N__30811\,
            I => \N__30781\
        );

    \I__6874\ : CascadeMux
    port map (
            O => \N__30810\,
            I => \N__30778\
        );

    \I__6873\ : Span4Mux_v
    port map (
            O => \N__30803\,
            I => \N__30775\
        );

    \I__6872\ : CascadeMux
    port map (
            O => \N__30802\,
            I => \N__30772\
        );

    \I__6871\ : Span4Mux_v
    port map (
            O => \N__30797\,
            I => \N__30769\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30766\
        );

    \I__6869\ : InMux
    port map (
            O => \N__30791\,
            I => \N__30763\
        );

    \I__6868\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30760\
        );

    \I__6867\ : CascadeMux
    port map (
            O => \N__30787\,
            I => \N__30757\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__30784\,
            I => \N__30754\
        );

    \I__6865\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30751\
        );

    \I__6864\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30747\
        );

    \I__6863\ : Span4Mux_h
    port map (
            O => \N__30775\,
            I => \N__30744\
        );

    \I__6862\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30741\
        );

    \I__6861\ : Span4Mux_v
    port map (
            O => \N__30769\,
            I => \N__30734\
        );

    \I__6860\ : Span4Mux_h
    port map (
            O => \N__30766\,
            I => \N__30734\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__30763\,
            I => \N__30734\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__30760\,
            I => \N__30731\
        );

    \I__6857\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30728\
        );

    \I__6856\ : Span12Mux_h
    port map (
            O => \N__30754\,
            I => \N__30723\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__30751\,
            I => \N__30723\
        );

    \I__6854\ : CascadeMux
    port map (
            O => \N__30750\,
            I => \N__30720\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__30747\,
            I => \N__30717\
        );

    \I__6852\ : Span4Mux_h
    port map (
            O => \N__30744\,
            I => \N__30714\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__30741\,
            I => \N__30711\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__30734\,
            I => \N__30704\
        );

    \I__6849\ : Span4Mux_h
    port map (
            O => \N__30731\,
            I => \N__30704\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__30728\,
            I => \N__30704\
        );

    \I__6847\ : Span12Mux_h
    port map (
            O => \N__30723\,
            I => \N__30701\
        );

    \I__6846\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30698\
        );

    \I__6845\ : Span12Mux_s11_h
    port map (
            O => \N__30717\,
            I => \N__30695\
        );

    \I__6844\ : Span4Mux_h
    port map (
            O => \N__30714\,
            I => \N__30688\
        );

    \I__6843\ : Span4Mux_v
    port map (
            O => \N__30711\,
            I => \N__30688\
        );

    \I__6842\ : Span4Mux_v
    port map (
            O => \N__30704\,
            I => \N__30688\
        );

    \I__6841\ : Span12Mux_v
    port map (
            O => \N__30701\,
            I => \N__30683\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__30698\,
            I => \N__30683\
        );

    \I__6839\ : Odrv12
    port map (
            O => \N__30695\,
            I => \M_this_ppu_spr_addr_2\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__30688\,
            I => \M_this_ppu_spr_addr_2\
        );

    \I__6837\ : Odrv12
    port map (
            O => \N__30683\,
            I => \M_this_ppu_spr_addr_2\
        );

    \I__6836\ : CascadeMux
    port map (
            O => \N__30676\,
            I => \N__30673\
        );

    \I__6835\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30670\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__30670\,
            I => \this_ppu.M_oam_cache_read_data_i_9\
        );

    \I__6833\ : CascadeMux
    port map (
            O => \N__30667\,
            I => \this_ppu.N_424_cascade_\
        );

    \I__6832\ : InMux
    port map (
            O => \N__30664\,
            I => \N__30661\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__30661\,
            I => \N__30658\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__30658\,
            I => \this_ppu.N_449\
        );

    \I__6829\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30652\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__30652\,
            I => \M_this_state_q_RNI1G0LZ0Z_1\
        );

    \I__6827\ : CascadeMux
    port map (
            O => \N__30649\,
            I => \N__30646\
        );

    \I__6826\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30640\
        );

    \I__6825\ : InMux
    port map (
            O => \N__30645\,
            I => \N__30640\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__30640\,
            I => \N__30637\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__30637\,
            I => \this_ppu.N_341_0\
        );

    \I__6822\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30629\
        );

    \I__6821\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30622\
        );

    \I__6820\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30619\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__30629\,
            I => \N__30616\
        );

    \I__6818\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30611\
        );

    \I__6817\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30611\
        );

    \I__6816\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30608\
        );

    \I__6815\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30605\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__30622\,
            I => \N__30594\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__30619\,
            I => \N__30594\
        );

    \I__6812\ : Span4Mux_h
    port map (
            O => \N__30616\,
            I => \N__30594\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__30611\,
            I => \N__30594\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__30608\,
            I => \N__30594\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__30605\,
            I => \N__30591\
        );

    \I__6808\ : Span4Mux_v
    port map (
            O => \N__30594\,
            I => \N__30588\
        );

    \I__6807\ : Span4Mux_h
    port map (
            O => \N__30591\,
            I => \N__30585\
        );

    \I__6806\ : Span4Mux_h
    port map (
            O => \N__30588\,
            I => \N__30582\
        );

    \I__6805\ : Odrv4
    port map (
            O => \N__30585\,
            I => \this_ppu.N_934\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__30582\,
            I => \this_ppu.N_934\
        );

    \I__6803\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30573\
        );

    \I__6802\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30567\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__30573\,
            I => \N__30564\
        );

    \I__6800\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30561\
        );

    \I__6799\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30556\
        );

    \I__6798\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30556\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__30567\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6796\ : Odrv12
    port map (
            O => \N__30564\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__30561\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__30556\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__6793\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30544\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__30544\,
            I => \N__30540\
        );

    \I__6791\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30535\
        );

    \I__6790\ : Span4Mux_h
    port map (
            O => \N__30540\,
            I => \N__30532\
        );

    \I__6789\ : InMux
    port map (
            O => \N__30539\,
            I => \N__30529\
        );

    \I__6788\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30526\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__30535\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__30532\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__30529\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__30526\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__6783\ : InMux
    port map (
            O => \N__30517\,
            I => \N__30514\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__30514\,
            I => this_ppu_un20_i_a4_0_a2_0_a2_0_2
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__30511\,
            I => \N_311_0_cascade_\
        );

    \I__6780\ : InMux
    port map (
            O => \N__30508\,
            I => \N__30505\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__30505\,
            I => \M_this_state_q_RNI244K2Z0Z_10\
        );

    \I__6778\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30495\
        );

    \I__6777\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30491\
        );

    \I__6776\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30486\
        );

    \I__6775\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30486\
        );

    \I__6774\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30483\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30480\
        );

    \I__6772\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30477\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__30491\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__30486\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__30483\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__30480\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__30477\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__6766\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30463\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__30463\,
            I => \M_this_state_q_RNIR71EZ0Z_10\
        );

    \I__6764\ : CascadeMux
    port map (
            O => \N__30460\,
            I => \N__30457\
        );

    \I__6763\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30454\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__30454\,
            I => \this_ppu.hspr_cry_0_c_inv_RNI1203\
        );

    \I__6761\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30439\
        );

    \I__6760\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30436\
        );

    \I__6759\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30427\
        );

    \I__6758\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30427\
        );

    \I__6757\ : InMux
    port map (
            O => \N__30447\,
            I => \N__30427\
        );

    \I__6756\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30427\
        );

    \I__6755\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30418\
        );

    \I__6754\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30418\
        );

    \I__6753\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30418\
        );

    \I__6752\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30418\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__30439\,
            I => \N__30409\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30406\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__30427\,
            I => \N__30401\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30401\
        );

    \I__6747\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30396\
        );

    \I__6746\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30396\
        );

    \I__6745\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30387\
        );

    \I__6744\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30387\
        );

    \I__6743\ : InMux
    port map (
            O => \N__30413\,
            I => \N__30387\
        );

    \I__6742\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30387\
        );

    \I__6741\ : Odrv12
    port map (
            O => \N__30409\,
            I => \N_332_0\
        );

    \I__6740\ : Odrv4
    port map (
            O => \N__30406\,
            I => \N_332_0\
        );

    \I__6739\ : Odrv4
    port map (
            O => \N__30401\,
            I => \N_332_0\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__30396\,
            I => \N_332_0\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N_332_0\
        );

    \I__6736\ : CascadeMux
    port map (
            O => \N__30376\,
            I => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_7_cascade_\
        );

    \I__6735\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30370\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__30370\,
            I => \this_ppu.N_405\
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__30367\,
            I => \N__30361\
        );

    \I__6732\ : InMux
    port map (
            O => \N__30366\,
            I => \N__30356\
        );

    \I__6731\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30351\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30364\,
            I => \N__30351\
        );

    \I__6729\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30344\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30360\,
            I => \N__30344\
        );

    \I__6727\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30344\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__30356\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30351\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__30344\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__6723\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_13_cascade_\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__30334\,
            I => \N__30331\
        );

    \I__6721\ : InMux
    port map (
            O => \N__30331\,
            I => \N__30326\
        );

    \I__6720\ : InMux
    port map (
            O => \N__30330\,
            I => \N__30323\
        );

    \I__6719\ : InMux
    port map (
            O => \N__30329\,
            I => \N__30320\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__30326\,
            I => \N__30315\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__30323\,
            I => \N__30315\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30320\,
            I => \N__30310\
        );

    \I__6715\ : Span4Mux_h
    port map (
            O => \N__30315\,
            I => \N__30310\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__30310\,
            I => \this_ppu.N_324_0\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__30307\,
            I => \N__30304\
        );

    \I__6712\ : CascadeBuf
    port map (
            O => \N__30304\,
            I => \N__30301\
        );

    \I__6711\ : CascadeMux
    port map (
            O => \N__30301\,
            I => \N__30296\
        );

    \I__6710\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30293\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__30299\,
            I => \N__30290\
        );

    \I__6708\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30287\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30283\
        );

    \I__6706\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30280\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__30287\,
            I => \N__30277\
        );

    \I__6704\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30274\
        );

    \I__6703\ : Span4Mux_h
    port map (
            O => \N__30283\,
            I => \N__30271\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__30280\,
            I => \N__30266\
        );

    \I__6701\ : Span4Mux_h
    port map (
            O => \N__30277\,
            I => \N__30266\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__30274\,
            I => \this_ppu.M_oamidx_qZ0Z_1\
        );

    \I__6699\ : Odrv4
    port map (
            O => \N__30271\,
            I => \this_ppu.M_oamidx_qZ0Z_1\
        );

    \I__6698\ : Odrv4
    port map (
            O => \N__30266\,
            I => \this_ppu.M_oamidx_qZ0Z_1\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__30259\,
            I => \N__30256\
        );

    \I__6696\ : InMux
    port map (
            O => \N__30256\,
            I => \N__30253\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__30253\,
            I => \N__30250\
        );

    \I__6694\ : Odrv12
    port map (
            O => \N__30250\,
            I => \this_ppu.un1_M_oamidx_q_cry_0_THRU_CO\
        );

    \I__6693\ : InMux
    port map (
            O => \N__30247\,
            I => \this_ppu.un1_M_oamidx_q_cry_0\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__30244\,
            I => \N__30241\
        );

    \I__6691\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30238\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__30238\,
            I => \this_ppu.un1_M_oamidx_q_cry_1_THRU_CO\
        );

    \I__6689\ : InMux
    port map (
            O => \N__30235\,
            I => \this_ppu.un1_M_oamidx_q_cry_1\
        );

    \I__6688\ : InMux
    port map (
            O => \N__30232\,
            I => \this_ppu.un1_M_oamidx_q_cry_2\
        );

    \I__6687\ : CascadeMux
    port map (
            O => \N__30229\,
            I => \N__30226\
        );

    \I__6686\ : CascadeBuf
    port map (
            O => \N__30226\,
            I => \N__30223\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__6684\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30214\
        );

    \I__6683\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30211\
        );

    \I__6682\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30206\
        );

    \I__6681\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30206\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__30214\,
            I => \N__30203\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__30211\,
            I => \this_ppu.M_oamidx_qZ1Z_2\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__30206\,
            I => \this_ppu.M_oamidx_qZ1Z_2\
        );

    \I__6677\ : Odrv12
    port map (
            O => \N__30203\,
            I => \this_ppu.M_oamidx_qZ1Z_2\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__6675\ : CascadeBuf
    port map (
            O => \N__30193\,
            I => \N__30190\
        );

    \I__6674\ : CascadeMux
    port map (
            O => \N__30190\,
            I => \N__30187\
        );

    \I__6673\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30184\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__30184\,
            I => \N__30179\
        );

    \I__6671\ : CascadeMux
    port map (
            O => \N__30183\,
            I => \N__30175\
        );

    \I__6670\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30172\
        );

    \I__6669\ : Span4Mux_v
    port map (
            O => \N__30179\,
            I => \N__30169\
        );

    \I__6668\ : InMux
    port map (
            O => \N__30178\,
            I => \N__30165\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30160\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30155\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__30169\,
            I => \N__30155\
        );

    \I__6664\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30152\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__30165\,
            I => \N__30149\
        );

    \I__6662\ : InMux
    port map (
            O => \N__30164\,
            I => \N__30146\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30143\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__30160\,
            I => \N__30138\
        );

    \I__6659\ : Span4Mux_h
    port map (
            O => \N__30155\,
            I => \N__30138\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__30152\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__30149\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__30146\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__30143\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__6654\ : Odrv4
    port map (
            O => \N__30138\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__30127\,
            I => \N__30124\
        );

    \I__6652\ : CascadeBuf
    port map (
            O => \N__30124\,
            I => \N__30121\
        );

    \I__6651\ : CascadeMux
    port map (
            O => \N__30121\,
            I => \N__30116\
        );

    \I__6650\ : CascadeMux
    port map (
            O => \N__30120\,
            I => \N__30113\
        );

    \I__6649\ : CascadeMux
    port map (
            O => \N__30119\,
            I => \N__30110\
        );

    \I__6648\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30107\
        );

    \I__6647\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30102\
        );

    \I__6646\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30102\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__30107\,
            I => \N__30099\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30094\
        );

    \I__6643\ : Span4Mux_h
    port map (
            O => \N__30099\,
            I => \N__30094\
        );

    \I__6642\ : Odrv4
    port map (
            O => \N__30094\,
            I => \this_ppu.M_oamidx_qZ0Z_3\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__30091\,
            I => \N__30088\
        );

    \I__6640\ : CascadeBuf
    port map (
            O => \N__30088\,
            I => \N__30085\
        );

    \I__6639\ : CascadeMux
    port map (
            O => \N__30085\,
            I => \N__30082\
        );

    \I__6638\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30078\
        );

    \I__6637\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30074\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__30078\,
            I => \N__30071\
        );

    \I__6635\ : CascadeMux
    port map (
            O => \N__30077\,
            I => \N__30067\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__30074\,
            I => \N__30063\
        );

    \I__6633\ : Span4Mux_v
    port map (
            O => \N__30071\,
            I => \N__30060\
        );

    \I__6632\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30057\
        );

    \I__6631\ : InMux
    port map (
            O => \N__30067\,
            I => \N__30054\
        );

    \I__6630\ : InMux
    port map (
            O => \N__30066\,
            I => \N__30051\
        );

    \I__6629\ : Span4Mux_v
    port map (
            O => \N__30063\,
            I => \N__30046\
        );

    \I__6628\ : Span4Mux_h
    port map (
            O => \N__30060\,
            I => \N__30046\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__30057\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__30054\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__30051\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__30046\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__6623\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30034\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__6621\ : Span4Mux_h
    port map (
            O => \N__30031\,
            I => \N__30028\
        );

    \I__6620\ : Odrv4
    port map (
            O => \N__30028\,
            I => \this_ppu.M_state_q_srsts_0_a3_0_o2_0_6\
        );

    \I__6619\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30016\
        );

    \I__6618\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30011\
        );

    \I__6617\ : InMux
    port map (
            O => \N__30023\,
            I => \N__30011\
        );

    \I__6616\ : CascadeMux
    port map (
            O => \N__30022\,
            I => \N__30007\
        );

    \I__6615\ : InMux
    port map (
            O => \N__30021\,
            I => \N__30004\
        );

    \I__6614\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30001\
        );

    \I__6613\ : InMux
    port map (
            O => \N__30019\,
            I => \N__29995\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__30016\,
            I => \N__29990\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__30011\,
            I => \N__29990\
        );

    \I__6610\ : InMux
    port map (
            O => \N__30010\,
            I => \N__29987\
        );

    \I__6609\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29984\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__30004\,
            I => \N__29977\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__30001\,
            I => \N__29977\
        );

    \I__6606\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29974\
        );

    \I__6605\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29969\
        );

    \I__6604\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29969\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__29995\,
            I => \N__29965\
        );

    \I__6602\ : Span4Mux_v
    port map (
            O => \N__29990\,
            I => \N__29962\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__29987\,
            I => \N__29957\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__29984\,
            I => \N__29957\
        );

    \I__6599\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29954\
        );

    \I__6598\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29951\
        );

    \I__6597\ : Span4Mux_v
    port map (
            O => \N__29977\,
            I => \N__29944\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__29974\,
            I => \N__29944\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__29969\,
            I => \N__29944\
        );

    \I__6594\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29941\
        );

    \I__6593\ : Span4Mux_v
    port map (
            O => \N__29965\,
            I => \N__29938\
        );

    \I__6592\ : Span4Mux_h
    port map (
            O => \N__29962\,
            I => \N__29931\
        );

    \I__6591\ : Span4Mux_h
    port map (
            O => \N__29957\,
            I => \N__29931\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__29954\,
            I => \N__29931\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__29951\,
            I => \N__29928\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__29944\,
            I => \N__29925\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__29941\,
            I => \N__29922\
        );

    \I__6586\ : Span4Mux_h
    port map (
            O => \N__29938\,
            I => \N__29917\
        );

    \I__6585\ : Span4Mux_v
    port map (
            O => \N__29931\,
            I => \N__29917\
        );

    \I__6584\ : Span4Mux_h
    port map (
            O => \N__29928\,
            I => \N__29914\
        );

    \I__6583\ : Span4Mux_h
    port map (
            O => \N__29925\,
            I => \N__29911\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__29922\,
            I => \N__29906\
        );

    \I__6581\ : Span4Mux_h
    port map (
            O => \N__29917\,
            I => \N__29906\
        );

    \I__6580\ : Span4Mux_v
    port map (
            O => \N__29914\,
            I => \N__29901\
        );

    \I__6579\ : Span4Mux_v
    port map (
            O => \N__29911\,
            I => \N__29901\
        );

    \I__6578\ : Odrv4
    port map (
            O => \N__29906\,
            I => \this_ppu.N_228_0_i_1_0\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__29901\,
            I => \this_ppu.N_228_0_i_1_0\
        );

    \I__6576\ : CascadeMux
    port map (
            O => \N__29896\,
            I => \N__29893\
        );

    \I__6575\ : CascadeBuf
    port map (
            O => \N__29893\,
            I => \N__29889\
        );

    \I__6574\ : InMux
    port map (
            O => \N__29892\,
            I => \N__29886\
        );

    \I__6573\ : CascadeMux
    port map (
            O => \N__29889\,
            I => \N__29881\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__29886\,
            I => \N__29878\
        );

    \I__6571\ : CascadeMux
    port map (
            O => \N__29885\,
            I => \N__29875\
        );

    \I__6570\ : CascadeMux
    port map (
            O => \N__29884\,
            I => \N__29872\
        );

    \I__6569\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29869\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__29878\,
            I => \N__29866\
        );

    \I__6567\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29861\
        );

    \I__6566\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29861\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__29869\,
            I => \N__29858\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__29866\,
            I => \this_ppu.M_oamidx_qZ0Z_0\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__29861\,
            I => \this_ppu.M_oamidx_qZ0Z_0\
        );

    \I__6562\ : Odrv12
    port map (
            O => \N__29858\,
            I => \this_ppu.M_oamidx_qZ0Z_0\
        );

    \I__6561\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29848\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__29848\,
            I => \N__29844\
        );

    \I__6559\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29840\
        );

    \I__6558\ : Span4Mux_h
    port map (
            O => \N__29844\,
            I => \N__29837\
        );

    \I__6557\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29834\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__29840\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__29837\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__29834\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__6553\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29824\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__29824\,
            I => \this_ppu.N_255\
        );

    \I__6551\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29817\
        );

    \I__6550\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29814\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__29817\,
            I => \N__29810\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__29814\,
            I => \N__29807\
        );

    \I__6547\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29804\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__29810\,
            I => \this_ppu.N_756_0\
        );

    \I__6545\ : Odrv4
    port map (
            O => \N__29807\,
            I => \this_ppu.N_756_0\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__29804\,
            I => \this_ppu.N_756_0\
        );

    \I__6543\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29791\
        );

    \I__6542\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29791\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__29791\,
            I => \this_ppu.un1_M_vaddress_q_c2\
        );

    \I__6540\ : InMux
    port map (
            O => \N__29788\,
            I => \N__29779\
        );

    \I__6539\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29779\
        );

    \I__6538\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29779\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__29779\,
            I => \this_ppu.un1_M_vaddress_q_c5\
        );

    \I__6536\ : SRMux
    port map (
            O => \N__29776\,
            I => \N__29773\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__29773\,
            I => \N__29770\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__29770\,
            I => \N__29766\
        );

    \I__6533\ : SRMux
    port map (
            O => \N__29769\,
            I => \N__29763\
        );

    \I__6532\ : Span4Mux_h
    port map (
            O => \N__29766\,
            I => \N__29760\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__29763\,
            I => \N__29757\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__29760\,
            I => \N__29751\
        );

    \I__6529\ : Span4Mux_v
    port map (
            O => \N__29757\,
            I => \N__29751\
        );

    \I__6528\ : SRMux
    port map (
            O => \N__29756\,
            I => \N__29748\
        );

    \I__6527\ : Sp12to4
    port map (
            O => \N__29751\,
            I => \N__29745\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__29748\,
            I => \N__29742\
        );

    \I__6525\ : Odrv12
    port map (
            O => \N__29745\,
            I => \this_ppu.M_last_q_RNIITCPC\
        );

    \I__6524\ : Odrv4
    port map (
            O => \N__29742\,
            I => \this_ppu.M_last_q_RNIITCPC\
        );

    \I__6523\ : InMux
    port map (
            O => \N__29737\,
            I => \this_ppu.un1_M_oam_cache_read_data_2_cry_8\
        );

    \I__6522\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29731\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29726\
        );

    \I__6520\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29723\
        );

    \I__6519\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29720\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__29726\,
            I => \N__29715\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29715\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__29720\,
            I => \N__29712\
        );

    \I__6515\ : Odrv4
    port map (
            O => \N__29715\,
            I => \this_ppu.N_242_0\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__29712\,
            I => \this_ppu.N_242_0\
        );

    \I__6513\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29704\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29701\
        );

    \I__6511\ : Span4Mux_v
    port map (
            O => \N__29701\,
            I => \N__29698\
        );

    \I__6510\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29695\
        );

    \I__6509\ : Odrv4
    port map (
            O => \N__29695\,
            I => \this_ppu.oam_cache.mem_4\
        );

    \I__6508\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29689\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__29689\,
            I => \N__29686\
        );

    \I__6506\ : Odrv12
    port map (
            O => \N__29686\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_4\
        );

    \I__6505\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29679\
        );

    \I__6504\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29676\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__29679\,
            I => \N__29671\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__29676\,
            I => \N__29667\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29664\
        );

    \I__6500\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29661\
        );

    \I__6499\ : Span4Mux_h
    port map (
            O => \N__29671\,
            I => \N__29658\
        );

    \I__6498\ : InMux
    port map (
            O => \N__29670\,
            I => \N__29655\
        );

    \I__6497\ : Span4Mux_v
    port map (
            O => \N__29667\,
            I => \N__29650\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__29664\,
            I => \N__29650\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__29661\,
            I => \this_ppu.M_hoffset_d_0_sqmuxa_7\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__29658\,
            I => \this_ppu.M_hoffset_d_0_sqmuxa_7\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__29655\,
            I => \this_ppu.M_hoffset_d_0_sqmuxa_7\
        );

    \I__6492\ : Odrv4
    port map (
            O => \N__29650\,
            I => \this_ppu.M_hoffset_d_0_sqmuxa_7\
        );

    \I__6491\ : InMux
    port map (
            O => \N__29641\,
            I => \N__29637\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29634\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__29637\,
            I => \N__29629\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29626\
        );

    \I__6487\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29622\
        );

    \I__6486\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29619\
        );

    \I__6485\ : Span4Mux_h
    port map (
            O => \N__29629\,
            I => \N__29614\
        );

    \I__6484\ : Span4Mux_v
    port map (
            O => \N__29626\,
            I => \N__29614\
        );

    \I__6483\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29611\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__29622\,
            I => \N__29608\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__29619\,
            I => \N__29605\
        );

    \I__6480\ : Span4Mux_v
    port map (
            O => \N__29614\,
            I => \N__29602\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__29611\,
            I => \N__29599\
        );

    \I__6478\ : Span12Mux_v
    port map (
            O => \N__29608\,
            I => \N__29596\
        );

    \I__6477\ : Sp12to4
    port map (
            O => \N__29605\,
            I => \N__29593\
        );

    \I__6476\ : Span4Mux_v
    port map (
            O => \N__29602\,
            I => \N__29588\
        );

    \I__6475\ : Span4Mux_v
    port map (
            O => \N__29599\,
            I => \N__29588\
        );

    \I__6474\ : Odrv12
    port map (
            O => \N__29596\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__6473\ : Odrv12
    port map (
            O => \N__29593\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__29588\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__6471\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29576\
        );

    \I__6470\ : InMux
    port map (
            O => \N__29580\,
            I => \N__29573\
        );

    \I__6469\ : InMux
    port map (
            O => \N__29579\,
            I => \N__29570\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__29576\,
            I => \N__29567\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__29573\,
            I => \N__29564\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29561\
        );

    \I__6465\ : Span12Mux_h
    port map (
            O => \N__29567\,
            I => \N__29557\
        );

    \I__6464\ : Span12Mux_v
    port map (
            O => \N__29564\,
            I => \N__29553\
        );

    \I__6463\ : Span4Mux_h
    port map (
            O => \N__29561\,
            I => \N__29550\
        );

    \I__6462\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29547\
        );

    \I__6461\ : Span12Mux_v
    port map (
            O => \N__29557\,
            I => \N__29544\
        );

    \I__6460\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29541\
        );

    \I__6459\ : Odrv12
    port map (
            O => \N__29553\,
            I => \this_ppu.N_772_0\
        );

    \I__6458\ : Odrv4
    port map (
            O => \N__29550\,
            I => \this_ppu.N_772_0\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__29547\,
            I => \this_ppu.N_772_0\
        );

    \I__6456\ : Odrv12
    port map (
            O => \N__29544\,
            I => \this_ppu.N_772_0\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__29541\,
            I => \this_ppu.N_772_0\
        );

    \I__6454\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29527\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__29527\,
            I => \N__29524\
        );

    \I__6452\ : Odrv12
    port map (
            O => \N__29524\,
            I => \this_ppu.N_760_0\
        );

    \I__6451\ : InMux
    port map (
            O => \N__29521\,
            I => \N__29515\
        );

    \I__6450\ : InMux
    port map (
            O => \N__29520\,
            I => \N__29511\
        );

    \I__6449\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29506\
        );

    \I__6448\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29506\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__29515\,
            I => \N__29503\
        );

    \I__6446\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29500\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__29511\,
            I => \N__29497\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29494\
        );

    \I__6443\ : Span4Mux_v
    port map (
            O => \N__29503\,
            I => \N__29489\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__29500\,
            I => \N__29489\
        );

    \I__6441\ : Span4Mux_v
    port map (
            O => \N__29497\,
            I => \N__29486\
        );

    \I__6440\ : Odrv12
    port map (
            O => \N__29494\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__29489\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__29486\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__29479\,
            I => \this_ppu.N_799_cascade_\
        );

    \I__6436\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29471\
        );

    \I__6435\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29468\
        );

    \I__6434\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29465\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__29471\,
            I => \N__29462\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29468\,
            I => \this_ppu.N_779_0\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__29465\,
            I => \this_ppu.N_779_0\
        );

    \I__6430\ : Odrv4
    port map (
            O => \N__29462\,
            I => \this_ppu.N_779_0\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__29455\,
            I => \N__29452\
        );

    \I__6428\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29444\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__29451\,
            I => \N__29440\
        );

    \I__6426\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29437\
        );

    \I__6425\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29433\
        );

    \I__6424\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29430\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__29447\,
            I => \N__29427\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__29444\,
            I => \N__29424\
        );

    \I__6421\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29419\
        );

    \I__6420\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29419\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29416\
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__29436\,
            I => \N__29412\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__29433\,
            I => \N__29407\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__29430\,
            I => \N__29407\
        );

    \I__6415\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29404\
        );

    \I__6414\ : Span4Mux_v
    port map (
            O => \N__29424\,
            I => \N__29399\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__29419\,
            I => \N__29399\
        );

    \I__6412\ : Span4Mux_v
    port map (
            O => \N__29416\,
            I => \N__29396\
        );

    \I__6411\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29393\
        );

    \I__6410\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29390\
        );

    \I__6409\ : Span4Mux_v
    port map (
            O => \N__29407\,
            I => \N__29385\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__29404\,
            I => \N__29385\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__29399\,
            I => \N__29380\
        );

    \I__6406\ : Span4Mux_h
    port map (
            O => \N__29396\,
            I => \N__29380\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__29393\,
            I => \N__29377\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__29390\,
            I => \N__29374\
        );

    \I__6403\ : Span4Mux_h
    port map (
            O => \N__29385\,
            I => \N__29371\
        );

    \I__6402\ : Odrv4
    port map (
            O => \N__29380\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__29377\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__6400\ : Odrv4
    port map (
            O => \N__29374\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__6399\ : Odrv4
    port map (
            O => \N__29371\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__6398\ : InMux
    port map (
            O => \N__29362\,
            I => \N__29359\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__29359\,
            I => \this_ppu.N_267\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__29356\,
            I => \N__29353\
        );

    \I__6395\ : InMux
    port map (
            O => \N__29353\,
            I => \N__29349\
        );

    \I__6394\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29346\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__29349\,
            I => \N__29342\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29339\
        );

    \I__6391\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29334\
        );

    \I__6390\ : Span4Mux_h
    port map (
            O => \N__29342\,
            I => \N__29331\
        );

    \I__6389\ : Span4Mux_v
    port map (
            O => \N__29339\,
            I => \N__29327\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__29338\,
            I => \N__29324\
        );

    \I__6387\ : CascadeMux
    port map (
            O => \N__29337\,
            I => \N__29320\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__29334\,
            I => \N__29316\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__29331\,
            I => \N__29313\
        );

    \I__6384\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29310\
        );

    \I__6383\ : Span4Mux_h
    port map (
            O => \N__29327\,
            I => \N__29307\
        );

    \I__6382\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29300\
        );

    \I__6381\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29300\
        );

    \I__6380\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29300\
        );

    \I__6379\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29297\
        );

    \I__6378\ : Span12Mux_h
    port map (
            O => \N__29316\,
            I => \N__29294\
        );

    \I__6377\ : Span4Mux_h
    port map (
            O => \N__29313\,
            I => \N__29289\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__29310\,
            I => \N__29289\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__29307\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__29300\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__29297\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__6372\ : Odrv12
    port map (
            O => \N__29294\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__6371\ : Odrv4
    port map (
            O => \N__29289\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__29278\,
            I => \N__29275\
        );

    \I__6369\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29272\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__29272\,
            I => \N__29268\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__29271\,
            I => \N__29265\
        );

    \I__6366\ : Span4Mux_h
    port map (
            O => \N__29268\,
            I => \N__29262\
        );

    \I__6365\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29259\
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__29262\,
            I => \M_this_scroll_qZ0Z_8\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__29259\,
            I => \M_this_scroll_qZ0Z_8\
        );

    \I__6362\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29251\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__29251\,
            I => \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_12\
        );

    \I__6360\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29245\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__29245\,
            I => dma_axb3
        );

    \I__6358\ : CascadeMux
    port map (
            O => \N__29242\,
            I => \this_ppu_un20_i_a4_0_a3_0_a2_3_0_cascade_\
        );

    \I__6357\ : IoInMux
    port map (
            O => \N__29239\,
            I => \N__29236\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__29236\,
            I => \N__29233\
        );

    \I__6355\ : IoSpan4Mux
    port map (
            O => \N__29233\,
            I => \N__29230\
        );

    \I__6354\ : Span4Mux_s2_h
    port map (
            O => \N__29230\,
            I => \N__29226\
        );

    \I__6353\ : InMux
    port map (
            O => \N__29229\,
            I => \N__29220\
        );

    \I__6352\ : Span4Mux_h
    port map (
            O => \N__29226\,
            I => \N__29217\
        );

    \I__6351\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29214\
        );

    \I__6350\ : CascadeMux
    port map (
            O => \N__29224\,
            I => \N__29211\
        );

    \I__6349\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29208\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__29220\,
            I => \N__29205\
        );

    \I__6347\ : Span4Mux_h
    port map (
            O => \N__29217\,
            I => \N__29200\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29200\
        );

    \I__6345\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29197\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29194\
        );

    \I__6343\ : Span4Mux_v
    port map (
            O => \N__29205\,
            I => \N__29191\
        );

    \I__6342\ : Span4Mux_v
    port map (
            O => \N__29200\,
            I => \N__29186\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29186\
        );

    \I__6340\ : Span4Mux_v
    port map (
            O => \N__29194\,
            I => \N__29183\
        );

    \I__6339\ : Span4Mux_h
    port map (
            O => \N__29191\,
            I => \N__29180\
        );

    \I__6338\ : Span4Mux_h
    port map (
            O => \N__29186\,
            I => \N__29177\
        );

    \I__6337\ : Sp12to4
    port map (
            O => \N__29183\,
            I => \N__29174\
        );

    \I__6336\ : Span4Mux_h
    port map (
            O => \N__29180\,
            I => \N__29169\
        );

    \I__6335\ : Span4Mux_v
    port map (
            O => \N__29177\,
            I => \N__29169\
        );

    \I__6334\ : Span12Mux_s9_h
    port map (
            O => \N__29174\,
            I => \N__29166\
        );

    \I__6333\ : Span4Mux_h
    port map (
            O => \N__29169\,
            I => \N__29163\
        );

    \I__6332\ : Odrv12
    port map (
            O => \N__29166\,
            I => dma_0
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__29163\,
            I => dma_0
        );

    \I__6330\ : InMux
    port map (
            O => \N__29158\,
            I => \N__29155\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__29155\,
            I => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_10\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__29152\,
            I => \this_ppu.N_414_1_cascade_\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__29149\,
            I => \N__29145\
        );

    \I__6326\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29142\
        );

    \I__6325\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29136\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__29142\,
            I => \N__29133\
        );

    \I__6323\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29130\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__29140\,
            I => \N__29127\
        );

    \I__6321\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29124\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29121\
        );

    \I__6319\ : Span4Mux_v
    port map (
            O => \N__29133\,
            I => \N__29116\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__29130\,
            I => \N__29116\
        );

    \I__6317\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29112\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__29124\,
            I => \N__29109\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__29121\,
            I => \N__29106\
        );

    \I__6314\ : Span4Mux_v
    port map (
            O => \N__29116\,
            I => \N__29103\
        );

    \I__6313\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29100\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__29112\,
            I => \N__29095\
        );

    \I__6311\ : Span12Mux_v
    port map (
            O => \N__29109\,
            I => \N__29095\
        );

    \I__6310\ : Span4Mux_h
    port map (
            O => \N__29106\,
            I => \N__29090\
        );

    \I__6309\ : Span4Mux_h
    port map (
            O => \N__29103\,
            I => \N__29090\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__29100\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__6307\ : Odrv12
    port map (
            O => \N__29095\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__29090\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__6305\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29080\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29077\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__29077\,
            I => \M_this_data_tmp_qZ0Z_9\
        );

    \I__6302\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29071\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29068\
        );

    \I__6300\ : Odrv12
    port map (
            O => \N__29068\,
            I => \M_this_oam_ram_write_data_9\
        );

    \I__6299\ : CEMux
    port map (
            O => \N__29065\,
            I => \N__29061\
        );

    \I__6298\ : CEMux
    port map (
            O => \N__29064\,
            I => \N__29058\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__29061\,
            I => \N__29054\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__29058\,
            I => \N__29050\
        );

    \I__6295\ : CEMux
    port map (
            O => \N__29057\,
            I => \N__29047\
        );

    \I__6294\ : Span4Mux_h
    port map (
            O => \N__29054\,
            I => \N__29043\
        );

    \I__6293\ : CEMux
    port map (
            O => \N__29053\,
            I => \N__29040\
        );

    \I__6292\ : Span4Mux_v
    port map (
            O => \N__29050\,
            I => \N__29036\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__29047\,
            I => \N__29033\
        );

    \I__6290\ : CEMux
    port map (
            O => \N__29046\,
            I => \N__29030\
        );

    \I__6289\ : Span4Mux_h
    port map (
            O => \N__29043\,
            I => \N__29025\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__29040\,
            I => \N__29025\
        );

    \I__6287\ : CEMux
    port map (
            O => \N__29039\,
            I => \N__29022\
        );

    \I__6286\ : Span4Mux_h
    port map (
            O => \N__29036\,
            I => \N__29015\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__29033\,
            I => \N__29015\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__29030\,
            I => \N__29015\
        );

    \I__6283\ : Span4Mux_v
    port map (
            O => \N__29025\,
            I => \N__29010\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__29010\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__29015\,
            I => \N_1294_0\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__29010\,
            I => \N_1294_0\
        );

    \I__6279\ : InMux
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__6277\ : Odrv12
    port map (
            O => \N__28999\,
            I => \M_this_data_tmp_qZ0Z_14\
        );

    \I__6276\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__6274\ : Span4Mux_v
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__6273\ : Span4Mux_h
    port map (
            O => \N__28987\,
            I => \N__28984\
        );

    \I__6272\ : Odrv4
    port map (
            O => \N__28984\,
            I => \M_this_oam_ram_write_data_14\
        );

    \I__6271\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28978\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__28978\,
            I => \N__28975\
        );

    \I__6269\ : Span12Mux_v
    port map (
            O => \N__28975\,
            I => \N__28972\
        );

    \I__6268\ : Odrv12
    port map (
            O => \N__28972\,
            I => \this_ppu.oam_cache.mem_6\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28966\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__28966\,
            I => \N__28963\
        );

    \I__6265\ : Odrv12
    port map (
            O => \N__28963\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_6\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__28960\,
            I => \this_ppu.un20_i_a4_0_a3_0_a2_1Z0Z_3_cascade_\
        );

    \I__6263\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28951\
        );

    \I__6262\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28951\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28944\
        );

    \I__6260\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28941\
        );

    \I__6259\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28938\
        );

    \I__6258\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28933\
        );

    \I__6257\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28933\
        );

    \I__6256\ : Span4Mux_h
    port map (
            O => \N__28944\,
            I => \N__28930\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__28941\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__28938\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__28933\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__28930\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__28921\,
            I => \N__28917\
        );

    \I__6250\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28914\
        );

    \I__6249\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28911\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__28914\,
            I => \N_260\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N_260\
        );

    \I__6246\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28903\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__28903\,
            I => \this_ppu.N_406\
        );

    \I__6244\ : SRMux
    port map (
            O => \N__28900\,
            I => \N__28867\
        );

    \I__6243\ : SRMux
    port map (
            O => \N__28899\,
            I => \N__28867\
        );

    \I__6242\ : SRMux
    port map (
            O => \N__28898\,
            I => \N__28867\
        );

    \I__6241\ : SRMux
    port map (
            O => \N__28897\,
            I => \N__28867\
        );

    \I__6240\ : SRMux
    port map (
            O => \N__28896\,
            I => \N__28867\
        );

    \I__6239\ : SRMux
    port map (
            O => \N__28895\,
            I => \N__28867\
        );

    \I__6238\ : SRMux
    port map (
            O => \N__28894\,
            I => \N__28867\
        );

    \I__6237\ : SRMux
    port map (
            O => \N__28893\,
            I => \N__28867\
        );

    \I__6236\ : SRMux
    port map (
            O => \N__28892\,
            I => \N__28867\
        );

    \I__6235\ : SRMux
    port map (
            O => \N__28891\,
            I => \N__28867\
        );

    \I__6234\ : SRMux
    port map (
            O => \N__28890\,
            I => \N__28867\
        );

    \I__6233\ : GlobalMux
    port map (
            O => \N__28867\,
            I => \N__28864\
        );

    \I__6232\ : gio2CtrlBuf
    port map (
            O => \N__28864\,
            I => \N_504_g\
        );

    \I__6231\ : CascadeMux
    port map (
            O => \N__28861\,
            I => \N__28858\
        );

    \I__6230\ : CascadeBuf
    port map (
            O => \N__28858\,
            I => \N__28855\
        );

    \I__6229\ : CascadeMux
    port map (
            O => \N__28855\,
            I => \N__28852\
        );

    \I__6228\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28849\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__6226\ : Odrv12
    port map (
            O => \N__28846\,
            I => \this_ppu.N_17_0\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__28843\,
            I => \this_ppu.N_329_0_cascade_\
        );

    \I__6224\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28836\
        );

    \I__6223\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28833\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__28836\,
            I => \this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__28833\,
            I => \this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__28828\,
            I => \N__28825\
        );

    \I__6219\ : CascadeBuf
    port map (
            O => \N__28825\,
            I => \N__28822\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__28822\,
            I => \N__28819\
        );

    \I__6217\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28816\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28813\
        );

    \I__6215\ : Span4Mux_h
    port map (
            O => \N__28813\,
            I => \N__28810\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__28810\,
            I => \this_ppu.N_21_0\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28807\,
            I => \N__28801\
        );

    \I__6212\ : InMux
    port map (
            O => \N__28806\,
            I => \N__28798\
        );

    \I__6211\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28795\
        );

    \I__6210\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28792\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__28801\,
            I => \this_ppu.un1_M_oamcurr_q_2_c3\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__28798\,
            I => \this_ppu.un1_M_oamcurr_q_2_c3\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__28795\,
            I => \this_ppu.un1_M_oamcurr_q_2_c3\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__28792\,
            I => \this_ppu.un1_M_oamcurr_q_2_c3\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__28783\,
            I => \N__28780\
        );

    \I__6204\ : CascadeBuf
    port map (
            O => \N__28780\,
            I => \N__28777\
        );

    \I__6203\ : CascadeMux
    port map (
            O => \N__28777\,
            I => \N__28774\
        );

    \I__6202\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28771\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__28771\,
            I => \N__28768\
        );

    \I__6200\ : Odrv12
    port map (
            O => \N__28768\,
            I => \this_ppu.N_23_0\
        );

    \I__6199\ : InMux
    port map (
            O => \N__28765\,
            I => \N__28756\
        );

    \I__6198\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28756\
        );

    \I__6197\ : InMux
    port map (
            O => \N__28763\,
            I => \N__28756\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__28756\,
            I => \this_ppu.N_329_0\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__28753\,
            I => \N__28750\
        );

    \I__6194\ : CascadeBuf
    port map (
            O => \N__28750\,
            I => \N__28747\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__28747\,
            I => \N__28744\
        );

    \I__6192\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28741\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__28741\,
            I => \N__28737\
        );

    \I__6190\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28730\
        );

    \I__6189\ : Span4Mux_h
    port map (
            O => \N__28737\,
            I => \N__28724\
        );

    \I__6188\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28719\
        );

    \I__6187\ : InMux
    port map (
            O => \N__28735\,
            I => \N__28719\
        );

    \I__6186\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28714\
        );

    \I__6185\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28714\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__28730\,
            I => \N__28711\
        );

    \I__6183\ : InMux
    port map (
            O => \N__28729\,
            I => \N__28706\
        );

    \I__6182\ : InMux
    port map (
            O => \N__28728\,
            I => \N__28706\
        );

    \I__6181\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28703\
        );

    \I__6180\ : Span4Mux_v
    port map (
            O => \N__28724\,
            I => \N__28700\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__28719\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__28714\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__28711\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__28706\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__28703\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__28700\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__28687\,
            I => \N__28684\
        );

    \I__6172\ : CascadeBuf
    port map (
            O => \N__28684\,
            I => \N__28681\
        );

    \I__6171\ : CascadeMux
    port map (
            O => \N__28681\,
            I => \N__28678\
        );

    \I__6170\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28675\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__28675\,
            I => \N__28669\
        );

    \I__6168\ : CascadeMux
    port map (
            O => \N__28674\,
            I => \N__28666\
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__28673\,
            I => \N__28663\
        );

    \I__6166\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28658\
        );

    \I__6165\ : Span4Mux_v
    port map (
            O => \N__28669\,
            I => \N__28654\
        );

    \I__6164\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28651\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28648\
        );

    \I__6162\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28643\
        );

    \I__6161\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28643\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28640\
        );

    \I__6159\ : InMux
    port map (
            O => \N__28657\,
            I => \N__28637\
        );

    \I__6158\ : Span4Mux_h
    port map (
            O => \N__28654\,
            I => \N__28634\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__28651\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__28648\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__28643\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__6154\ : Odrv4
    port map (
            O => \N__28640\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__28637\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__6152\ : Odrv4
    port map (
            O => \N__28634\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__6151\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28612\
        );

    \I__6150\ : InMux
    port map (
            O => \N__28620\,
            I => \N__28612\
        );

    \I__6149\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28607\
        );

    \I__6148\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28607\
        );

    \I__6147\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28604\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__28612\,
            I => \this_ppu.un1_M_state_q_2_0\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__28607\,
            I => \this_ppu.un1_M_state_q_2_0\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__28604\,
            I => \this_ppu.un1_M_state_q_2_0\
        );

    \I__6143\ : CascadeMux
    port map (
            O => \N__28597\,
            I => \N__28594\
        );

    \I__6142\ : CascadeBuf
    port map (
            O => \N__28594\,
            I => \N__28591\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__28591\,
            I => \N__28588\
        );

    \I__6140\ : InMux
    port map (
            O => \N__28588\,
            I => \N__28585\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28582\
        );

    \I__6138\ : Odrv12
    port map (
            O => \N__28582\,
            I => \this_ppu.N_19_0\
        );

    \I__6137\ : CascadeMux
    port map (
            O => \N__28579\,
            I => \this_ppu.un1_M_vaddress_q_c2_cascade_\
        );

    \I__6136\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28573\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__28573\,
            I => \M_this_data_tmp_qZ0Z_8\
        );

    \I__6134\ : InMux
    port map (
            O => \N__28570\,
            I => \N__28567\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__28567\,
            I => \N__28564\
        );

    \I__6132\ : Span4Mux_h
    port map (
            O => \N__28564\,
            I => \N__28561\
        );

    \I__6131\ : Span4Mux_h
    port map (
            O => \N__28561\,
            I => \N__28558\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__28558\,
            I => \M_this_oam_ram_write_data_8\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__28555\,
            I => \this_ppu.N_61_i_cascade_\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__28552\,
            I => \N__28549\
        );

    \I__6127\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__28546\,
            I => \N__28542\
        );

    \I__6125\ : InMux
    port map (
            O => \N__28545\,
            I => \N__28539\
        );

    \I__6124\ : Span12Mux_h
    port map (
            O => \N__28542\,
            I => \N__28536\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28533\
        );

    \I__6122\ : Odrv12
    port map (
            O => \N__28536\,
            I => \this_ppu.N_769_0\
        );

    \I__6121\ : Odrv4
    port map (
            O => \N__28533\,
            I => \this_ppu.N_769_0\
        );

    \I__6120\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28525\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__28525\,
            I => \N__28522\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__28522\,
            I => \this_ppu.M_state_q_srsts_i_i_o2_4_2\
        );

    \I__6117\ : CascadeMux
    port map (
            O => \N__28519\,
            I => \N__28516\
        );

    \I__6116\ : InMux
    port map (
            O => \N__28516\,
            I => \N__28512\
        );

    \I__6115\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28508\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__28512\,
            I => \N__28504\
        );

    \I__6113\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28501\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__28508\,
            I => \N__28498\
        );

    \I__6111\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28495\
        );

    \I__6110\ : Span4Mux_h
    port map (
            O => \N__28504\,
            I => \N__28492\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__28501\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__6108\ : Odrv4
    port map (
            O => \N__28498\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__28495\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__6106\ : Odrv4
    port map (
            O => \N__28492\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__28483\,
            I => \this_ppu.un1_M_state_q_2_0_cascade_\
        );

    \I__6104\ : CascadeMux
    port map (
            O => \N__28480\,
            I => \N__28477\
        );

    \I__6103\ : CascadeBuf
    port map (
            O => \N__28477\,
            I => \N__28474\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__28474\,
            I => \N__28471\
        );

    \I__6101\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28468\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__28468\,
            I => \N__28465\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__28465\,
            I => \N__28459\
        );

    \I__6098\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28456\
        );

    \I__6097\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28453\
        );

    \I__6096\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28450\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__28459\,
            I => \N__28447\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__28456\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__28453\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__28450\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__6091\ : Odrv4
    port map (
            O => \N__28447\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__6090\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28429\
        );

    \I__6089\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28426\
        );

    \I__6088\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28415\
        );

    \I__6087\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28415\
        );

    \I__6086\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28415\
        );

    \I__6085\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28415\
        );

    \I__6084\ : InMux
    port map (
            O => \N__28432\,
            I => \N__28415\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__28429\,
            I => \this_ppu.M_oamcurr_qc_0_1\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__28426\,
            I => \this_ppu.M_oamcurr_qc_0_1\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__28415\,
            I => \this_ppu.M_oamcurr_qc_0_1\
        );

    \I__6080\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28404\
        );

    \I__6079\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28401\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__28404\,
            I => \this_ppu.un1_M_oamcurr_q_2_c5\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__28401\,
            I => \this_ppu.un1_M_oamcurr_q_2_c5\
        );

    \I__6076\ : CascadeMux
    port map (
            O => \N__28396\,
            I => \N__28392\
        );

    \I__6075\ : CascadeMux
    port map (
            O => \N__28395\,
            I => \N__28389\
        );

    \I__6074\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28384\
        );

    \I__6073\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28384\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__28384\,
            I => \this_ppu.M_oamcurr_qZ0Z_6\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__28381\,
            I => \N__28376\
        );

    \I__6070\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28372\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28369\
        );

    \I__6068\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28366\
        );

    \I__6067\ : InMux
    port map (
            O => \N__28375\,
            I => \N__28363\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__28372\,
            I => \N__28360\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__28369\,
            I => \N__28357\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__28366\,
            I => \N__28353\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__28363\,
            I => \N__28348\
        );

    \I__6062\ : Span4Mux_v
    port map (
            O => \N__28360\,
            I => \N__28348\
        );

    \I__6061\ : Span4Mux_v
    port map (
            O => \N__28357\,
            I => \N__28344\
        );

    \I__6060\ : CascadeMux
    port map (
            O => \N__28356\,
            I => \N__28341\
        );

    \I__6059\ : Span12Mux_s10_v
    port map (
            O => \N__28353\,
            I => \N__28338\
        );

    \I__6058\ : Sp12to4
    port map (
            O => \N__28348\,
            I => \N__28335\
        );

    \I__6057\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28332\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__28344\,
            I => \N__28329\
        );

    \I__6055\ : InMux
    port map (
            O => \N__28341\,
            I => \N__28326\
        );

    \I__6054\ : Odrv12
    port map (
            O => \N__28338\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__6053\ : Odrv12
    port map (
            O => \N__28335\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__28332\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__6051\ : Odrv4
    port map (
            O => \N__28329\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__28326\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__28315\,
            I => \N__28312\
        );

    \I__6048\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28309\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__28309\,
            I => \M_this_scroll_qZ0Z_10\
        );

    \I__6046\ : InMux
    port map (
            O => \N__28306\,
            I => \this_ppu.un1_M_hoffset_d_cry_1\
        );

    \I__6045\ : CascadeMux
    port map (
            O => \N__28303\,
            I => \N__28300\
        );

    \I__6044\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28296\
        );

    \I__6043\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28292\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__28296\,
            I => \N__28289\
        );

    \I__6041\ : CascadeMux
    port map (
            O => \N__28295\,
            I => \N__28286\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__28292\,
            I => \N__28282\
        );

    \I__6039\ : Span4Mux_h
    port map (
            O => \N__28289\,
            I => \N__28279\
        );

    \I__6038\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28272\
        );

    \I__6037\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28269\
        );

    \I__6036\ : Span4Mux_v
    port map (
            O => \N__28282\,
            I => \N__28266\
        );

    \I__6035\ : Span4Mux_h
    port map (
            O => \N__28279\,
            I => \N__28263\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28260\
        );

    \I__6033\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28257\
        );

    \I__6032\ : InMux
    port map (
            O => \N__28276\,
            I => \N__28254\
        );

    \I__6031\ : InMux
    port map (
            O => \N__28275\,
            I => \N__28251\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__28272\,
            I => \N__28246\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__28269\,
            I => \N__28246\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__28266\,
            I => \N__28243\
        );

    \I__6027\ : Span4Mux_v
    port map (
            O => \N__28263\,
            I => \N__28236\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__28260\,
            I => \N__28236\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28236\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__28254\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__28251\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__6022\ : Odrv4
    port map (
            O => \N__28246\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__28243\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__6020\ : Odrv4
    port map (
            O => \N__28236\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__6019\ : CascadeMux
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__6018\ : InMux
    port map (
            O => \N__28222\,
            I => \N__28219\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__28219\,
            I => \M_this_scroll_qZ0Z_11\
        );

    \I__6016\ : InMux
    port map (
            O => \N__28216\,
            I => \this_ppu.un1_M_hoffset_d_cry_2\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__28213\,
            I => \N__28210\
        );

    \I__6014\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__28207\,
            I => \N__28203\
        );

    \I__6012\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28200\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__28203\,
            I => \N__28197\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__28200\,
            I => \N__28191\
        );

    \I__6009\ : Span4Mux_v
    port map (
            O => \N__28197\,
            I => \N__28188\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__28196\,
            I => \N__28185\
        );

    \I__6007\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28180\
        );

    \I__6006\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28180\
        );

    \I__6005\ : Span4Mux_v
    port map (
            O => \N__28191\,
            I => \N__28177\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__28188\,
            I => \N__28174\
        );

    \I__6003\ : InMux
    port map (
            O => \N__28185\,
            I => \N__28171\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28166\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__28177\,
            I => \N__28166\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__28174\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__28171\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__28166\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__28159\,
            I => \N__28156\
        );

    \I__5996\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28153\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__28153\,
            I => \N__28150\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__28150\,
            I => \M_this_scroll_qZ0Z_12\
        );

    \I__5993\ : InMux
    port map (
            O => \N__28147\,
            I => \this_ppu.un1_M_hoffset_d_cry_3\
        );

    \I__5992\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28141\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__28141\,
            I => \M_this_scroll_qZ0Z_13\
        );

    \I__5990\ : CascadeMux
    port map (
            O => \N__28138\,
            I => \N__28135\
        );

    \I__5989\ : InMux
    port map (
            O => \N__28135\,
            I => \N__28132\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__28132\,
            I => \N__28128\
        );

    \I__5987\ : CascadeMux
    port map (
            O => \N__28131\,
            I => \N__28125\
        );

    \I__5986\ : Span4Mux_h
    port map (
            O => \N__28128\,
            I => \N__28122\
        );

    \I__5985\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28119\
        );

    \I__5984\ : Span4Mux_h
    port map (
            O => \N__28122\,
            I => \N__28114\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28111\
        );

    \I__5982\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28106\
        );

    \I__5981\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28106\
        );

    \I__5980\ : Sp12to4
    port map (
            O => \N__28114\,
            I => \N__28101\
        );

    \I__5979\ : Span12Mux_h
    port map (
            O => \N__28111\,
            I => \N__28101\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__28106\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__5977\ : Odrv12
    port map (
            O => \N__28101\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__5976\ : InMux
    port map (
            O => \N__28096\,
            I => \this_ppu.un1_M_hoffset_d_cry_4\
        );

    \I__5975\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28090\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__28090\,
            I => \M_this_scroll_qZ0Z_14\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__28087\,
            I => \N__28083\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__28086\,
            I => \N__28080\
        );

    \I__5971\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28077\
        );

    \I__5970\ : InMux
    port map (
            O => \N__28080\,
            I => \N__28074\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__28077\,
            I => \N__28071\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__28074\,
            I => \N__28068\
        );

    \I__5967\ : Sp12to4
    port map (
            O => \N__28071\,
            I => \N__28063\
        );

    \I__5966\ : Span4Mux_v
    port map (
            O => \N__28068\,
            I => \N__28060\
        );

    \I__5965\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28057\
        );

    \I__5964\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28054\
        );

    \I__5963\ : Span12Mux_s9_v
    port map (
            O => \N__28063\,
            I => \N__28051\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__28060\,
            I => \N__28048\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__28057\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__28054\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__5959\ : Odrv12
    port map (
            O => \N__28051\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__28048\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__5957\ : InMux
    port map (
            O => \N__28039\,
            I => \this_ppu.un1_M_hoffset_d_cry_5\
        );

    \I__5956\ : InMux
    port map (
            O => \N__28036\,
            I => \N__28033\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__28033\,
            I => \N__28029\
        );

    \I__5954\ : InMux
    port map (
            O => \N__28032\,
            I => \N__28026\
        );

    \I__5953\ : Span4Mux_v
    port map (
            O => \N__28029\,
            I => \N__28023\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__28026\,
            I => \N__28018\
        );

    \I__5951\ : Span4Mux_v
    port map (
            O => \N__28023\,
            I => \N__28018\
        );

    \I__5950\ : Odrv4
    port map (
            O => \N__28018\,
            I => \this_ppu.M_haddress_qZ0Z_7\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__28015\,
            I => \N__28012\
        );

    \I__5948\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28009\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__28009\,
            I => \M_this_scroll_qZ0Z_15\
        );

    \I__5946\ : InMux
    port map (
            O => \N__28006\,
            I => \this_ppu.un1_M_hoffset_d_cry_6\
        );

    \I__5945\ : InMux
    port map (
            O => \N__28003\,
            I => \bfn_19_18_0_\
        );

    \I__5944\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27997\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__5942\ : Span4Mux_h
    port map (
            O => \N__27994\,
            I => \N__27991\
        );

    \I__5941\ : Span4Mux_h
    port map (
            O => \N__27991\,
            I => \N__27988\
        );

    \I__5940\ : Odrv4
    port map (
            O => \N__27988\,
            I => \this_ppu.oam_cache.mem_1\
        );

    \I__5939\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27982\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__27982\,
            I => \N__27979\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__27979\,
            I => \N__27976\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__27976\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_1\
        );

    \I__5935\ : CEMux
    port map (
            O => \N__27973\,
            I => \N__27969\
        );

    \I__5934\ : CEMux
    port map (
            O => \N__27972\,
            I => \N__27966\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N_1310_0\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__27966\,
            I => \N_1310_0\
        );

    \I__5931\ : CascadeMux
    port map (
            O => \N__27961\,
            I => \N__27958\
        );

    \I__5930\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27955\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__27955\,
            I => \N__27951\
        );

    \I__5928\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27948\
        );

    \I__5927\ : Sp12to4
    port map (
            O => \N__27951\,
            I => \N__27945\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__27948\,
            I => \N__27939\
        );

    \I__5925\ : Span12Mux_h
    port map (
            O => \N__27945\,
            I => \N__27935\
        );

    \I__5924\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27930\
        );

    \I__5923\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27930\
        );

    \I__5922\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27927\
        );

    \I__5921\ : Span12Mux_v
    port map (
            O => \N__27939\,
            I => \N__27924\
        );

    \I__5920\ : InMux
    port map (
            O => \N__27938\,
            I => \N__27921\
        );

    \I__5919\ : Odrv12
    port map (
            O => \N__27935\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__27930\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__27927\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5916\ : Odrv12
    port map (
            O => \N__27924\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__27921\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__27910\,
            I => \N__27907\
        );

    \I__5913\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27904\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__27904\,
            I => \M_this_scroll_qZ0Z_9\
        );

    \I__5911\ : InMux
    port map (
            O => \N__27901\,
            I => \this_ppu.un1_M_hoffset_d_cry_0\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__27898\,
            I => \N__27894\
        );

    \I__5909\ : CascadeMux
    port map (
            O => \N__27897\,
            I => \N__27889\
        );

    \I__5908\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27884\
        );

    \I__5907\ : CascadeMux
    port map (
            O => \N__27893\,
            I => \N__27881\
        );

    \I__5906\ : CascadeMux
    port map (
            O => \N__27892\,
            I => \N__27876\
        );

    \I__5905\ : InMux
    port map (
            O => \N__27889\,
            I => \N__27872\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__27888\,
            I => \N__27869\
        );

    \I__5903\ : CascadeMux
    port map (
            O => \N__27887\,
            I => \N__27865\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__27884\,
            I => \N__27862\
        );

    \I__5901\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27859\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__27880\,
            I => \N__27856\
        );

    \I__5899\ : CascadeMux
    port map (
            O => \N__27879\,
            I => \N__27848\
        );

    \I__5898\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27844\
        );

    \I__5897\ : CascadeMux
    port map (
            O => \N__27875\,
            I => \N__27841\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__27872\,
            I => \N__27838\
        );

    \I__5895\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27835\
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__27868\,
            I => \N__27832\
        );

    \I__5893\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27829\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__27862\,
            I => \N__27826\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__27859\,
            I => \N__27823\
        );

    \I__5890\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27820\
        );

    \I__5889\ : CascadeMux
    port map (
            O => \N__27855\,
            I => \N__27817\
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__27854\,
            I => \N__27814\
        );

    \I__5887\ : CascadeMux
    port map (
            O => \N__27853\,
            I => \N__27811\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__27852\,
            I => \N__27808\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__27851\,
            I => \N__27805\
        );

    \I__5884\ : InMux
    port map (
            O => \N__27848\,
            I => \N__27802\
        );

    \I__5883\ : CascadeMux
    port map (
            O => \N__27847\,
            I => \N__27799\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__27844\,
            I => \N__27796\
        );

    \I__5881\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27793\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__27838\,
            I => \N__27790\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__27835\,
            I => \N__27787\
        );

    \I__5878\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27784\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__27829\,
            I => \N__27781\
        );

    \I__5876\ : Span4Mux_v
    port map (
            O => \N__27826\,
            I => \N__27776\
        );

    \I__5875\ : Span4Mux_h
    port map (
            O => \N__27823\,
            I => \N__27776\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__27820\,
            I => \N__27773\
        );

    \I__5873\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27770\
        );

    \I__5872\ : InMux
    port map (
            O => \N__27814\,
            I => \N__27767\
        );

    \I__5871\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27764\
        );

    \I__5870\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27761\
        );

    \I__5869\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27758\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__27802\,
            I => \N__27755\
        );

    \I__5867\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27752\
        );

    \I__5866\ : Span4Mux_h
    port map (
            O => \N__27796\,
            I => \N__27749\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__27793\,
            I => \N__27746\
        );

    \I__5864\ : Span4Mux_v
    port map (
            O => \N__27790\,
            I => \N__27741\
        );

    \I__5863\ : Span4Mux_h
    port map (
            O => \N__27787\,
            I => \N__27741\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27738\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__27781\,
            I => \N__27735\
        );

    \I__5860\ : Span4Mux_v
    port map (
            O => \N__27776\,
            I => \N__27730\
        );

    \I__5859\ : Span4Mux_h
    port map (
            O => \N__27773\,
            I => \N__27730\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__27770\,
            I => \N__27727\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__27767\,
            I => \N__27718\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__27764\,
            I => \N__27718\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__27761\,
            I => \N__27718\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__27758\,
            I => \N__27718\
        );

    \I__5853\ : Sp12to4
    port map (
            O => \N__27755\,
            I => \N__27713\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__27752\,
            I => \N__27713\
        );

    \I__5851\ : Span4Mux_v
    port map (
            O => \N__27749\,
            I => \N__27708\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__27746\,
            I => \N__27708\
        );

    \I__5849\ : Span4Mux_v
    port map (
            O => \N__27741\,
            I => \N__27703\
        );

    \I__5848\ : Span4Mux_h
    port map (
            O => \N__27738\,
            I => \N__27703\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__27735\,
            I => \N__27696\
        );

    \I__5846\ : Span4Mux_v
    port map (
            O => \N__27730\,
            I => \N__27696\
        );

    \I__5845\ : Span4Mux_h
    port map (
            O => \N__27727\,
            I => \N__27696\
        );

    \I__5844\ : Span12Mux_v
    port map (
            O => \N__27718\,
            I => \N__27690\
        );

    \I__5843\ : Span12Mux_v
    port map (
            O => \N__27713\,
            I => \N__27690\
        );

    \I__5842\ : Span4Mux_h
    port map (
            O => \N__27708\,
            I => \N__27685\
        );

    \I__5841\ : Span4Mux_h
    port map (
            O => \N__27703\,
            I => \N__27685\
        );

    \I__5840\ : Span4Mux_h
    port map (
            O => \N__27696\,
            I => \N__27682\
        );

    \I__5839\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27679\
        );

    \I__5838\ : Odrv12
    port map (
            O => \N__27690\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__27685\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__27682\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__27679\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__5834\ : InMux
    port map (
            O => \N__27670\,
            I => \un1_M_this_spr_address_q_cry_6\
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__27667\,
            I => \N__27663\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__27666\,
            I => \N__27659\
        );

    \I__5831\ : InMux
    port map (
            O => \N__27663\,
            I => \N__27655\
        );

    \I__5830\ : CascadeMux
    port map (
            O => \N__27662\,
            I => \N__27652\
        );

    \I__5829\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27647\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__27658\,
            I => \N__27644\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__27655\,
            I => \N__27639\
        );

    \I__5826\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27636\
        );

    \I__5825\ : CascadeMux
    port map (
            O => \N__27651\,
            I => \N__27633\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__27650\,
            I => \N__27630\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__27647\,
            I => \N__27626\
        );

    \I__5822\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27623\
        );

    \I__5821\ : CascadeMux
    port map (
            O => \N__27643\,
            I => \N__27620\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__27642\,
            I => \N__27616\
        );

    \I__5819\ : Span4Mux_h
    port map (
            O => \N__27639\,
            I => \N__27606\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__27636\,
            I => \N__27606\
        );

    \I__5817\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27603\
        );

    \I__5816\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27600\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__27629\,
            I => \N__27597\
        );

    \I__5814\ : Span4Mux_v
    port map (
            O => \N__27626\,
            I => \N__27592\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__27623\,
            I => \N__27592\
        );

    \I__5812\ : InMux
    port map (
            O => \N__27620\,
            I => \N__27589\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__27619\,
            I => \N__27586\
        );

    \I__5810\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27583\
        );

    \I__5809\ : CascadeMux
    port map (
            O => \N__27615\,
            I => \N__27580\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__27614\,
            I => \N__27577\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__27613\,
            I => \N__27574\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__27612\,
            I => \N__27571\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__27611\,
            I => \N__27568\
        );

    \I__5804\ : Span4Mux_v
    port map (
            O => \N__27606\,
            I => \N__27563\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__27603\,
            I => \N__27563\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27560\
        );

    \I__5801\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27557\
        );

    \I__5800\ : Span4Mux_h
    port map (
            O => \N__27592\,
            I => \N__27552\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27552\
        );

    \I__5798\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27549\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__27583\,
            I => \N__27546\
        );

    \I__5796\ : InMux
    port map (
            O => \N__27580\,
            I => \N__27543\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27540\
        );

    \I__5794\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27536\
        );

    \I__5793\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27533\
        );

    \I__5792\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27530\
        );

    \I__5791\ : Span4Mux_v
    port map (
            O => \N__27563\,
            I => \N__27525\
        );

    \I__5790\ : Span4Mux_v
    port map (
            O => \N__27560\,
            I => \N__27525\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__27557\,
            I => \N__27522\
        );

    \I__5788\ : Span4Mux_v
    port map (
            O => \N__27552\,
            I => \N__27517\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__27549\,
            I => \N__27517\
        );

    \I__5786\ : Span4Mux_v
    port map (
            O => \N__27546\,
            I => \N__27510\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__27543\,
            I => \N__27510\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27510\
        );

    \I__5783\ : CascadeMux
    port map (
            O => \N__27539\,
            I => \N__27507\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__27536\,
            I => \N__27504\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__27533\,
            I => \N__27501\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__27530\,
            I => \N__27498\
        );

    \I__5779\ : Sp12to4
    port map (
            O => \N__27525\,
            I => \N__27493\
        );

    \I__5778\ : Sp12to4
    port map (
            O => \N__27522\,
            I => \N__27493\
        );

    \I__5777\ : Span4Mux_v
    port map (
            O => \N__27517\,
            I => \N__27488\
        );

    \I__5776\ : Span4Mux_v
    port map (
            O => \N__27510\,
            I => \N__27488\
        );

    \I__5775\ : InMux
    port map (
            O => \N__27507\,
            I => \N__27485\
        );

    \I__5774\ : Span12Mux_h
    port map (
            O => \N__27504\,
            I => \N__27481\
        );

    \I__5773\ : Span12Mux_h
    port map (
            O => \N__27501\,
            I => \N__27476\
        );

    \I__5772\ : Span12Mux_h
    port map (
            O => \N__27498\,
            I => \N__27476\
        );

    \I__5771\ : Span12Mux_h
    port map (
            O => \N__27493\,
            I => \N__27469\
        );

    \I__5770\ : Sp12to4
    port map (
            O => \N__27488\,
            I => \N__27469\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__27485\,
            I => \N__27469\
        );

    \I__5768\ : InMux
    port map (
            O => \N__27484\,
            I => \N__27466\
        );

    \I__5767\ : Odrv12
    port map (
            O => \N__27481\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__5766\ : Odrv12
    port map (
            O => \N__27476\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__5765\ : Odrv12
    port map (
            O => \N__27469\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__27466\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__5763\ : InMux
    port map (
            O => \N__27457\,
            I => \bfn_19_14_0_\
        );

    \I__5762\ : CascadeMux
    port map (
            O => \N__27454\,
            I => \N__27450\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__27453\,
            I => \N__27446\
        );

    \I__5760\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27442\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__27449\,
            I => \N__27439\
        );

    \I__5758\ : InMux
    port map (
            O => \N__27446\,
            I => \N__27435\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__27445\,
            I => \N__27432\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27428\
        );

    \I__5755\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27425\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__27438\,
            I => \N__27422\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__27435\,
            I => \N__27417\
        );

    \I__5752\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27414\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__27431\,
            I => \N__27411\
        );

    \I__5750\ : Span4Mux_h
    port map (
            O => \N__27428\,
            I => \N__27403\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__27425\,
            I => \N__27403\
        );

    \I__5748\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27400\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__27421\,
            I => \N__27397\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__27420\,
            I => \N__27394\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__27417\,
            I => \N__27388\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__27414\,
            I => \N__27388\
        );

    \I__5743\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27385\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__27410\,
            I => \N__27382\
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__27409\,
            I => \N__27378\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__27408\,
            I => \N__27373\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__27403\,
            I => \N__27368\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27368\
        );

    \I__5737\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27365\
        );

    \I__5736\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27362\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__27393\,
            I => \N__27359\
        );

    \I__5734\ : Span4Mux_h
    port map (
            O => \N__27388\,
            I => \N__27354\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__27385\,
            I => \N__27354\
        );

    \I__5732\ : InMux
    port map (
            O => \N__27382\,
            I => \N__27351\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__27381\,
            I => \N__27348\
        );

    \I__5730\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27345\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__27377\,
            I => \N__27342\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__27376\,
            I => \N__27339\
        );

    \I__5727\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27336\
        );

    \I__5726\ : Span4Mux_h
    port map (
            O => \N__27368\,
            I => \N__27331\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__27365\,
            I => \N__27331\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27328\
        );

    \I__5723\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27325\
        );

    \I__5722\ : Span4Mux_v
    port map (
            O => \N__27354\,
            I => \N__27320\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__27351\,
            I => \N__27320\
        );

    \I__5720\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27317\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27314\
        );

    \I__5718\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27311\
        );

    \I__5717\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27308\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__27336\,
            I => \N__27304\
        );

    \I__5715\ : Span4Mux_v
    port map (
            O => \N__27331\,
            I => \N__27297\
        );

    \I__5714\ : Span4Mux_v
    port map (
            O => \N__27328\,
            I => \N__27297\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27297\
        );

    \I__5712\ : Span4Mux_h
    port map (
            O => \N__27320\,
            I => \N__27292\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__27317\,
            I => \N__27292\
        );

    \I__5710\ : Span4Mux_v
    port map (
            O => \N__27314\,
            I => \N__27285\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__27311\,
            I => \N__27285\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27285\
        );

    \I__5707\ : CascadeMux
    port map (
            O => \N__27307\,
            I => \N__27282\
        );

    \I__5706\ : Span12Mux_h
    port map (
            O => \N__27304\,
            I => \N__27279\
        );

    \I__5705\ : Sp12to4
    port map (
            O => \N__27297\,
            I => \N__27276\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__27292\,
            I => \N__27271\
        );

    \I__5703\ : Span4Mux_v
    port map (
            O => \N__27285\,
            I => \N__27271\
        );

    \I__5702\ : InMux
    port map (
            O => \N__27282\,
            I => \N__27268\
        );

    \I__5701\ : Span12Mux_v
    port map (
            O => \N__27279\,
            I => \N__27258\
        );

    \I__5700\ : Span12Mux_h
    port map (
            O => \N__27276\,
            I => \N__27258\
        );

    \I__5699\ : Sp12to4
    port map (
            O => \N__27271\,
            I => \N__27258\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__27268\,
            I => \N__27258\
        );

    \I__5697\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27255\
        );

    \I__5696\ : Odrv12
    port map (
            O => \N__27258\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__27255\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__5694\ : InMux
    port map (
            O => \N__27250\,
            I => \un1_M_this_spr_address_q_cry_8\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__27247\,
            I => \N__27244\
        );

    \I__5692\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27240\
        );

    \I__5691\ : CascadeMux
    port map (
            O => \N__27243\,
            I => \N__27237\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__27240\,
            I => \N__27230\
        );

    \I__5689\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27227\
        );

    \I__5688\ : CascadeMux
    port map (
            O => \N__27236\,
            I => \N__27224\
        );

    \I__5687\ : CascadeMux
    port map (
            O => \N__27235\,
            I => \N__27218\
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__27234\,
            I => \N__27215\
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__27233\,
            I => \N__27210\
        );

    \I__5684\ : Span4Mux_h
    port map (
            O => \N__27230\,
            I => \N__27204\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__27227\,
            I => \N__27204\
        );

    \I__5682\ : InMux
    port map (
            O => \N__27224\,
            I => \N__27201\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__27223\,
            I => \N__27198\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__27222\,
            I => \N__27195\
        );

    \I__5679\ : CascadeMux
    port map (
            O => \N__27221\,
            I => \N__27190\
        );

    \I__5678\ : InMux
    port map (
            O => \N__27218\,
            I => \N__27187\
        );

    \I__5677\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27183\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__27214\,
            I => \N__27180\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__27213\,
            I => \N__27177\
        );

    \I__5674\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27173\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__27209\,
            I => \N__27170\
        );

    \I__5672\ : Span4Mux_v
    port map (
            O => \N__27204\,
            I => \N__27165\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__27201\,
            I => \N__27165\
        );

    \I__5670\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27162\
        );

    \I__5669\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27159\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__27194\,
            I => \N__27156\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__27193\,
            I => \N__27153\
        );

    \I__5666\ : InMux
    port map (
            O => \N__27190\,
            I => \N__27150\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__27187\,
            I => \N__27147\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__27186\,
            I => \N__27144\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__27183\,
            I => \N__27141\
        );

    \I__5662\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27138\
        );

    \I__5661\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27135\
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__27176\,
            I => \N__27132\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__27173\,
            I => \N__27129\
        );

    \I__5658\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27126\
        );

    \I__5657\ : Span4Mux_h
    port map (
            O => \N__27165\,
            I => \N__27123\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__27162\,
            I => \N__27120\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__27159\,
            I => \N__27117\
        );

    \I__5654\ : InMux
    port map (
            O => \N__27156\,
            I => \N__27114\
        );

    \I__5653\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27111\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__27150\,
            I => \N__27108\
        );

    \I__5651\ : Span4Mux_v
    port map (
            O => \N__27147\,
            I => \N__27105\
        );

    \I__5650\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27102\
        );

    \I__5649\ : Span4Mux_h
    port map (
            O => \N__27141\,
            I => \N__27099\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__27138\,
            I => \N__27096\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__27135\,
            I => \N__27093\
        );

    \I__5646\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27090\
        );

    \I__5645\ : Span12Mux_s1_v
    port map (
            O => \N__27129\,
            I => \N__27085\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__27126\,
            I => \N__27085\
        );

    \I__5643\ : Span4Mux_v
    port map (
            O => \N__27123\,
            I => \N__27080\
        );

    \I__5642\ : Span4Mux_h
    port map (
            O => \N__27120\,
            I => \N__27080\
        );

    \I__5641\ : Sp12to4
    port map (
            O => \N__27117\,
            I => \N__27077\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__27114\,
            I => \N__27074\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__27111\,
            I => \N__27071\
        );

    \I__5638\ : Span12Mux_h
    port map (
            O => \N__27108\,
            I => \N__27064\
        );

    \I__5637\ : Sp12to4
    port map (
            O => \N__27105\,
            I => \N__27064\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__27102\,
            I => \N__27064\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__27099\,
            I => \N__27059\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__27096\,
            I => \N__27059\
        );

    \I__5633\ : Span4Mux_h
    port map (
            O => \N__27093\,
            I => \N__27056\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__27090\,
            I => \N__27053\
        );

    \I__5631\ : Span12Mux_v
    port map (
            O => \N__27085\,
            I => \N__27049\
        );

    \I__5630\ : Span4Mux_h
    port map (
            O => \N__27080\,
            I => \N__27046\
        );

    \I__5629\ : Span12Mux_h
    port map (
            O => \N__27077\,
            I => \N__27041\
        );

    \I__5628\ : Span12Mux_h
    port map (
            O => \N__27074\,
            I => \N__27041\
        );

    \I__5627\ : Span12Mux_h
    port map (
            O => \N__27071\,
            I => \N__27036\
        );

    \I__5626\ : Span12Mux_h
    port map (
            O => \N__27064\,
            I => \N__27036\
        );

    \I__5625\ : Span4Mux_v
    port map (
            O => \N__27059\,
            I => \N__27029\
        );

    \I__5624\ : Span4Mux_v
    port map (
            O => \N__27056\,
            I => \N__27029\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__27053\,
            I => \N__27029\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27026\
        );

    \I__5621\ : Odrv12
    port map (
            O => \N__27049\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__27046\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__5619\ : Odrv12
    port map (
            O => \N__27041\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__5618\ : Odrv12
    port map (
            O => \N__27036\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__27029\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__27026\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__5615\ : InMux
    port map (
            O => \N__27013\,
            I => \un1_M_this_spr_address_q_cry_9\
        );

    \I__5614\ : InMux
    port map (
            O => \N__27010\,
            I => \un1_M_this_spr_address_q_cry_10\
        );

    \I__5613\ : InMux
    port map (
            O => \N__27007\,
            I => \un1_M_this_spr_address_q_cry_11\
        );

    \I__5612\ : InMux
    port map (
            O => \N__27004\,
            I => \un1_M_this_spr_address_q_cry_12\
        );

    \I__5611\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26998\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__26998\,
            I => \M_this_data_tmp_qZ0Z_18\
        );

    \I__5609\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26992\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__26992\,
            I => \N__26989\
        );

    \I__5607\ : Span4Mux_h
    port map (
            O => \N__26989\,
            I => \N__26986\
        );

    \I__5606\ : Span4Mux_h
    port map (
            O => \N__26986\,
            I => \N__26983\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__26983\,
            I => \M_this_oam_ram_write_data_18\
        );

    \I__5604\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26977\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__26977\,
            I => \M_this_data_tmp_qZ0Z_21\
        );

    \I__5602\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26971\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__26971\,
            I => \N__26968\
        );

    \I__5600\ : Span4Mux_v
    port map (
            O => \N__26968\,
            I => \N__26965\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__26965\,
            I => \N__26962\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__26962\,
            I => \M_this_oam_ram_write_data_21\
        );

    \I__5597\ : CascadeMux
    port map (
            O => \N__26959\,
            I => \N__26951\
        );

    \I__5596\ : CascadeMux
    port map (
            O => \N__26958\,
            I => \N__26948\
        );

    \I__5595\ : CascadeMux
    port map (
            O => \N__26957\,
            I => \N__26941\
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__26956\,
            I => \N__26938\
        );

    \I__5593\ : CascadeMux
    port map (
            O => \N__26955\,
            I => \N__26933\
        );

    \I__5592\ : CascadeMux
    port map (
            O => \N__26954\,
            I => \N__26930\
        );

    \I__5591\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26927\
        );

    \I__5590\ : InMux
    port map (
            O => \N__26948\,
            I => \N__26924\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__26947\,
            I => \N__26921\
        );

    \I__5588\ : CascadeMux
    port map (
            O => \N__26946\,
            I => \N__26918\
        );

    \I__5587\ : CascadeMux
    port map (
            O => \N__26945\,
            I => \N__26915\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__26944\,
            I => \N__26912\
        );

    \I__5585\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26908\
        );

    \I__5584\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26905\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__26937\,
            I => \N__26902\
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__26936\,
            I => \N__26899\
        );

    \I__5581\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26894\
        );

    \I__5580\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26890\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__26927\,
            I => \N__26885\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__26924\,
            I => \N__26885\
        );

    \I__5577\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26882\
        );

    \I__5576\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26879\
        );

    \I__5575\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26876\
        );

    \I__5574\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26873\
        );

    \I__5573\ : CascadeMux
    port map (
            O => \N__26911\,
            I => \N__26870\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__26908\,
            I => \N__26865\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__26905\,
            I => \N__26865\
        );

    \I__5570\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26862\
        );

    \I__5569\ : InMux
    port map (
            O => \N__26899\,
            I => \N__26859\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__26898\,
            I => \N__26856\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__26897\,
            I => \N__26853\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__26894\,
            I => \N__26850\
        );

    \I__5565\ : CascadeMux
    port map (
            O => \N__26893\,
            I => \N__26847\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__26890\,
            I => \N__26844\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__26885\,
            I => \N__26837\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__26882\,
            I => \N__26837\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__26879\,
            I => \N__26837\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__26876\,
            I => \N__26832\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__26873\,
            I => \N__26832\
        );

    \I__5558\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26829\
        );

    \I__5557\ : Span4Mux_v
    port map (
            O => \N__26865\,
            I => \N__26822\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__26862\,
            I => \N__26822\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__26859\,
            I => \N__26822\
        );

    \I__5554\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26819\
        );

    \I__5553\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26816\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__26850\,
            I => \N__26813\
        );

    \I__5551\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26810\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__26844\,
            I => \N__26805\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__26837\,
            I => \N__26805\
        );

    \I__5548\ : Span4Mux_v
    port map (
            O => \N__26832\,
            I => \N__26800\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__26829\,
            I => \N__26800\
        );

    \I__5546\ : Span4Mux_v
    port map (
            O => \N__26822\,
            I => \N__26793\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__26819\,
            I => \N__26793\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__26816\,
            I => \N__26793\
        );

    \I__5543\ : Span4Mux_h
    port map (
            O => \N__26813\,
            I => \N__26790\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__26810\,
            I => \N__26787\
        );

    \I__5541\ : Span4Mux_h
    port map (
            O => \N__26805\,
            I => \N__26784\
        );

    \I__5540\ : Span4Mux_v
    port map (
            O => \N__26800\,
            I => \N__26781\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__26793\,
            I => \N__26778\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__26790\,
            I => \N__26773\
        );

    \I__5537\ : Span4Mux_h
    port map (
            O => \N__26787\,
            I => \N__26773\
        );

    \I__5536\ : Span4Mux_h
    port map (
            O => \N__26784\,
            I => \N__26769\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__26781\,
            I => \N__26764\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__26778\,
            I => \N__26764\
        );

    \I__5533\ : Span4Mux_h
    port map (
            O => \N__26773\,
            I => \N__26761\
        );

    \I__5532\ : InMux
    port map (
            O => \N__26772\,
            I => \N__26758\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__26769\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__26764\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__26761\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__26758\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__26749\,
            I => \N__26742\
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__26748\,
            I => \N__26737\
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__26747\,
            I => \N__26732\
        );

    \I__5524\ : CascadeMux
    port map (
            O => \N__26746\,
            I => \N__26727\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__26745\,
            I => \N__26722\
        );

    \I__5522\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26718\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__26741\,
            I => \N__26715\
        );

    \I__5520\ : CascadeMux
    port map (
            O => \N__26740\,
            I => \N__26712\
        );

    \I__5519\ : InMux
    port map (
            O => \N__26737\,
            I => \N__26709\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__26736\,
            I => \N__26706\
        );

    \I__5517\ : CascadeMux
    port map (
            O => \N__26735\,
            I => \N__26703\
        );

    \I__5516\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26700\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__26731\,
            I => \N__26697\
        );

    \I__5514\ : CascadeMux
    port map (
            O => \N__26730\,
            I => \N__26694\
        );

    \I__5513\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26691\
        );

    \I__5512\ : CascadeMux
    port map (
            O => \N__26726\,
            I => \N__26688\
        );

    \I__5511\ : CascadeMux
    port map (
            O => \N__26725\,
            I => \N__26685\
        );

    \I__5510\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26682\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__26721\,
            I => \N__26679\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26676\
        );

    \I__5507\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26673\
        );

    \I__5506\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26668\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__26709\,
            I => \N__26665\
        );

    \I__5504\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26662\
        );

    \I__5503\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26659\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__26700\,
            I => \N__26656\
        );

    \I__5501\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26653\
        );

    \I__5500\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26650\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__26691\,
            I => \N__26647\
        );

    \I__5498\ : InMux
    port map (
            O => \N__26688\,
            I => \N__26644\
        );

    \I__5497\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26641\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__26682\,
            I => \N__26638\
        );

    \I__5495\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26635\
        );

    \I__5494\ : Span4Mux_v
    port map (
            O => \N__26676\,
            I => \N__26630\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__26673\,
            I => \N__26630\
        );

    \I__5492\ : CascadeMux
    port map (
            O => \N__26672\,
            I => \N__26627\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__26671\,
            I => \N__26624\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__26668\,
            I => \N__26617\
        );

    \I__5489\ : Span4Mux_v
    port map (
            O => \N__26665\,
            I => \N__26617\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26617\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__26659\,
            I => \N__26614\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__26656\,
            I => \N__26611\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__26653\,
            I => \N__26608\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__26650\,
            I => \N__26603\
        );

    \I__5483\ : Span4Mux_v
    port map (
            O => \N__26647\,
            I => \N__26603\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__26644\,
            I => \N__26596\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__26641\,
            I => \N__26596\
        );

    \I__5480\ : Span4Mux_v
    port map (
            O => \N__26638\,
            I => \N__26596\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__26635\,
            I => \N__26591\
        );

    \I__5478\ : Span4Mux_h
    port map (
            O => \N__26630\,
            I => \N__26591\
        );

    \I__5477\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26588\
        );

    \I__5476\ : InMux
    port map (
            O => \N__26624\,
            I => \N__26585\
        );

    \I__5475\ : Span4Mux_v
    port map (
            O => \N__26617\,
            I => \N__26580\
        );

    \I__5474\ : Span4Mux_v
    port map (
            O => \N__26614\,
            I => \N__26580\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__26611\,
            I => \N__26577\
        );

    \I__5472\ : Sp12to4
    port map (
            O => \N__26608\,
            I => \N__26573\
        );

    \I__5471\ : Span4Mux_v
    port map (
            O => \N__26603\,
            I => \N__26568\
        );

    \I__5470\ : Span4Mux_v
    port map (
            O => \N__26596\,
            I => \N__26568\
        );

    \I__5469\ : Sp12to4
    port map (
            O => \N__26591\,
            I => \N__26565\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__26588\,
            I => \N__26562\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__26585\,
            I => \N__26557\
        );

    \I__5466\ : Sp12to4
    port map (
            O => \N__26580\,
            I => \N__26557\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__26577\,
            I => \N__26554\
        );

    \I__5464\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26551\
        );

    \I__5463\ : Span12Mux_v
    port map (
            O => \N__26573\,
            I => \N__26544\
        );

    \I__5462\ : Sp12to4
    port map (
            O => \N__26568\,
            I => \N__26544\
        );

    \I__5461\ : Span12Mux_v
    port map (
            O => \N__26565\,
            I => \N__26544\
        );

    \I__5460\ : Span12Mux_h
    port map (
            O => \N__26562\,
            I => \N__26539\
        );

    \I__5459\ : Span12Mux_h
    port map (
            O => \N__26557\,
            I => \N__26539\
        );

    \I__5458\ : Span4Mux_h
    port map (
            O => \N__26554\,
            I => \N__26536\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__26551\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__5456\ : Odrv12
    port map (
            O => \N__26544\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__5455\ : Odrv12
    port map (
            O => \N__26539\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__5454\ : Odrv4
    port map (
            O => \N__26536\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__5453\ : InMux
    port map (
            O => \N__26527\,
            I => \un1_M_this_spr_address_q_cry_0\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__26524\,
            I => \N__26518\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__26523\,
            I => \N__26515\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__26522\,
            I => \N__26509\
        );

    \I__5449\ : CascadeMux
    port map (
            O => \N__26521\,
            I => \N__26505\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26502\
        );

    \I__5447\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26499\
        );

    \I__5446\ : CascadeMux
    port map (
            O => \N__26514\,
            I => \N__26496\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__26513\,
            I => \N__26493\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__26512\,
            I => \N__26490\
        );

    \I__5443\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26486\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__26508\,
            I => \N__26483\
        );

    \I__5441\ : InMux
    port map (
            O => \N__26505\,
            I => \N__26479\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26474\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__26499\,
            I => \N__26474\
        );

    \I__5438\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26471\
        );

    \I__5437\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26468\
        );

    \I__5436\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26460\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__26489\,
            I => \N__26457\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26453\
        );

    \I__5433\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26450\
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__26482\,
            I => \N__26447\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__26479\,
            I => \N__26444\
        );

    \I__5430\ : Span4Mux_v
    port map (
            O => \N__26474\,
            I => \N__26437\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__26471\,
            I => \N__26437\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26437\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__26467\,
            I => \N__26434\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__26466\,
            I => \N__26431\
        );

    \I__5425\ : CascadeMux
    port map (
            O => \N__26465\,
            I => \N__26428\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__26464\,
            I => \N__26425\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__26463\,
            I => \N__26422\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__26460\,
            I => \N__26419\
        );

    \I__5421\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26416\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__26456\,
            I => \N__26413\
        );

    \I__5419\ : Span4Mux_h
    port map (
            O => \N__26453\,
            I => \N__26410\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__26450\,
            I => \N__26407\
        );

    \I__5417\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26404\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__26444\,
            I => \N__26399\
        );

    \I__5415\ : Span4Mux_v
    port map (
            O => \N__26437\,
            I => \N__26399\
        );

    \I__5414\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26396\
        );

    \I__5413\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26393\
        );

    \I__5412\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26390\
        );

    \I__5411\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26387\
        );

    \I__5410\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26384\
        );

    \I__5409\ : Span4Mux_v
    port map (
            O => \N__26419\,
            I => \N__26379\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__26416\,
            I => \N__26379\
        );

    \I__5407\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26376\
        );

    \I__5406\ : Span4Mux_h
    port map (
            O => \N__26410\,
            I => \N__26373\
        );

    \I__5405\ : Span4Mux_h
    port map (
            O => \N__26407\,
            I => \N__26370\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26367\
        );

    \I__5403\ : Span4Mux_h
    port map (
            O => \N__26399\,
            I => \N__26364\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__26396\,
            I => \N__26357\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__26393\,
            I => \N__26357\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26357\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__26387\,
            I => \N__26348\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__26384\,
            I => \N__26348\
        );

    \I__5397\ : Sp12to4
    port map (
            O => \N__26379\,
            I => \N__26348\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__26376\,
            I => \N__26348\
        );

    \I__5395\ : Span4Mux_h
    port map (
            O => \N__26373\,
            I => \N__26341\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__26370\,
            I => \N__26341\
        );

    \I__5393\ : Span4Mux_h
    port map (
            O => \N__26367\,
            I => \N__26341\
        );

    \I__5392\ : Sp12to4
    port map (
            O => \N__26364\,
            I => \N__26333\
        );

    \I__5391\ : Span12Mux_v
    port map (
            O => \N__26357\,
            I => \N__26333\
        );

    \I__5390\ : Span12Mux_v
    port map (
            O => \N__26348\,
            I => \N__26333\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__26341\,
            I => \N__26330\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26327\
        );

    \I__5387\ : Odrv12
    port map (
            O => \N__26333\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5386\ : Odrv4
    port map (
            O => \N__26330\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__26327\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5384\ : InMux
    port map (
            O => \N__26320\,
            I => \un1_M_this_spr_address_q_cry_1\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__26317\,
            I => \N__26313\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__26316\,
            I => \N__26309\
        );

    \I__5381\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26304\
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__26312\,
            I => \N__26301\
        );

    \I__5379\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26294\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__26308\,
            I => \N__26291\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__26307\,
            I => \N__26288\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26304\,
            I => \N__26285\
        );

    \I__5375\ : InMux
    port map (
            O => \N__26301\,
            I => \N__26282\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__26300\,
            I => \N__26279\
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__26299\,
            I => \N__26275\
        );

    \I__5372\ : CascadeMux
    port map (
            O => \N__26298\,
            I => \N__26271\
        );

    \I__5371\ : CascadeMux
    port map (
            O => \N__26297\,
            I => \N__26268\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__26294\,
            I => \N__26265\
        );

    \I__5369\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26262\
        );

    \I__5368\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26258\
        );

    \I__5367\ : Span4Mux_h
    port map (
            O => \N__26285\,
            I => \N__26255\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26282\,
            I => \N__26252\
        );

    \I__5365\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26249\
        );

    \I__5364\ : CascadeMux
    port map (
            O => \N__26278\,
            I => \N__26246\
        );

    \I__5363\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26243\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__26274\,
            I => \N__26240\
        );

    \I__5361\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26236\
        );

    \I__5360\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26232\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__26265\,
            I => \N__26228\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__26262\,
            I => \N__26225\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__26261\,
            I => \N__26222\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__26258\,
            I => \N__26219\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__26255\,
            I => \N__26213\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__26252\,
            I => \N__26213\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__26249\,
            I => \N__26210\
        );

    \I__5352\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26207\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__26243\,
            I => \N__26204\
        );

    \I__5350\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26201\
        );

    \I__5349\ : CascadeMux
    port map (
            O => \N__26239\,
            I => \N__26198\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__26236\,
            I => \N__26195\
        );

    \I__5347\ : CascadeMux
    port map (
            O => \N__26235\,
            I => \N__26192\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__26232\,
            I => \N__26189\
        );

    \I__5345\ : CascadeMux
    port map (
            O => \N__26231\,
            I => \N__26186\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__26228\,
            I => \N__26181\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__26225\,
            I => \N__26181\
        );

    \I__5342\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26178\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__26219\,
            I => \N__26175\
        );

    \I__5340\ : CascadeMux
    port map (
            O => \N__26218\,
            I => \N__26172\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__26213\,
            I => \N__26167\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__26210\,
            I => \N__26167\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__26207\,
            I => \N__26164\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__26204\,
            I => \N__26161\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__26201\,
            I => \N__26158\
        );

    \I__5334\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26155\
        );

    \I__5333\ : Span4Mux_s3_v
    port map (
            O => \N__26195\,
            I => \N__26152\
        );

    \I__5332\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26149\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__26189\,
            I => \N__26146\
        );

    \I__5330\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26143\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__26181\,
            I => \N__26138\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__26178\,
            I => \N__26138\
        );

    \I__5327\ : Span4Mux_v
    port map (
            O => \N__26175\,
            I => \N__26135\
        );

    \I__5326\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26132\
        );

    \I__5325\ : Span4Mux_h
    port map (
            O => \N__26167\,
            I => \N__26129\
        );

    \I__5324\ : Span4Mux_h
    port map (
            O => \N__26164\,
            I => \N__26126\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__26161\,
            I => \N__26121\
        );

    \I__5322\ : Span4Mux_h
    port map (
            O => \N__26158\,
            I => \N__26121\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__26155\,
            I => \N__26118\
        );

    \I__5320\ : Sp12to4
    port map (
            O => \N__26152\,
            I => \N__26113\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__26149\,
            I => \N__26113\
        );

    \I__5318\ : Sp12to4
    port map (
            O => \N__26146\,
            I => \N__26108\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__26143\,
            I => \N__26108\
        );

    \I__5316\ : Sp12to4
    port map (
            O => \N__26138\,
            I => \N__26105\
        );

    \I__5315\ : Sp12to4
    port map (
            O => \N__26135\,
            I => \N__26100\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26100\
        );

    \I__5313\ : Span4Mux_h
    port map (
            O => \N__26129\,
            I => \N__26091\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__26126\,
            I => \N__26091\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__26121\,
            I => \N__26091\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__26118\,
            I => \N__26091\
        );

    \I__5309\ : Span12Mux_h
    port map (
            O => \N__26113\,
            I => \N__26085\
        );

    \I__5308\ : Span12Mux_h
    port map (
            O => \N__26108\,
            I => \N__26085\
        );

    \I__5307\ : Span12Mux_h
    port map (
            O => \N__26105\,
            I => \N__26080\
        );

    \I__5306\ : Span12Mux_h
    port map (
            O => \N__26100\,
            I => \N__26080\
        );

    \I__5305\ : Span4Mux_h
    port map (
            O => \N__26091\,
            I => \N__26077\
        );

    \I__5304\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26074\
        );

    \I__5303\ : Odrv12
    port map (
            O => \N__26085\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__5302\ : Odrv12
    port map (
            O => \N__26080\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__5301\ : Odrv4
    port map (
            O => \N__26077\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__26074\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__5299\ : InMux
    port map (
            O => \N__26065\,
            I => \un1_M_this_spr_address_q_cry_2\
        );

    \I__5298\ : CascadeMux
    port map (
            O => \N__26062\,
            I => \N__26056\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__26061\,
            I => \N__26053\
        );

    \I__5296\ : CascadeMux
    port map (
            O => \N__26060\,
            I => \N__26046\
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__26059\,
            I => \N__26043\
        );

    \I__5294\ : InMux
    port map (
            O => \N__26056\,
            I => \N__26036\
        );

    \I__5293\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26033\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__26052\,
            I => \N__26030\
        );

    \I__5291\ : CascadeMux
    port map (
            O => \N__26051\,
            I => \N__26027\
        );

    \I__5290\ : CascadeMux
    port map (
            O => \N__26050\,
            I => \N__26024\
        );

    \I__5289\ : CascadeMux
    port map (
            O => \N__26049\,
            I => \N__26021\
        );

    \I__5288\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26018\
        );

    \I__5287\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26015\
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__26042\,
            I => \N__26012\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__26041\,
            I => \N__26009\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__26040\,
            I => \N__26004\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__26039\,
            I => \N__26001\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__26036\,
            I => \N__25994\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__26033\,
            I => \N__25994\
        );

    \I__5280\ : InMux
    port map (
            O => \N__26030\,
            I => \N__25991\
        );

    \I__5279\ : InMux
    port map (
            O => \N__26027\,
            I => \N__25988\
        );

    \I__5278\ : InMux
    port map (
            O => \N__26024\,
            I => \N__25985\
        );

    \I__5277\ : InMux
    port map (
            O => \N__26021\,
            I => \N__25982\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__26018\,
            I => \N__25977\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__26015\,
            I => \N__25977\
        );

    \I__5274\ : InMux
    port map (
            O => \N__26012\,
            I => \N__25974\
        );

    \I__5273\ : InMux
    port map (
            O => \N__26009\,
            I => \N__25971\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__26008\,
            I => \N__25968\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__26007\,
            I => \N__25965\
        );

    \I__5270\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25962\
        );

    \I__5269\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25959\
        );

    \I__5268\ : CascadeMux
    port map (
            O => \N__26000\,
            I => \N__25956\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__25999\,
            I => \N__25953\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__25994\,
            I => \N__25946\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25946\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25946\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__25985\,
            I => \N__25941\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__25982\,
            I => \N__25941\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__25977\,
            I => \N__25934\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__25974\,
            I => \N__25934\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__25971\,
            I => \N__25934\
        );

    \I__5258\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25931\
        );

    \I__5257\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25928\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__25962\,
            I => \N__25923\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__25959\,
            I => \N__25923\
        );

    \I__5254\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25920\
        );

    \I__5253\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25917\
        );

    \I__5252\ : Span4Mux_v
    port map (
            O => \N__25946\,
            I => \N__25912\
        );

    \I__5251\ : Span4Mux_v
    port map (
            O => \N__25941\,
            I => \N__25912\
        );

    \I__5250\ : Span4Mux_v
    port map (
            O => \N__25934\,
            I => \N__25905\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__25931\,
            I => \N__25905\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__25928\,
            I => \N__25905\
        );

    \I__5247\ : Span4Mux_v
    port map (
            O => \N__25923\,
            I => \N__25898\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__25920\,
            I => \N__25898\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__25917\,
            I => \N__25898\
        );

    \I__5244\ : Span4Mux_h
    port map (
            O => \N__25912\,
            I => \N__25895\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__25905\,
            I => \N__25890\
        );

    \I__5242\ : Span4Mux_v
    port map (
            O => \N__25898\,
            I => \N__25890\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__25895\,
            I => \N__25884\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__25890\,
            I => \N__25884\
        );

    \I__5239\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25881\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__25884\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__25881\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__5236\ : InMux
    port map (
            O => \N__25876\,
            I => \un1_M_this_spr_address_q_cry_3\
        );

    \I__5235\ : CascadeMux
    port map (
            O => \N__25873\,
            I => \N__25870\
        );

    \I__5234\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25861\
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__25869\,
            I => \N__25858\
        );

    \I__5232\ : CascadeMux
    port map (
            O => \N__25868\,
            I => \N__25854\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__25867\,
            I => \N__25850\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__25866\,
            I => \N__25847\
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__25865\,
            I => \N__25844\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__25864\,
            I => \N__25837\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__25861\,
            I => \N__25833\
        );

    \I__5226\ : InMux
    port map (
            O => \N__25858\,
            I => \N__25830\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__25857\,
            I => \N__25827\
        );

    \I__5224\ : InMux
    port map (
            O => \N__25854\,
            I => \N__25824\
        );

    \I__5223\ : CascadeMux
    port map (
            O => \N__25853\,
            I => \N__25821\
        );

    \I__5222\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25818\
        );

    \I__5221\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25815\
        );

    \I__5220\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25812\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__25843\,
            I => \N__25809\
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__25842\,
            I => \N__25806\
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__25841\,
            I => \N__25803\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__25840\,
            I => \N__25800\
        );

    \I__5215\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25797\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__25836\,
            I => \N__25794\
        );

    \I__5213\ : Span4Mux_v
    port map (
            O => \N__25833\,
            I => \N__25787\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__25830\,
            I => \N__25787\
        );

    \I__5211\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25784\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__25824\,
            I => \N__25781\
        );

    \I__5209\ : InMux
    port map (
            O => \N__25821\,
            I => \N__25778\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__25818\,
            I => \N__25775\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__25815\,
            I => \N__25770\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__25812\,
            I => \N__25770\
        );

    \I__5205\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25767\
        );

    \I__5204\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25764\
        );

    \I__5203\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25761\
        );

    \I__5202\ : InMux
    port map (
            O => \N__25800\,
            I => \N__25758\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__25797\,
            I => \N__25755\
        );

    \I__5200\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25752\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__25793\,
            I => \N__25749\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__25792\,
            I => \N__25746\
        );

    \I__5197\ : Span4Mux_v
    port map (
            O => \N__25787\,
            I => \N__25743\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__25784\,
            I => \N__25736\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__25781\,
            I => \N__25736\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__25778\,
            I => \N__25736\
        );

    \I__5193\ : Span4Mux_s3_v
    port map (
            O => \N__25775\,
            I => \N__25733\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__25770\,
            I => \N__25728\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__25767\,
            I => \N__25728\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__25764\,
            I => \N__25723\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__25761\,
            I => \N__25723\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25720\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__25755\,
            I => \N__25717\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25714\
        );

    \I__5185\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25711\
        );

    \I__5184\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25708\
        );

    \I__5183\ : Span4Mux_v
    port map (
            O => \N__25743\,
            I => \N__25703\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__25736\,
            I => \N__25703\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__25733\,
            I => \N__25698\
        );

    \I__5180\ : Span4Mux_h
    port map (
            O => \N__25728\,
            I => \N__25698\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__25723\,
            I => \N__25693\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__25720\,
            I => \N__25693\
        );

    \I__5177\ : Span4Mux_v
    port map (
            O => \N__25717\,
            I => \N__25688\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__25714\,
            I => \N__25688\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__25711\,
            I => \N__25684\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__25708\,
            I => \N__25679\
        );

    \I__5173\ : Sp12to4
    port map (
            O => \N__25703\,
            I => \N__25679\
        );

    \I__5172\ : Sp12to4
    port map (
            O => \N__25698\,
            I => \N__25676\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__25693\,
            I => \N__25673\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__25688\,
            I => \N__25670\
        );

    \I__5169\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25667\
        );

    \I__5168\ : Span12Mux_h
    port map (
            O => \N__25684\,
            I => \N__25662\
        );

    \I__5167\ : Span12Mux_h
    port map (
            O => \N__25679\,
            I => \N__25662\
        );

    \I__5166\ : Span12Mux_v
    port map (
            O => \N__25676\,
            I => \N__25659\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__25673\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__25670\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__25667\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5162\ : Odrv12
    port map (
            O => \N__25662\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5161\ : Odrv12
    port map (
            O => \N__25659\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5160\ : InMux
    port map (
            O => \N__25648\,
            I => \un1_M_this_spr_address_q_cry_4\
        );

    \I__5159\ : CascadeMux
    port map (
            O => \N__25645\,
            I => \N__25642\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25634\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__25641\,
            I => \N__25631\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__25640\,
            I => \N__25627\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__25639\,
            I => \N__25623\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__25638\,
            I => \N__25620\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__25637\,
            I => \N__25615\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__25634\,
            I => \N__25611\
        );

    \I__5151\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25608\
        );

    \I__5150\ : CascadeMux
    port map (
            O => \N__25630\,
            I => \N__25605\
        );

    \I__5149\ : InMux
    port map (
            O => \N__25627\,
            I => \N__25601\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__25626\,
            I => \N__25598\
        );

    \I__5147\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25594\
        );

    \I__5146\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25591\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__25619\,
            I => \N__25588\
        );

    \I__5144\ : CascadeMux
    port map (
            O => \N__25618\,
            I => \N__25585\
        );

    \I__5143\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25581\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__25614\,
            I => \N__25578\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__25611\,
            I => \N__25574\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__25608\,
            I => \N__25571\
        );

    \I__5139\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25568\
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__25604\,
            I => \N__25565\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__25601\,
            I => \N__25562\
        );

    \I__5136\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25559\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__25597\,
            I => \N__25556\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__25594\,
            I => \N__25552\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__25591\,
            I => \N__25549\
        );

    \I__5132\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25546\
        );

    \I__5131\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25543\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__25584\,
            I => \N__25540\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__25581\,
            I => \N__25537\
        );

    \I__5128\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25534\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__25577\,
            I => \N__25531\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__25574\,
            I => \N__25526\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__25571\,
            I => \N__25526\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__25568\,
            I => \N__25523\
        );

    \I__5123\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25520\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__25562\,
            I => \N__25517\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__25559\,
            I => \N__25514\
        );

    \I__5120\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25511\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__25555\,
            I => \N__25508\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__25552\,
            I => \N__25505\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__25549\,
            I => \N__25502\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__25546\,
            I => \N__25499\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__25543\,
            I => \N__25496\
        );

    \I__5114\ : InMux
    port map (
            O => \N__25540\,
            I => \N__25493\
        );

    \I__5113\ : Span4Mux_h
    port map (
            O => \N__25537\,
            I => \N__25490\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__25534\,
            I => \N__25487\
        );

    \I__5111\ : InMux
    port map (
            O => \N__25531\,
            I => \N__25484\
        );

    \I__5110\ : Span4Mux_v
    port map (
            O => \N__25526\,
            I => \N__25479\
        );

    \I__5109\ : Span4Mux_h
    port map (
            O => \N__25523\,
            I => \N__25479\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__25520\,
            I => \N__25476\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__25517\,
            I => \N__25471\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__25514\,
            I => \N__25471\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__25511\,
            I => \N__25468\
        );

    \I__5104\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25465\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__25505\,
            I => \N__25458\
        );

    \I__5102\ : Span4Mux_v
    port map (
            O => \N__25502\,
            I => \N__25458\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__25499\,
            I => \N__25458\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__25496\,
            I => \N__25455\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__25493\,
            I => \N__25452\
        );

    \I__5098\ : Span4Mux_v
    port map (
            O => \N__25490\,
            I => \N__25447\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__25487\,
            I => \N__25447\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__25484\,
            I => \N__25444\
        );

    \I__5095\ : Span4Mux_h
    port map (
            O => \N__25479\,
            I => \N__25441\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__25476\,
            I => \N__25438\
        );

    \I__5093\ : Span4Mux_v
    port map (
            O => \N__25471\,
            I => \N__25433\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__25468\,
            I => \N__25433\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__25465\,
            I => \N__25430\
        );

    \I__5090\ : Span4Mux_h
    port map (
            O => \N__25458\,
            I => \N__25427\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__25455\,
            I => \N__25422\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__25452\,
            I => \N__25422\
        );

    \I__5087\ : Span4Mux_v
    port map (
            O => \N__25447\,
            I => \N__25417\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__25444\,
            I => \N__25417\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__25441\,
            I => \N__25408\
        );

    \I__5084\ : Span4Mux_v
    port map (
            O => \N__25438\,
            I => \N__25408\
        );

    \I__5083\ : Span4Mux_v
    port map (
            O => \N__25433\,
            I => \N__25408\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__25430\,
            I => \N__25408\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__25427\,
            I => \N__25400\
        );

    \I__5080\ : Span4Mux_h
    port map (
            O => \N__25422\,
            I => \N__25400\
        );

    \I__5079\ : Span4Mux_h
    port map (
            O => \N__25417\,
            I => \N__25400\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__25408\,
            I => \N__25397\
        );

    \I__5077\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25394\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__25400\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__25397\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__25394\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__5073\ : InMux
    port map (
            O => \N__25387\,
            I => \un1_M_this_spr_address_q_cry_5\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__25384\,
            I => \N__25381\
        );

    \I__5071\ : CascadeBuf
    port map (
            O => \N__25381\,
            I => \N__25378\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__25378\,
            I => \N__25374\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__25377\,
            I => \N__25371\
        );

    \I__5068\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25368\
        );

    \I__5067\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25363\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__25368\,
            I => \N__25360\
        );

    \I__5065\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25357\
        );

    \I__5064\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25354\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__25363\,
            I => \N__25351\
        );

    \I__5062\ : Span12Mux_h
    port map (
            O => \N__25360\,
            I => \N__25348\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__25357\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__25354\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__25351\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__5058\ : Odrv12
    port map (
            O => \N__25348\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__5057\ : InMux
    port map (
            O => \N__25339\,
            I => \N__25336\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__25336\,
            I => \N__25333\
        );

    \I__5055\ : Span4Mux_v
    port map (
            O => \N__25333\,
            I => \N__25330\
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__25330\,
            I => \M_this_data_tmp_qZ0Z_13\
        );

    \I__5053\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25324\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__25324\,
            I => \N__25321\
        );

    \I__5051\ : Span4Mux_v
    port map (
            O => \N__25321\,
            I => \N__25318\
        );

    \I__5050\ : Span4Mux_h
    port map (
            O => \N__25318\,
            I => \N__25315\
        );

    \I__5049\ : Odrv4
    port map (
            O => \N__25315\,
            I => \M_this_oam_ram_write_data_13\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__25312\,
            I => \N__25309\
        );

    \I__5047\ : CascadeBuf
    port map (
            O => \N__25309\,
            I => \N__25306\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__25306\,
            I => \N__25303\
        );

    \I__5045\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25300\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__25300\,
            I => \N__25297\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__25297\,
            I => \N__25291\
        );

    \I__5042\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25288\
        );

    \I__5041\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25285\
        );

    \I__5040\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25282\
        );

    \I__5039\ : Span4Mux_h
    port map (
            O => \N__25291\,
            I => \N__25279\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__25288\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__25285\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__25282\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__25279\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__25270\,
            I => \N__25267\
        );

    \I__5033\ : CascadeBuf
    port map (
            O => \N__25267\,
            I => \N__25264\
        );

    \I__5032\ : CascadeMux
    port map (
            O => \N__25264\,
            I => \N__25261\
        );

    \I__5031\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25258\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25255\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__25255\,
            I => \N__25251\
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__25254\,
            I => \N__25248\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__25251\,
            I => \N__25244\
        );

    \I__5026\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25241\
        );

    \I__5025\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25238\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__25244\,
            I => \N__25235\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__25241\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__25238\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5021\ : Odrv4
    port map (
            O => \N__25235\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5020\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25224\
        );

    \I__5019\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25221\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__25224\,
            I => \N__25215\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__25221\,
            I => \N__25215\
        );

    \I__5016\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25212\
        );

    \I__5015\ : Sp12to4
    port map (
            O => \N__25215\,
            I => \N__25207\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__25212\,
            I => \N__25207\
        );

    \I__5013\ : Odrv12
    port map (
            O => \N__25207\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__5012\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25198\
        );

    \I__5011\ : InMux
    port map (
            O => \N__25203\,
            I => \N__25198\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__25198\,
            I => \un1_M_this_oam_address_q_c4\
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__25195\,
            I => \N__25192\
        );

    \I__5008\ : CascadeBuf
    port map (
            O => \N__25192\,
            I => \N__25189\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__25189\,
            I => \N__25186\
        );

    \I__5006\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25183\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__25183\,
            I => \N__25180\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__25180\,
            I => \N__25175\
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__25179\,
            I => \N__25172\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25169\
        );

    \I__5001\ : Span4Mux_h
    port map (
            O => \N__25175\,
            I => \N__25166\
        );

    \I__5000\ : InMux
    port map (
            O => \N__25172\,
            I => \N__25163\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__25169\,
            I => \N__25158\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__25166\,
            I => \N__25158\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25163\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__25158\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__4995\ : CascadeMux
    port map (
            O => \N__25153\,
            I => \un1_M_this_oam_address_q_c4_cascade_\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__25150\,
            I => \N__25147\
        );

    \I__4993\ : CascadeBuf
    port map (
            O => \N__25147\,
            I => \N__25144\
        );

    \I__4992\ : CascadeMux
    port map (
            O => \N__25144\,
            I => \N__25141\
        );

    \I__4991\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25138\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__25138\,
            I => \N__25135\
        );

    \I__4989\ : Span4Mux_v
    port map (
            O => \N__25135\,
            I => \N__25132\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__4987\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25121\
        );

    \I__4986\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25121\
        );

    \I__4985\ : InMux
    port map (
            O => \N__25129\,
            I => \N__25118\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__25126\,
            I => \N__25115\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__25121\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__25118\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__25115\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__4980\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25104\
        );

    \I__4979\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25101\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__25104\,
            I => \un1_M_this_oam_address_q_c6\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__25101\,
            I => \un1_M_this_oam_address_q_c6\
        );

    \I__4976\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25086\
        );

    \I__4975\ : InMux
    port map (
            O => \N__25095\,
            I => \N__25086\
        );

    \I__4974\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25081\
        );

    \I__4973\ : InMux
    port map (
            O => \N__25093\,
            I => \N__25081\
        );

    \I__4972\ : InMux
    port map (
            O => \N__25092\,
            I => \N__25078\
        );

    \I__4971\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25075\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__25086\,
            I => \this_ppu.N_268_i_0_0\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__25081\,
            I => \this_ppu.N_268_i_0_0\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__25078\,
            I => \this_ppu.N_268_i_0_0\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__25075\,
            I => \this_ppu.N_268_i_0_0\
        );

    \I__4966\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25052\
        );

    \I__4965\ : InMux
    port map (
            O => \N__25065\,
            I => \N__25052\
        );

    \I__4964\ : InMux
    port map (
            O => \N__25064\,
            I => \N__25052\
        );

    \I__4963\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25052\
        );

    \I__4962\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25049\
        );

    \I__4961\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25046\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__25052\,
            I => \this_ppu.N_1323_0\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__25049\,
            I => \this_ppu.N_1323_0\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__25046\,
            I => \this_ppu.N_1323_0\
        );

    \I__4957\ : InMux
    port map (
            O => \N__25039\,
            I => \N__25035\
        );

    \I__4956\ : InMux
    port map (
            O => \N__25038\,
            I => \N__25031\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__25035\,
            I => \N__25028\
        );

    \I__4954\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25025\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__25031\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__4952\ : Odrv4
    port map (
            O => \N__25028\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__25025\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__25018\,
            I => \N__25015\
        );

    \I__4949\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25007\
        );

    \I__4948\ : CascadeMux
    port map (
            O => \N__25014\,
            I => \N__25003\
        );

    \I__4947\ : InMux
    port map (
            O => \N__25013\,
            I => \N__24998\
        );

    \I__4946\ : InMux
    port map (
            O => \N__25012\,
            I => \N__24998\
        );

    \I__4945\ : InMux
    port map (
            O => \N__25011\,
            I => \N__24995\
        );

    \I__4944\ : CascadeMux
    port map (
            O => \N__25010\,
            I => \N__24990\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__25007\,
            I => \N__24987\
        );

    \I__4942\ : InMux
    port map (
            O => \N__25006\,
            I => \N__24984\
        );

    \I__4941\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24981\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__24998\,
            I => \N__24976\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__24995\,
            I => \N__24976\
        );

    \I__4938\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24969\
        );

    \I__4937\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24969\
        );

    \I__4936\ : InMux
    port map (
            O => \N__24990\,
            I => \N__24969\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__24987\,
            I => \N__24966\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__24984\,
            I => \N__24963\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__24981\,
            I => \N__24956\
        );

    \I__4932\ : Sp12to4
    port map (
            O => \N__24976\,
            I => \N__24956\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__24969\,
            I => \N__24956\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__24966\,
            I => \N_611\
        );

    \I__4929\ : Odrv12
    port map (
            O => \N__24963\,
            I => \N_611\
        );

    \I__4928\ : Odrv12
    port map (
            O => \N__24956\,
            I => \N_611\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__24949\,
            I => \N__24946\
        );

    \I__4926\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__24943\,
            I => \N__24940\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__24940\,
            I => \M_this_data_count_q_s_13\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__4922\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24930\
        );

    \I__4921\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24927\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__24930\,
            I => \N__24924\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24919\
        );

    \I__4918\ : Span4Mux_h
    port map (
            O => \N__24924\,
            I => \N__24919\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__24919\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__4916\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24913\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__24913\,
            I => \M_this_data_count_q_s_8\
        );

    \I__4914\ : CascadeMux
    port map (
            O => \N__24910\,
            I => \N__24905\
        );

    \I__4913\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24889\
        );

    \I__4912\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24889\
        );

    \I__4911\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24889\
        );

    \I__4910\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24889\
        );

    \I__4909\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24886\
        );

    \I__4908\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24877\
        );

    \I__4907\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24877\
        );

    \I__4906\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24877\
        );

    \I__4905\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24877\
        );

    \I__4904\ : InMux
    port map (
            O => \N__24898\,
            I => \N__24870\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__24889\,
            I => \N__24865\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__24886\,
            I => \N__24865\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24862\
        );

    \I__4900\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24853\
        );

    \I__4899\ : InMux
    port map (
            O => \N__24875\,
            I => \N__24853\
        );

    \I__4898\ : InMux
    port map (
            O => \N__24874\,
            I => \N__24853\
        );

    \I__4897\ : InMux
    port map (
            O => \N__24873\,
            I => \N__24853\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__24870\,
            I => \N__24850\
        );

    \I__4895\ : Span4Mux_v
    port map (
            O => \N__24865\,
            I => \N__24847\
        );

    \I__4894\ : Span4Mux_h
    port map (
            O => \N__24862\,
            I => \N__24842\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__24853\,
            I => \N__24842\
        );

    \I__4892\ : Odrv12
    port map (
            O => \N__24850\,
            I => \N_660_i\
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__24847\,
            I => \N_660_i\
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__24842\,
            I => \N_660_i\
        );

    \I__4889\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24831\
        );

    \I__4888\ : InMux
    port map (
            O => \N__24834\,
            I => \N__24828\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__24831\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__24828\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__4885\ : CEMux
    port map (
            O => \N__24823\,
            I => \N__24820\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__24820\,
            I => \N__24816\
        );

    \I__4883\ : CEMux
    port map (
            O => \N__24819\,
            I => \N__24812\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__24816\,
            I => \N__24808\
        );

    \I__4881\ : CEMux
    port map (
            O => \N__24815\,
            I => \N__24805\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__24812\,
            I => \N__24801\
        );

    \I__4879\ : CEMux
    port map (
            O => \N__24811\,
            I => \N__24798\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__24808\,
            I => \N__24793\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__24805\,
            I => \N__24793\
        );

    \I__4876\ : CEMux
    port map (
            O => \N__24804\,
            I => \N__24790\
        );

    \I__4875\ : Span4Mux_h
    port map (
            O => \N__24801\,
            I => \N__24785\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__24798\,
            I => \N__24785\
        );

    \I__4873\ : Span4Mux_v
    port map (
            O => \N__24793\,
            I => \N__24782\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__24790\,
            I => \N__24779\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__24785\,
            I => \N__24776\
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__24782\,
            I => \N_257\
        );

    \I__4869\ : Odrv12
    port map (
            O => \N__24779\,
            I => \N_257\
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__24776\,
            I => \N_257\
        );

    \I__4867\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__24766\,
            I => \N__24761\
        );

    \I__4865\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24758\
        );

    \I__4864\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24754\
        );

    \I__4863\ : Span4Mux_v
    port map (
            O => \N__24761\,
            I => \N__24749\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__24758\,
            I => \N__24749\
        );

    \I__4861\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24746\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__24754\,
            I => \N__24743\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__24749\,
            I => \N__24740\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__24746\,
            I => \N__24737\
        );

    \I__4857\ : Sp12to4
    port map (
            O => \N__24743\,
            I => \N__24734\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__24740\,
            I => \N__24731\
        );

    \I__4855\ : Span4Mux_h
    port map (
            O => \N__24737\,
            I => \N__24726\
        );

    \I__4854\ : Span12Mux_v
    port map (
            O => \N__24734\,
            I => \N__24723\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__24731\,
            I => \N__24720\
        );

    \I__4852\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24715\
        );

    \I__4851\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24715\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__24726\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4849\ : Odrv12
    port map (
            O => \N__24723\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__24720\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__24715\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__4846\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24703\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__24703\,
            I => \N__24695\
        );

    \I__4844\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24692\
        );

    \I__4843\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24689\
        );

    \I__4842\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24684\
        );

    \I__4841\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24684\
        );

    \I__4840\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24681\
        );

    \I__4839\ : Span4Mux_v
    port map (
            O => \N__24695\,
            I => \N__24678\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__24692\,
            I => \N__24675\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__24689\,
            I => \N__24672\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__24684\,
            I => \N__24669\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__24681\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__24678\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4833\ : Odrv12
    port map (
            O => \N__24675\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__24672\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4831\ : Odrv12
    port map (
            O => \N__24669\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4830\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24652\
        );

    \I__4829\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24649\
        );

    \I__4828\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24646\
        );

    \I__4827\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24640\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__24652\,
            I => \N__24635\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__24649\,
            I => \N__24635\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24632\
        );

    \I__4823\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24627\
        );

    \I__4822\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24627\
        );

    \I__4821\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24624\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24619\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__24635\,
            I => \N__24619\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__24632\,
            I => \N__24614\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__24627\,
            I => \N__24614\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__24624\,
            I => \N__24607\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__24619\,
            I => \N__24607\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__24614\,
            I => \N__24607\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__24607\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__4812\ : CascadeMux
    port map (
            O => \N__24604\,
            I => \N__24599\
        );

    \I__4811\ : CascadeMux
    port map (
            O => \N__24603\,
            I => \N__24596\
        );

    \I__4810\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24592\
        );

    \I__4809\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24589\
        );

    \I__4808\ : InMux
    port map (
            O => \N__24596\,
            I => \N__24586\
        );

    \I__4807\ : CascadeMux
    port map (
            O => \N__24595\,
            I => \N__24583\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__24592\,
            I => \N__24575\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__24589\,
            I => \N__24575\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__24586\,
            I => \N__24575\
        );

    \I__4803\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24572\
        );

    \I__4802\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24568\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__24575\,
            I => \N__24565\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__24572\,
            I => \N__24562\
        );

    \I__4799\ : InMux
    port map (
            O => \N__24571\,
            I => \N__24559\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24556\
        );

    \I__4797\ : Span4Mux_h
    port map (
            O => \N__24565\,
            I => \N__24553\
        );

    \I__4796\ : Sp12to4
    port map (
            O => \N__24562\,
            I => \N__24548\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__24559\,
            I => \N__24548\
        );

    \I__4794\ : Odrv12
    port map (
            O => \N__24556\,
            I => \N_314_1\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__24553\,
            I => \N_314_1\
        );

    \I__4792\ : Odrv12
    port map (
            O => \N__24548\,
            I => \N_314_1\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__24541\,
            I => \N__24537\
        );

    \I__4790\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24532\
        );

    \I__4789\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24532\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__24532\,
            I => \N__24527\
        );

    \I__4787\ : InMux
    port map (
            O => \N__24531\,
            I => \N__24524\
        );

    \I__4786\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24521\
        );

    \I__4785\ : Span4Mux_v
    port map (
            O => \N__24527\,
            I => \N__24518\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__24524\,
            I => \N__24515\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__24521\,
            I => \N__24512\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__24518\,
            I => \N__24508\
        );

    \I__4781\ : Span4Mux_v
    port map (
            O => \N__24515\,
            I => \N__24503\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__24512\,
            I => \N__24503\
        );

    \I__4779\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24500\
        );

    \I__4778\ : Sp12to4
    port map (
            O => \N__24508\,
            I => \N__24493\
        );

    \I__4777\ : Sp12to4
    port map (
            O => \N__24503\,
            I => \N__24493\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__24500\,
            I => \N__24493\
        );

    \I__4775\ : Span12Mux_h
    port map (
            O => \N__24493\,
            I => \N__24490\
        );

    \I__4774\ : Odrv12
    port map (
            O => \N__24490\,
            I => port_enb_c
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \N__24484\
        );

    \I__4772\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__4770\ : Span4Mux_v
    port map (
            O => \N__24478\,
            I => \N__24471\
        );

    \I__4769\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24468\
        );

    \I__4768\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24461\
        );

    \I__4767\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24461\
        );

    \I__4766\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24461\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__24471\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__24468\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__24461\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4762\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24451\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__24451\,
            I => \N__24446\
        );

    \I__4760\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24443\
        );

    \I__4759\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24438\
        );

    \I__4758\ : Span4Mux_v
    port map (
            O => \N__24446\,
            I => \N__24433\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__24443\,
            I => \N__24433\
        );

    \I__4756\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24428\
        );

    \I__4755\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24428\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__24438\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__24433\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__24428\,
            I => \M_this_delay_clk_out_0\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__24421\,
            I => \N_309_0_cascade_\
        );

    \I__4750\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24415\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__24415\,
            I => \M_this_data_count_q_cry_0_THRU_CO\
        );

    \I__4748\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24407\
        );

    \I__4747\ : InMux
    port map (
            O => \N__24411\,
            I => \N__24404\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24401\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__24407\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__24404\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__24401\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__4742\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24391\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__24391\,
            I => \M_this_data_count_q_cry_5_THRU_CO\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__24388\,
            I => \N__24383\
        );

    \I__4739\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24380\
        );

    \I__4738\ : InMux
    port map (
            O => \N__24386\,
            I => \N__24377\
        );

    \I__4737\ : InMux
    port map (
            O => \N__24383\,
            I => \N__24374\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__24380\,
            I => \N__24371\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__24377\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__24374\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4733\ : Odrv4
    port map (
            O => \N__24371\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__4732\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24361\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__24361\,
            I => \M_this_data_count_q_cry_6_THRU_CO\
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__24358\,
            I => \N__24353\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__24357\,
            I => \N__24350\
        );

    \I__4728\ : InMux
    port map (
            O => \N__24356\,
            I => \N__24347\
        );

    \I__4727\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24344\
        );

    \I__4726\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24341\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__24347\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__24344\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__24341\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__24334\,
            I => \N__24331\
        );

    \I__4721\ : CascadeBuf
    port map (
            O => \N__24331\,
            I => \N__24328\
        );

    \I__4720\ : CascadeMux
    port map (
            O => \N__24328\,
            I => \N__24325\
        );

    \I__4719\ : InMux
    port map (
            O => \N__24325\,
            I => \N__24322\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__24322\,
            I => \N__24319\
        );

    \I__4717\ : Sp12to4
    port map (
            O => \N__24319\,
            I => \N__24314\
        );

    \I__4716\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24311\
        );

    \I__4715\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24308\
        );

    \I__4714\ : Span12Mux_h
    port map (
            O => \N__24314\,
            I => \N__24305\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__24311\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__24308\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__4711\ : Odrv12
    port map (
            O => \N__24305\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__24298\,
            I => \N__24295\
        );

    \I__4709\ : CascadeBuf
    port map (
            O => \N__24295\,
            I => \N__24292\
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__24292\,
            I => \N__24289\
        );

    \I__4707\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24286\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24282\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__24285\,
            I => \N__24279\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__24282\,
            I => \N__24276\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24273\
        );

    \I__4702\ : Span4Mux_h
    port map (
            O => \N__24276\,
            I => \N__24270\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__24273\,
            I => \N__24265\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__24270\,
            I => \N__24265\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__24265\,
            I => \M_this_oam_address_qZ0Z_7\
        );

    \I__4698\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24252\
        );

    \I__4697\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24249\
        );

    \I__4696\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24244\
        );

    \I__4695\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24244\
        );

    \I__4694\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24235\
        );

    \I__4693\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24235\
        );

    \I__4692\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24235\
        );

    \I__4691\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24235\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__24252\,
            I => \N__24230\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__24249\,
            I => \N__24223\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__24244\,
            I => \N__24223\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__24235\,
            I => \N__24223\
        );

    \I__4686\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24218\
        );

    \I__4685\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24218\
        );

    \I__4684\ : Span4Mux_v
    port map (
            O => \N__24230\,
            I => \N__24215\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__24223\,
            I => \N__24210\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24210\
        );

    \I__4681\ : Sp12to4
    port map (
            O => \N__24215\,
            I => \N__24207\
        );

    \I__4680\ : Span4Mux_v
    port map (
            O => \N__24210\,
            I => \N__24204\
        );

    \I__4679\ : Span12Mux_h
    port map (
            O => \N__24207\,
            I => \N__24201\
        );

    \I__4678\ : Span4Mux_v
    port map (
            O => \N__24204\,
            I => \N__24198\
        );

    \I__4677\ : Odrv12
    port map (
            O => \N__24201\,
            I => rst_n_c
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__24198\,
            I => rst_n_c
        );

    \I__4675\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24190\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__24190\,
            I => \this_reset_cond.M_stage_qZ0Z_6\
        );

    \I__4673\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24184\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__24184\,
            I => \this_reset_cond.M_stage_qZ0Z_7\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__24181\,
            I => \this_ppu.N_760_0_cascade_\
        );

    \I__4670\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24175\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__24175\,
            I => \N__24168\
        );

    \I__4668\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24165\
        );

    \I__4667\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24158\
        );

    \I__4666\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24158\
        );

    \I__4665\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24158\
        );

    \I__4664\ : Span4Mux_v
    port map (
            O => \N__24168\,
            I => \N__24155\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__24165\,
            I => \N__24150\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__24158\,
            I => \N__24150\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__24155\,
            I => \N__24147\
        );

    \I__4660\ : Span12Mux_h
    port map (
            O => \N__24150\,
            I => \N__24144\
        );

    \I__4659\ : Span4Mux_h
    port map (
            O => \N__24147\,
            I => \N__24141\
        );

    \I__4658\ : Span12Mux_v
    port map (
            O => \N__24144\,
            I => \N__24138\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__24141\,
            I => \this_ppu.N_762_0\
        );

    \I__4656\ : Odrv12
    port map (
            O => \N__24138\,
            I => \this_ppu.N_762_0\
        );

    \I__4655\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24130\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24127\
        );

    \I__4653\ : Span4Mux_h
    port map (
            O => \N__24127\,
            I => \N__24121\
        );

    \I__4652\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24118\
        );

    \I__4651\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24115\
        );

    \I__4650\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24112\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__24121\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__24118\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__24115\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__24112\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4645\ : CascadeMux
    port map (
            O => \N__24103\,
            I => \N__24100\
        );

    \I__4644\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24095\
        );

    \I__4643\ : CascadeMux
    port map (
            O => \N__24099\,
            I => \N__24092\
        );

    \I__4642\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24089\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__24095\,
            I => \N__24086\
        );

    \I__4640\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24082\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24079\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__24086\,
            I => \N__24076\
        );

    \I__4637\ : InMux
    port map (
            O => \N__24085\,
            I => \N__24073\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__24082\,
            I => \N__24070\
        );

    \I__4635\ : Sp12to4
    port map (
            O => \N__24079\,
            I => \N__24067\
        );

    \I__4634\ : Span4Mux_v
    port map (
            O => \N__24076\,
            I => \N__24063\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__24073\,
            I => \N__24058\
        );

    \I__4632\ : Span4Mux_h
    port map (
            O => \N__24070\,
            I => \N__24058\
        );

    \I__4631\ : Span12Mux_v
    port map (
            O => \N__24067\,
            I => \N__24055\
        );

    \I__4630\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24052\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__24063\,
            I => \this_ppu.M_last_q\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__24058\,
            I => \this_ppu.M_last_q\
        );

    \I__4627\ : Odrv12
    port map (
            O => \N__24055\,
            I => \this_ppu.M_last_q\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__24052\,
            I => \this_ppu.M_last_q\
        );

    \I__4625\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24040\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__24040\,
            I => \N__24035\
        );

    \I__4623\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24032\
        );

    \I__4622\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24028\
        );

    \I__4621\ : Span4Mux_h
    port map (
            O => \N__24035\,
            I => \N__24023\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__24032\,
            I => \N__24023\
        );

    \I__4619\ : InMux
    port map (
            O => \N__24031\,
            I => \N__24020\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__24028\,
            I => \N__24017\
        );

    \I__4617\ : Span4Mux_v
    port map (
            O => \N__24023\,
            I => \N__24014\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__24009\
        );

    \I__4615\ : Span4Mux_h
    port map (
            O => \N__24017\,
            I => \N__24009\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__24014\,
            I => \N__24006\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__24009\,
            I => \this_ppu.N_5_4\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__24006\,
            I => \this_ppu.N_5_4\
        );

    \I__4611\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23998\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__23998\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__23995\,
            I => \this_ppu.N_268_i_0_0_cascade_\
        );

    \I__4608\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23987\
        );

    \I__4607\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23984\
        );

    \I__4606\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23981\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__23987\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__23984\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__23981\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__4602\ : IoInMux
    port map (
            O => \N__23974\,
            I => \N__23970\
        );

    \I__4601\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23967\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__23970\,
            I => \N__23964\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__23967\,
            I => \N__23961\
        );

    \I__4598\ : IoSpan4Mux
    port map (
            O => \N__23964\,
            I => \N__23950\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__23961\,
            I => \N__23947\
        );

    \I__4596\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23938\
        );

    \I__4595\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23938\
        );

    \I__4594\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23938\
        );

    \I__4593\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23938\
        );

    \I__4592\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23933\
        );

    \I__4591\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23933\
        );

    \I__4590\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23930\
        );

    \I__4589\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23927\
        );

    \I__4588\ : Span4Mux_s1_h
    port map (
            O => \N__23950\,
            I => \N__23924\
        );

    \I__4587\ : Sp12to4
    port map (
            O => \N__23947\,
            I => \N__23919\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__23938\,
            I => \N__23919\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__23933\,
            I => \N__23916\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23913\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__23927\,
            I => \N__23910\
        );

    \I__4582\ : Sp12to4
    port map (
            O => \N__23924\,
            I => \N__23907\
        );

    \I__4581\ : Span12Mux_h
    port map (
            O => \N__23919\,
            I => \N__23904\
        );

    \I__4580\ : Span12Mux_s11_h
    port map (
            O => \N__23916\,
            I => \N__23899\
        );

    \I__4579\ : Span12Mux_v
    port map (
            O => \N__23913\,
            I => \N__23899\
        );

    \I__4578\ : Span12Mux_v
    port map (
            O => \N__23910\,
            I => \N__23894\
        );

    \I__4577\ : Span12Mux_h
    port map (
            O => \N__23907\,
            I => \N__23894\
        );

    \I__4576\ : Odrv12
    port map (
            O => \N__23904\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4575\ : Odrv12
    port map (
            O => \N__23899\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4574\ : Odrv12
    port map (
            O => \N__23894\,
            I => \M_this_reset_cond_out_0\
        );

    \I__4573\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23884\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__23884\,
            I => \N__23881\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__23881\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__23878\,
            I => \this_ppu.N_1323_0_cascade_\
        );

    \I__4569\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23870\
        );

    \I__4568\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23867\
        );

    \I__4567\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23864\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__23870\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__23867\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__23864\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__4563\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23853\
        );

    \I__4562\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23850\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__23853\,
            I => \N__23845\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__23850\,
            I => \N__23845\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__23845\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__4558\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__23839\,
            I => \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_3\
        );

    \I__4556\ : InMux
    port map (
            O => \N__23836\,
            I => \bfn_17_19_0_\
        );

    \I__4555\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__23827\,
            I => \M_this_data_count_q_cry_8_THRU_CO\
        );

    \I__4552\ : InMux
    port map (
            O => \N__23824\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__4551\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23817\
        );

    \I__4550\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23814\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__23817\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__23814\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__4547\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23806\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__23806\,
            I => \M_this_data_count_q_s_10\
        );

    \I__4545\ : InMux
    port map (
            O => \N__23803\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__23800\,
            I => \N__23797\
        );

    \I__4543\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23792\
        );

    \I__4542\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23787\
        );

    \I__4541\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23787\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__23792\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__23787\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__4538\ : CascadeMux
    port map (
            O => \N__23782\,
            I => \N__23779\
        );

    \I__4537\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23776\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__23776\,
            I => \M_this_data_count_q_cry_10_THRU_CO\
        );

    \I__4535\ : InMux
    port map (
            O => \N__23773\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__23770\,
            I => \N__23764\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__23769\,
            I => \N__23760\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__23768\,
            I => \N__23756\
        );

    \I__4531\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23736\
        );

    \I__4530\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23736\
        );

    \I__4529\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23736\
        );

    \I__4528\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23736\
        );

    \I__4527\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23736\
        );

    \I__4526\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23736\
        );

    \I__4525\ : CascadeMux
    port map (
            O => \N__23755\,
            I => \N__23732\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__23754\,
            I => \N__23729\
        );

    \I__4523\ : SRMux
    port map (
            O => \N__23753\,
            I => \N__23726\
        );

    \I__4522\ : SRMux
    port map (
            O => \N__23752\,
            I => \N__23723\
        );

    \I__4521\ : SRMux
    port map (
            O => \N__23751\,
            I => \N__23720\
        );

    \I__4520\ : IoInMux
    port map (
            O => \N__23750\,
            I => \N__23714\
        );

    \I__4519\ : CascadeMux
    port map (
            O => \N__23749\,
            I => \N__23709\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23705\
        );

    \I__4517\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23698\
        );

    \I__4516\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23698\
        );

    \I__4515\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23698\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23726\,
            I => \N__23689\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__23723\,
            I => \N__23689\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23686\
        );

    \I__4511\ : SRMux
    port map (
            O => \N__23719\,
            I => \N__23683\
        );

    \I__4510\ : SRMux
    port map (
            O => \N__23718\,
            I => \N__23680\
        );

    \I__4509\ : SRMux
    port map (
            O => \N__23717\,
            I => \N__23677\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__23714\,
            I => \N__23671\
        );

    \I__4507\ : SRMux
    port map (
            O => \N__23713\,
            I => \N__23668\
        );

    \I__4506\ : SRMux
    port map (
            O => \N__23712\,
            I => \N__23664\
        );

    \I__4505\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23657\
        );

    \I__4504\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23657\
        );

    \I__4503\ : Span4Mux_h
    port map (
            O => \N__23705\,
            I => \N__23652\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__23698\,
            I => \N__23652\
        );

    \I__4501\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23649\
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__23696\,
            I => \N__23645\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__23695\,
            I => \N__23641\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__23694\,
            I => \N__23637\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__23689\,
            I => \N__23627\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__23686\,
            I => \N__23627\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__23683\,
            I => \N__23627\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__23680\,
            I => \N__23627\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23677\,
            I => \N__23624\
        );

    \I__4492\ : SRMux
    port map (
            O => \N__23676\,
            I => \N__23621\
        );

    \I__4491\ : SRMux
    port map (
            O => \N__23675\,
            I => \N__23618\
        );

    \I__4490\ : SRMux
    port map (
            O => \N__23674\,
            I => \N__23615\
        );

    \I__4489\ : IoSpan4Mux
    port map (
            O => \N__23671\,
            I => \N__23610\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23607\
        );

    \I__4487\ : SRMux
    port map (
            O => \N__23667\,
            I => \N__23604\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__23664\,
            I => \N__23601\
        );

    \I__4485\ : SRMux
    port map (
            O => \N__23663\,
            I => \N__23598\
        );

    \I__4484\ : SRMux
    port map (
            O => \N__23662\,
            I => \N__23592\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23588\
        );

    \I__4482\ : Span4Mux_v
    port map (
            O => \N__23652\,
            I => \N__23583\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__23649\,
            I => \N__23583\
        );

    \I__4480\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23570\
        );

    \I__4479\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23570\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23644\,
            I => \N__23570\
        );

    \I__4477\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23570\
        );

    \I__4476\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23570\
        );

    \I__4475\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23570\
        );

    \I__4474\ : IoInMux
    port map (
            O => \N__23636\,
            I => \N__23567\
        );

    \I__4473\ : Span4Mux_v
    port map (
            O => \N__23627\,
            I => \N__23558\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__23624\,
            I => \N__23558\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__23621\,
            I => \N__23558\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__23618\,
            I => \N__23558\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23555\
        );

    \I__4468\ : SRMux
    port map (
            O => \N__23614\,
            I => \N__23552\
        );

    \I__4467\ : SRMux
    port map (
            O => \N__23613\,
            I => \N__23549\
        );

    \I__4466\ : Span4Mux_s3_h
    port map (
            O => \N__23610\,
            I => \N__23542\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__23607\,
            I => \N__23537\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__23604\,
            I => \N__23537\
        );

    \I__4463\ : Span4Mux_v
    port map (
            O => \N__23601\,
            I => \N__23532\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__23598\,
            I => \N__23532\
        );

    \I__4461\ : SRMux
    port map (
            O => \N__23597\,
            I => \N__23529\
        );

    \I__4460\ : SRMux
    port map (
            O => \N__23596\,
            I => \N__23526\
        );

    \I__4459\ : SRMux
    port map (
            O => \N__23595\,
            I => \N__23518\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__23592\,
            I => \N__23515\
        );

    \I__4457\ : SRMux
    port map (
            O => \N__23591\,
            I => \N__23510\
        );

    \I__4456\ : Span4Mux_v
    port map (
            O => \N__23588\,
            I => \N__23503\
        );

    \I__4455\ : Span4Mux_h
    port map (
            O => \N__23583\,
            I => \N__23503\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23503\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__23567\,
            I => \N__23500\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__23558\,
            I => \N__23491\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__23555\,
            I => \N__23491\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__23552\,
            I => \N__23491\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23491\
        );

    \I__4448\ : SRMux
    port map (
            O => \N__23548\,
            I => \N__23488\
        );

    \I__4447\ : SRMux
    port map (
            O => \N__23547\,
            I => \N__23485\
        );

    \I__4446\ : SRMux
    port map (
            O => \N__23546\,
            I => \N__23482\
        );

    \I__4445\ : SRMux
    port map (
            O => \N__23545\,
            I => \N__23478\
        );

    \I__4444\ : Span4Mux_h
    port map (
            O => \N__23542\,
            I => \N__23466\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__23537\,
            I => \N__23466\
        );

    \I__4442\ : Span4Mux_v
    port map (
            O => \N__23532\,
            I => \N__23466\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__23529\,
            I => \N__23466\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__23526\,
            I => \N__23463\
        );

    \I__4439\ : SRMux
    port map (
            O => \N__23525\,
            I => \N__23460\
        );

    \I__4438\ : SRMux
    port map (
            O => \N__23524\,
            I => \N__23457\
        );

    \I__4437\ : SRMux
    port map (
            O => \N__23523\,
            I => \N__23451\
        );

    \I__4436\ : SRMux
    port map (
            O => \N__23522\,
            I => \N__23448\
        );

    \I__4435\ : SRMux
    port map (
            O => \N__23521\,
            I => \N__23442\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__23518\,
            I => \N__23437\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__23515\,
            I => \N__23437\
        );

    \I__4432\ : SRMux
    port map (
            O => \N__23514\,
            I => \N__23434\
        );

    \I__4431\ : SRMux
    port map (
            O => \N__23513\,
            I => \N__23431\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__23510\,
            I => \N__23425\
        );

    \I__4429\ : Span4Mux_v
    port map (
            O => \N__23503\,
            I => \N__23422\
        );

    \I__4428\ : Span4Mux_s2_h
    port map (
            O => \N__23500\,
            I => \N__23419\
        );

    \I__4427\ : Span4Mux_v
    port map (
            O => \N__23491\,
            I => \N__23412\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__23488\,
            I => \N__23412\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__23485\,
            I => \N__23412\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23409\
        );

    \I__4423\ : SRMux
    port map (
            O => \N__23481\,
            I => \N__23406\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__23478\,
            I => \N__23402\
        );

    \I__4421\ : SRMux
    port map (
            O => \N__23477\,
            I => \N__23399\
        );

    \I__4420\ : SRMux
    port map (
            O => \N__23476\,
            I => \N__23396\
        );

    \I__4419\ : SRMux
    port map (
            O => \N__23475\,
            I => \N__23393\
        );

    \I__4418\ : Span4Mux_v
    port map (
            O => \N__23466\,
            I => \N__23384\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__23463\,
            I => \N__23384\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23384\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23384\
        );

    \I__4414\ : SRMux
    port map (
            O => \N__23456\,
            I => \N__23381\
        );

    \I__4413\ : SRMux
    port map (
            O => \N__23455\,
            I => \N__23378\
        );

    \I__4412\ : SRMux
    port map (
            O => \N__23454\,
            I => \N__23375\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__23451\,
            I => \N__23370\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__23448\,
            I => \N__23370\
        );

    \I__4409\ : SRMux
    port map (
            O => \N__23447\,
            I => \N__23367\
        );

    \I__4408\ : SRMux
    port map (
            O => \N__23446\,
            I => \N__23364\
        );

    \I__4407\ : SRMux
    port map (
            O => \N__23445\,
            I => \N__23360\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__23442\,
            I => \N__23351\
        );

    \I__4405\ : Sp12to4
    port map (
            O => \N__23437\,
            I => \N__23351\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__23434\,
            I => \N__23351\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N__23351\
        );

    \I__4402\ : SRMux
    port map (
            O => \N__23430\,
            I => \N__23348\
        );

    \I__4401\ : SRMux
    port map (
            O => \N__23429\,
            I => \N__23345\
        );

    \I__4400\ : SRMux
    port map (
            O => \N__23428\,
            I => \N__23342\
        );

    \I__4399\ : Span4Mux_h
    port map (
            O => \N__23425\,
            I => \N__23339\
        );

    \I__4398\ : Span4Mux_v
    port map (
            O => \N__23422\,
            I => \N__23336\
        );

    \I__4397\ : Span4Mux_h
    port map (
            O => \N__23419\,
            I => \N__23331\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__23412\,
            I => \N__23331\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__23409\,
            I => \N__23328\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__23406\,
            I => \N__23325\
        );

    \I__4393\ : SRMux
    port map (
            O => \N__23405\,
            I => \N__23322\
        );

    \I__4392\ : Span4Mux_s1_v
    port map (
            O => \N__23402\,
            I => \N__23315\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__23399\,
            I => \N__23315\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__23396\,
            I => \N__23315\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__23393\,
            I => \N__23312\
        );

    \I__4388\ : Span4Mux_v
    port map (
            O => \N__23384\,
            I => \N__23305\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23305\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23305\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__23375\,
            I => \N__23302\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__23370\,
            I => \N__23295\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23295\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__23364\,
            I => \N__23295\
        );

    \I__4381\ : SRMux
    port map (
            O => \N__23363\,
            I => \N__23292\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23289\
        );

    \I__4379\ : Span12Mux_v
    port map (
            O => \N__23351\,
            I => \N__23280\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__23348\,
            I => \N__23280\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23280\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23280\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__23339\,
            I => \N__23273\
        );

    \I__4374\ : Span4Mux_v
    port map (
            O => \N__23336\,
            I => \N__23273\
        );

    \I__4373\ : Span4Mux_h
    port map (
            O => \N__23331\,
            I => \N__23273\
        );

    \I__4372\ : Span4Mux_v
    port map (
            O => \N__23328\,
            I => \N__23268\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__23325\,
            I => \N__23268\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23263\
        );

    \I__4369\ : Sp12to4
    port map (
            O => \N__23315\,
            I => \N__23263\
        );

    \I__4368\ : Span4Mux_v
    port map (
            O => \N__23312\,
            I => \N__23258\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__23305\,
            I => \N__23258\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__23302\,
            I => \N__23251\
        );

    \I__4365\ : Span4Mux_v
    port map (
            O => \N__23295\,
            I => \N__23251\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__23292\,
            I => \N__23251\
        );

    \I__4363\ : Span4Mux_h
    port map (
            O => \N__23289\,
            I => \N__23248\
        );

    \I__4362\ : Span12Mux_v
    port map (
            O => \N__23280\,
            I => \N__23239\
        );

    \I__4361\ : Sp12to4
    port map (
            O => \N__23273\,
            I => \N__23239\
        );

    \I__4360\ : Sp12to4
    port map (
            O => \N__23268\,
            I => \N__23239\
        );

    \I__4359\ : Span12Mux_s5_v
    port map (
            O => \N__23263\,
            I => \N__23239\
        );

    \I__4358\ : Span4Mux_h
    port map (
            O => \N__23258\,
            I => \N__23234\
        );

    \I__4357\ : Span4Mux_h
    port map (
            O => \N__23251\,
            I => \N__23234\
        );

    \I__4356\ : Span4Mux_h
    port map (
            O => \N__23248\,
            I => \N__23231\
        );

    \I__4355\ : Odrv12
    port map (
            O => \N__23239\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__23234\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__23231\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__23224\,
            I => \N__23221\
        );

    \I__4351\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23216\
        );

    \I__4350\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23211\
        );

    \I__4349\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23211\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__23216\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__23211\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__4346\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23203\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__23203\,
            I => \M_this_data_count_q_cry_11_THRU_CO\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23200\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__4343\ : InMux
    port map (
            O => \N__23197\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__4342\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23189\
        );

    \I__4341\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23186\
        );

    \I__4340\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23183\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__23189\,
            I => \N__23180\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__23186\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__23183\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__23180\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__23173\,
            I => \N__23169\
        );

    \I__4334\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23163\
        );

    \I__4333\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23163\
        );

    \I__4332\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23160\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23157\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__23160\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__23157\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__23152\,
            I => \N__23149\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23144\
        );

    \I__4326\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23141\
        );

    \I__4325\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23138\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__23144\,
            I => \N__23133\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23133\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__23138\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__23133\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__4320\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23125\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__23125\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_11\
        );

    \I__4318\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23119\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__23116\,
            I => \N__23111\
        );

    \I__4315\ : InMux
    port map (
            O => \N__23115\,
            I => \N__23106\
        );

    \I__4314\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23106\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__23111\,
            I => \this_ppu.N_91\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__23106\,
            I => \this_ppu.N_91\
        );

    \I__4311\ : InMux
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__23095\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_11\
        );

    \I__4308\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23087\
        );

    \I__4307\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23082\
        );

    \I__4306\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23082\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__23087\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__23082\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__4303\ : InMux
    port map (
            O => \N__23077\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__4301\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23066\
        );

    \I__4300\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23061\
        );

    \I__4299\ : InMux
    port map (
            O => \N__23069\,
            I => \N__23061\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__23066\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__23061\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__4296\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23053\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__23053\,
            I => \M_this_data_count_q_cry_1_THRU_CO\
        );

    \I__4294\ : InMux
    port map (
            O => \N__23050\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__4293\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23042\
        );

    \I__4292\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23039\
        );

    \I__4291\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23036\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__23042\,
            I => \N__23033\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__23039\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__23036\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__23033\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__4286\ : InMux
    port map (
            O => \N__23026\,
            I => \N__23023\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__23023\,
            I => \M_this_data_count_q_cry_2_THRU_CO\
        );

    \I__4284\ : InMux
    port map (
            O => \N__23020\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__4283\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__23014\,
            I => \M_this_data_count_q_cry_3_THRU_CO\
        );

    \I__4281\ : InMux
    port map (
            O => \N__23011\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__4280\ : InMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__23005\,
            I => \M_this_data_count_q_cry_4_THRU_CO\
        );

    \I__4278\ : InMux
    port map (
            O => \N__23002\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__4277\ : InMux
    port map (
            O => \N__22999\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__4276\ : InMux
    port map (
            O => \N__22996\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__4275\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22990\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__22987\,
            I => \N__22984\
        );

    \I__4272\ : Span4Mux_h
    port map (
            O => \N__22984\,
            I => \N__22981\
        );

    \I__4271\ : Span4Mux_h
    port map (
            O => \N__22981\,
            I => \N__22978\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__22978\,
            I => \this_ppu.oam_cache.mem_5\
        );

    \I__4269\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22972\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__22972\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_5\
        );

    \I__4267\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22965\
        );

    \I__4266\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22961\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22957\
        );

    \I__4264\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22954\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__22961\,
            I => \N__22950\
        );

    \I__4262\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22947\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__22957\,
            I => \N__22942\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__22954\,
            I => \N__22939\
        );

    \I__4259\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22936\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__22950\,
            I => \N__22933\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22930\
        );

    \I__4256\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22927\
        );

    \I__4255\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22923\
        );

    \I__4254\ : Span4Mux_v
    port map (
            O => \N__22942\,
            I => \N__22918\
        );

    \I__4253\ : Span4Mux_h
    port map (
            O => \N__22939\,
            I => \N__22918\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__22936\,
            I => \N__22915\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__22933\,
            I => \N__22910\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__22930\,
            I => \N__22910\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__22927\,
            I => \N__22907\
        );

    \I__4248\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22904\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__22923\,
            I => \N__22901\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__22918\,
            I => \N__22896\
        );

    \I__4245\ : Span4Mux_h
    port map (
            O => \N__22915\,
            I => \N__22896\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__22910\,
            I => \N__22891\
        );

    \I__4243\ : Span4Mux_h
    port map (
            O => \N__22907\,
            I => \N__22891\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__22904\,
            I => \N__22888\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__22901\,
            I => \N__22885\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__22896\,
            I => \N__22882\
        );

    \I__4239\ : Span4Mux_v
    port map (
            O => \N__22891\,
            I => \N__22877\
        );

    \I__4238\ : Span4Mux_h
    port map (
            O => \N__22888\,
            I => \N__22877\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__22885\,
            I => \N__22870\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__22882\,
            I => \N__22870\
        );

    \I__4235\ : Span4Mux_h
    port map (
            O => \N__22877\,
            I => \N__22870\
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__22870\,
            I => \M_this_spr_ram_write_data_1\
        );

    \I__4233\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22853\
        );

    \I__4232\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22853\
        );

    \I__4231\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22844\
        );

    \I__4230\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22844\
        );

    \I__4229\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22844\
        );

    \I__4228\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22844\
        );

    \I__4227\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22835\
        );

    \I__4226\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22835\
        );

    \I__4225\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22835\
        );

    \I__4224\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22835\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__22853\,
            I => \N__22828\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__22844\,
            I => \N__22828\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__22835\,
            I => \N__22828\
        );

    \I__4220\ : Span4Mux_v
    port map (
            O => \N__22828\,
            I => \N__22824\
        );

    \I__4219\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22821\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__22824\,
            I => \N__22818\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22813\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__22818\,
            I => \N__22813\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__22813\,
            I => \N_609\
        );

    \I__4214\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22807\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__22807\,
            I => \this_reset_cond.M_stage_qZ0Z_5\
        );

    \I__4212\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22801\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__22801\,
            I => \this_reset_cond.M_stage_qZ0Z_3\
        );

    \I__4210\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__22795\,
            I => \this_reset_cond.M_stage_qZ0Z_4\
        );

    \I__4208\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22789\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__22789\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__4206\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22783\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__22783\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__4204\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22777\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__22777\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__4202\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22771\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__22771\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__4200\ : CEMux
    port map (
            O => \N__22768\,
            I => \N__22765\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__22765\,
            I => \N__22761\
        );

    \I__4198\ : CEMux
    port map (
            O => \N__22764\,
            I => \N__22758\
        );

    \I__4197\ : Span4Mux_v
    port map (
            O => \N__22761\,
            I => \N__22753\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__22758\,
            I => \N__22753\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__22753\,
            I => \N__22750\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__22747\,
            I => \this_spr_ram.mem_WE_10\
        );

    \I__4192\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22739\
        );

    \I__4191\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22736\
        );

    \I__4190\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22730\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__22739\,
            I => \N__22726\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__22736\,
            I => \N__22723\
        );

    \I__4187\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22720\
        );

    \I__4186\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22717\
        );

    \I__4185\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22714\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22711\
        );

    \I__4183\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22708\
        );

    \I__4182\ : Sp12to4
    port map (
            O => \N__22726\,
            I => \N__22704\
        );

    \I__4181\ : Span4Mux_h
    port map (
            O => \N__22723\,
            I => \N__22701\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__22720\,
            I => \N__22698\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__22717\,
            I => \N__22695\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__22714\,
            I => \N__22692\
        );

    \I__4177\ : Span12Mux_h
    port map (
            O => \N__22711\,
            I => \N__22689\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__22708\,
            I => \N__22686\
        );

    \I__4175\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22683\
        );

    \I__4174\ : Span12Mux_v
    port map (
            O => \N__22704\,
            I => \N__22680\
        );

    \I__4173\ : Span4Mux_h
    port map (
            O => \N__22701\,
            I => \N__22677\
        );

    \I__4172\ : Span12Mux_h
    port map (
            O => \N__22698\,
            I => \N__22670\
        );

    \I__4171\ : Span12Mux_h
    port map (
            O => \N__22695\,
            I => \N__22670\
        );

    \I__4170\ : Span12Mux_h
    port map (
            O => \N__22692\,
            I => \N__22670\
        );

    \I__4169\ : Span12Mux_v
    port map (
            O => \N__22689\,
            I => \N__22663\
        );

    \I__4168\ : Span12Mux_h
    port map (
            O => \N__22686\,
            I => \N__22663\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22663\
        );

    \I__4166\ : Odrv12
    port map (
            O => \N__22680\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__22677\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__4164\ : Odrv12
    port map (
            O => \N__22670\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__4163\ : Odrv12
    port map (
            O => \N__22663\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__22654\,
            I => \N__22651\
        );

    \I__4161\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22648\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__22648\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__22645\,
            I => \N__22641\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__22644\,
            I => \N__22637\
        );

    \I__4157\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22634\
        );

    \I__4156\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22629\
        );

    \I__4155\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22629\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__22634\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__22629\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__4152\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22621\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__22621\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__22618\,
            I => \N__22614\
        );

    \I__4149\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22610\
        );

    \I__4148\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22605\
        );

    \I__4147\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22605\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__22610\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__22605\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__4144\ : IoInMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__22594\,
            I => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\
        );

    \I__4141\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22588\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__22588\,
            I => \N__22585\
        );

    \I__4139\ : Span12Mux_h
    port map (
            O => \N__22585\,
            I => \N__22582\
        );

    \I__4138\ : Odrv12
    port map (
            O => \N__22582\,
            I => \this_spr_ram.mem_out_bus4_3\
        );

    \I__4137\ : InMux
    port map (
            O => \N__22579\,
            I => \N__22576\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__22576\,
            I => \N__22573\
        );

    \I__4135\ : Span12Mux_h
    port map (
            O => \N__22573\,
            I => \N__22570\
        );

    \I__4134\ : Odrv12
    port map (
            O => \N__22570\,
            I => \this_spr_ram.mem_out_bus0_3\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__22567\,
            I => \N__22564\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22561\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__22561\,
            I => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\
        );

    \I__4130\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22555\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__22555\,
            I => \this_reset_cond.M_stage_qZ0Z_8\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22549\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__22549\,
            I => \N__22546\
        );

    \I__4126\ : Span12Mux_v
    port map (
            O => \N__22546\,
            I => \N__22543\
        );

    \I__4125\ : Odrv12
    port map (
            O => \N__22543\,
            I => \this_spr_ram.mem_out_bus7_3\
        );

    \I__4124\ : InMux
    port map (
            O => \N__22540\,
            I => \N__22537\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__4122\ : Span4Mux_h
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__22528\,
            I => \this_spr_ram.mem_out_bus3_3\
        );

    \I__4119\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__22522\,
            I => \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\
        );

    \I__4117\ : InMux
    port map (
            O => \N__22519\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1\
        );

    \I__4116\ : InMux
    port map (
            O => \N__22516\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1\
        );

    \I__4115\ : InMux
    port map (
            O => \N__22513\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1\
        );

    \I__4114\ : InMux
    port map (
            O => \N__22510\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1\
        );

    \I__4113\ : InMux
    port map (
            O => \N__22507\,
            I => \this_ppu.un1_M_count_q_1_cry_6_s1\
        );

    \I__4112\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__22501\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_7\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__22498\,
            I => \N__22495\
        );

    \I__4109\ : InMux
    port map (
            O => \N__22495\,
            I => \N__22492\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__22492\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__22489\,
            I => \N__22485\
        );

    \I__4106\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22481\
        );

    \I__4105\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22478\
        );

    \I__4104\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22475\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__22481\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__22478\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__22475\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__22468\,
            I => \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_4_cascade_\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__22465\,
            I => \N__22462\
        );

    \I__4098\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22459\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__22459\,
            I => \N__22456\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__22456\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\
        );

    \I__4095\ : InMux
    port map (
            O => \N__22453\,
            I => \N__22449\
        );

    \I__4094\ : CascadeMux
    port map (
            O => \N__22452\,
            I => \N__22446\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__22449\,
            I => \N__22442\
        );

    \I__4092\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22439\
        );

    \I__4091\ : InMux
    port map (
            O => \N__22445\,
            I => \N__22436\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__22442\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__22439\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__22436\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__22429\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_11_cascade_\
        );

    \I__4086\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__22423\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_11\
        );

    \I__4084\ : InMux
    port map (
            O => \N__22420\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1\
        );

    \I__4083\ : InMux
    port map (
            O => \N__22417\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1\
        );

    \I__4082\ : SRMux
    port map (
            O => \N__22414\,
            I => \N__22410\
        );

    \I__4081\ : SRMux
    port map (
            O => \N__22413\,
            I => \N__22406\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22402\
        );

    \I__4079\ : SRMux
    port map (
            O => \N__22409\,
            I => \N__22399\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__22406\,
            I => \N__22396\
        );

    \I__4077\ : SRMux
    port map (
            O => \N__22405\,
            I => \N__22393\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__22402\,
            I => \N__22388\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__22399\,
            I => \N__22388\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__22396\,
            I => \N__22385\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22382\
        );

    \I__4072\ : Span4Mux_h
    port map (
            O => \N__22388\,
            I => \N__22379\
        );

    \I__4071\ : Odrv4
    port map (
            O => \N__22385\,
            I => \this_ppu.M_last_q_RNIGL6V4\
        );

    \I__4070\ : Odrv12
    port map (
            O => \N__22382\,
            I => \this_ppu.M_last_q_RNIGL6V4\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__22379\,
            I => \this_ppu.M_last_q_RNIGL6V4\
        );

    \I__4068\ : CEMux
    port map (
            O => \N__22372\,
            I => \N__22369\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__22369\,
            I => \N__22365\
        );

    \I__4066\ : CEMux
    port map (
            O => \N__22368\,
            I => \N__22362\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__22365\,
            I => \N__22357\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__22362\,
            I => \N__22357\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__22354\,
            I => \N__22351\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__22351\,
            I => \this_spr_ram.mem_WE_8\
        );

    \I__4060\ : InMux
    port map (
            O => \N__22348\,
            I => \N__22345\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__22345\,
            I => \N__22342\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__4057\ : Span4Mux_v
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__4056\ : Span4Mux_v
    port map (
            O => \N__22336\,
            I => \N__22333\
        );

    \I__4055\ : Span4Mux_h
    port map (
            O => \N__22333\,
            I => \N__22330\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__22330\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__4052\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22320\
        );

    \I__4051\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22315\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__22320\,
            I => \N__22312\
        );

    \I__4049\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22307\
        );

    \I__4048\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22307\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__22315\,
            I => \N__22304\
        );

    \I__4046\ : Span4Mux_h
    port map (
            O => \N__22312\,
            I => \N__22299\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22299\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__22304\,
            I => \N__22296\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__22299\,
            I => \this_spr_ram.mem_radregZ0Z_12\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__22296\,
            I => \this_spr_ram.mem_radregZ0Z_12\
        );

    \I__4041\ : InMux
    port map (
            O => \N__22291\,
            I => \N__22288\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__22288\,
            I => \N__22285\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__22285\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__4038\ : InMux
    port map (
            O => \N__22282\,
            I => \N__22279\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22276\
        );

    \I__4036\ : Span4Mux_v
    port map (
            O => \N__22276\,
            I => \N__22273\
        );

    \I__4035\ : Sp12to4
    port map (
            O => \N__22273\,
            I => \N__22270\
        );

    \I__4034\ : Span12Mux_h
    port map (
            O => \N__22270\,
            I => \N__22267\
        );

    \I__4033\ : Odrv12
    port map (
            O => \N__22267\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__4032\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22258\
        );

    \I__4031\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22255\
        );

    \I__4030\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22251\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__22261\,
            I => \N__22248\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__22258\,
            I => \N__22244\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__22255\,
            I => \N__22241\
        );

    \I__4026\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22238\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__22251\,
            I => \N__22235\
        );

    \I__4024\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22230\
        );

    \I__4023\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22227\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__22244\,
            I => \N__22224\
        );

    \I__4021\ : Span4Mux_h
    port map (
            O => \N__22241\,
            I => \N__22221\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__22238\,
            I => \N__22216\
        );

    \I__4019\ : Span4Mux_h
    port map (
            O => \N__22235\,
            I => \N__22216\
        );

    \I__4018\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22211\
        );

    \I__4017\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22211\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__22230\,
            I => \N__22208\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22205\
        );

    \I__4014\ : Span4Mux_v
    port map (
            O => \N__22224\,
            I => \N__22202\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__22221\,
            I => \N__22199\
        );

    \I__4012\ : Span4Mux_v
    port map (
            O => \N__22216\,
            I => \N__22196\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__22211\,
            I => \N__22193\
        );

    \I__4010\ : Span4Mux_v
    port map (
            O => \N__22208\,
            I => \N__22188\
        );

    \I__4009\ : Span4Mux_h
    port map (
            O => \N__22205\,
            I => \N__22188\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__22202\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__22199\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__22196\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__4005\ : Odrv12
    port map (
            O => \N__22193\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__22188\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__4003\ : CEMux
    port map (
            O => \N__22177\,
            I => \N__22174\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__22174\,
            I => \N__22170\
        );

    \I__4001\ : InMux
    port map (
            O => \N__22173\,
            I => \N__22167\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__22170\,
            I => \N__22154\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__22167\,
            I => \N__22154\
        );

    \I__3998\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22151\
        );

    \I__3997\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22146\
        );

    \I__3996\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22146\
        );

    \I__3995\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22143\
        );

    \I__3994\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22140\
        );

    \I__3993\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22137\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__22160\,
            I => \N__22132\
        );

    \I__3991\ : CEMux
    port map (
            O => \N__22159\,
            I => \N__22129\
        );

    \I__3990\ : Span4Mux_h
    port map (
            O => \N__22154\,
            I => \N__22124\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22124\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__22146\,
            I => \N__22119\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__22143\,
            I => \N__22119\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__22140\,
            I => \N__22114\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__22137\,
            I => \N__22114\
        );

    \I__3984\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22111\
        );

    \I__3983\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22108\
        );

    \I__3982\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22105\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__22129\,
            I => \N__22102\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__22124\,
            I => \N__22099\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__22119\,
            I => \N__22094\
        );

    \I__3978\ : Span4Mux_h
    port map (
            O => \N__22114\,
            I => \N__22094\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__22111\,
            I => \N__22087\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__22108\,
            I => \N__22087\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__22105\,
            I => \N__22087\
        );

    \I__3974\ : Span12Mux_v
    port map (
            O => \N__22102\,
            I => \N__22084\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__22099\,
            I => \N__22081\
        );

    \I__3972\ : Span4Mux_h
    port map (
            O => \N__22094\,
            I => \N__22078\
        );

    \I__3971\ : Span12Mux_h
    port map (
            O => \N__22087\,
            I => \N__22075\
        );

    \I__3970\ : Odrv12
    port map (
            O => \N__22084\,
            I => \M_this_state_d_0_sqmuxa\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__22081\,
            I => \M_this_state_d_0_sqmuxa\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__22078\,
            I => \M_this_state_d_0_sqmuxa\
        );

    \I__3967\ : Odrv12
    port map (
            O => \N__22075\,
            I => \M_this_state_d_0_sqmuxa\
        );

    \I__3966\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22063\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__3964\ : Span4Mux_v
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__3963\ : Sp12to4
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__3962\ : Odrv12
    port map (
            O => \N__22054\,
            I => \this_spr_ram.mem_out_bus6_1\
        );

    \I__3961\ : InMux
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__22048\,
            I => \N__22045\
        );

    \I__3959\ : Span4Mux_h
    port map (
            O => \N__22045\,
            I => \N__22042\
        );

    \I__3958\ : Span4Mux_v
    port map (
            O => \N__22042\,
            I => \N__22039\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__22039\,
            I => \N__22036\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__22036\,
            I => \this_spr_ram.mem_out_bus2_1\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__22033\,
            I => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0_cascade_\
        );

    \I__3954\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22027\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__22027\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1\
        );

    \I__3952\ : CEMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__22017\
        );

    \I__3950\ : CEMux
    port map (
            O => \N__22020\,
            I => \N__22014\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__22017\,
            I => \N__22009\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__22014\,
            I => \N__22009\
        );

    \I__3947\ : Span4Mux_h
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__22003\,
            I => \this_spr_ram.mem_WE_6\
        );

    \I__3944\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__21997\,
            I => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__21994\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\
        );

    \I__3941\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21987\
        );

    \I__3940\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21984\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21981\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__21984\,
            I => \N__21978\
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__21981\,
            I => \M_this_spr_ram_read_data_3\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__21978\,
            I => \M_this_spr_ram_read_data_3\
        );

    \I__3935\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21970\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__21970\,
            I => \N__21967\
        );

    \I__3933\ : Span4Mux_h
    port map (
            O => \N__21967\,
            I => \N__21964\
        );

    \I__3932\ : Span4Mux_h
    port map (
            O => \N__21964\,
            I => \N__21961\
        );

    \I__3931\ : Odrv4
    port map (
            O => \N__21961\,
            I => \this_spr_ram.mem_out_bus4_1\
        );

    \I__3930\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21955\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__21955\,
            I => \N__21952\
        );

    \I__3928\ : Sp12to4
    port map (
            O => \N__21952\,
            I => \N__21949\
        );

    \I__3927\ : Span12Mux_v
    port map (
            O => \N__21949\,
            I => \N__21946\
        );

    \I__3926\ : Odrv12
    port map (
            O => \N__21946\,
            I => \this_spr_ram.mem_out_bus0_1\
        );

    \I__3925\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21940\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__21940\,
            I => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21934\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__21934\,
            I => \this_ppu.un1_M_haddress_q_c6\
        );

    \I__3921\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21923\
        );

    \I__3920\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21923\
        );

    \I__3919\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21920\
        );

    \I__3918\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21917\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__21923\,
            I => \this_ppu.N_754_0\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__21920\,
            I => \this_ppu.N_754_0\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__21917\,
            I => \this_ppu.N_754_0\
        );

    \I__3914\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21906\
        );

    \I__3913\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21903\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__21906\,
            I => \this_ppu.un1_M_haddress_q_c2\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__21903\,
            I => \this_ppu.un1_M_haddress_q_c2\
        );

    \I__3910\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__21895\,
            I => \this_ppu.M_state_qZ0Z_8\
        );

    \I__3908\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__3906\ : Span4Mux_v
    port map (
            O => \N__21886\,
            I => \N__21883\
        );

    \I__3905\ : Sp12to4
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__21880\,
            I => \this_spr_ram.mem_out_bus6_3\
        );

    \I__3903\ : InMux
    port map (
            O => \N__21877\,
            I => \N__21874\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__21874\,
            I => \N__21871\
        );

    \I__3901\ : Span4Mux_v
    port map (
            O => \N__21871\,
            I => \N__21868\
        );

    \I__3900\ : Span4Mux_h
    port map (
            O => \N__21868\,
            I => \N__21865\
        );

    \I__3899\ : Span4Mux_h
    port map (
            O => \N__21865\,
            I => \N__21862\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__21862\,
            I => \this_spr_ram.mem_out_bus2_3\
        );

    \I__3897\ : InMux
    port map (
            O => \N__21859\,
            I => \N__21856\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__21856\,
            I => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\
        );

    \I__3895\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21850\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21846\
        );

    \I__3893\ : InMux
    port map (
            O => \N__21849\,
            I => \N__21843\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__21846\,
            I => \M_this_spr_ram_read_data_1\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__21843\,
            I => \M_this_spr_ram_read_data_1\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__21838\,
            I => \this_ppu.un1_M_haddress_q_c3_cascade_\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__21835\,
            I => \this_ppu.un1_M_haddress_q_c6_cascade_\
        );

    \I__3888\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21829\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__21829\,
            I => \this_ppu.un1_M_haddress_q_c3\
        );

    \I__3886\ : InMux
    port map (
            O => \N__21826\,
            I => \N__21823\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__3883\ : Sp12to4
    port map (
            O => \N__21817\,
            I => \N__21814\
        );

    \I__3882\ : Span12Mux_h
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__21811\,
            I => \this_spr_ram.mem_out_bus7_1\
        );

    \I__3880\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21805\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__21805\,
            I => \N__21802\
        );

    \I__3878\ : Span4Mux_h
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__21796\,
            I => \this_spr_ram.mem_out_bus3_1\
        );

    \I__3875\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21790\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__21784\,
            I => \N__21781\
        );

    \I__3871\ : Span4Mux_h
    port map (
            O => \N__21781\,
            I => \N__21778\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__21778\,
            I => \this_spr_ram.mem_out_bus6_0\
        );

    \I__3869\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21772\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__21772\,
            I => \N__21769\
        );

    \I__3867\ : Span4Mux_h
    port map (
            O => \N__21769\,
            I => \N__21766\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__21766\,
            I => \N__21763\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__21763\,
            I => \N__21760\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__21760\,
            I => \this_spr_ram.mem_out_bus2_0\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__21757\,
            I => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\
        );

    \I__3862\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21751\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__21751\,
            I => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\
        );

    \I__3860\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21745\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__21745\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__3858\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21739\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__21739\,
            I => \N__21736\
        );

    \I__3856\ : Span12Mux_h
    port map (
            O => \N__21736\,
            I => \N__21733\
        );

    \I__3855\ : Odrv12
    port map (
            O => \N__21733\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__3854\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21727\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21724\
        );

    \I__3852\ : Span12Mux_v
    port map (
            O => \N__21724\,
            I => \N__21721\
        );

    \I__3851\ : Span12Mux_h
    port map (
            O => \N__21721\,
            I => \N__21718\
        );

    \I__3850\ : Odrv12
    port map (
            O => \N__21718\,
            I => \this_ppu.oam_cache.mem_2\
        );

    \I__3849\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__3847\ : Odrv12
    port map (
            O => \N__21709\,
            I => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_2\
        );

    \I__3846\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21703\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__21703\,
            I => \N__21700\
        );

    \I__3844\ : Odrv12
    port map (
            O => \N__21700\,
            I => \M_this_map_ram_write_data_6\
        );

    \I__3843\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21694\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__21694\,
            I => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0\
        );

    \I__3841\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21688\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__21688\,
            I => \N__21685\
        );

    \I__3839\ : Span4Mux_h
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__21679\,
            I => \N__21676\
        );

    \I__3836\ : Span4Mux_v
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__21673\,
            I => \this_spr_ram.mem_out_bus7_2\
        );

    \I__3834\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21667\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21664\
        );

    \I__3832\ : Span4Mux_h
    port map (
            O => \N__21664\,
            I => \N__21661\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__21658\,
            I => \this_spr_ram.mem_out_bus3_2\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__21655\,
            I => \this_spr_ram.mem_mem_3_1_RNISI5GZ0_cascade_\
        );

    \I__3828\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__21649\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2\
        );

    \I__3826\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__21640\,
            I => \M_this_spr_ram_read_data_2\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__21637\,
            I => \M_this_spr_ram_read_data_2_cascade_\
        );

    \I__3822\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21631\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__21631\,
            I => \N__21628\
        );

    \I__3820\ : Span4Mux_h
    port map (
            O => \N__21628\,
            I => \N__21625\
        );

    \I__3819\ : Span4Mux_h
    port map (
            O => \N__21625\,
            I => \N__21622\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__21622\,
            I => \N__21619\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__21619\,
            I => \this_spr_ram.mem_out_bus6_2\
        );

    \I__3816\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__21613\,
            I => \N__21610\
        );

    \I__3814\ : Span4Mux_h
    port map (
            O => \N__21610\,
            I => \N__21607\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__3812\ : Span4Mux_h
    port map (
            O => \N__21604\,
            I => \N__21601\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__21601\,
            I => \this_spr_ram.mem_out_bus2_2\
        );

    \I__3810\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__21595\,
            I => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0\
        );

    \I__3808\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__21589\,
            I => \N__21586\
        );

    \I__3806\ : Span4Mux_h
    port map (
            O => \N__21586\,
            I => \N__21583\
        );

    \I__3805\ : Sp12to4
    port map (
            O => \N__21583\,
            I => \N__21580\
        );

    \I__3804\ : Span12Mux_v
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__3803\ : Odrv12
    port map (
            O => \N__21577\,
            I => \this_spr_ram.mem_out_bus7_0\
        );

    \I__3802\ : InMux
    port map (
            O => \N__21574\,
            I => \N__21571\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__21571\,
            I => \N__21568\
        );

    \I__3800\ : Span4Mux_h
    port map (
            O => \N__21568\,
            I => \N__21565\
        );

    \I__3799\ : Span4Mux_h
    port map (
            O => \N__21565\,
            I => \N__21562\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__21562\,
            I => \this_spr_ram.mem_out_bus3_0\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__21559\,
            I => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0_cascade_\
        );

    \I__3796\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21552\
        );

    \I__3795\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21549\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__21552\,
            I => \M_this_spr_ram_read_data_0\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__21549\,
            I => \M_this_spr_ram_read_data_0\
        );

    \I__3792\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21541\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__21538\,
            I => \N__21535\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__21535\,
            I => \N__21532\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__21532\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__3787\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21524\
        );

    \I__3786\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21519\
        );

    \I__3785\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21519\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__21524\,
            I => \this_ppu.N_806\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__21519\,
            I => \this_ppu.N_806\
        );

    \I__3782\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21511\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__21511\,
            I => \N__21508\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__3779\ : Span4Mux_h
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__21502\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__3777\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21496\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__3775\ : Span4Mux_h
    port map (
            O => \N__21493\,
            I => \N__21490\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__21490\,
            I => \N__21487\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__21487\,
            I => \this_spr_ram.mem_out_bus4_0\
        );

    \I__3772\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21481\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21478\
        );

    \I__3770\ : Span12Mux_v
    port map (
            O => \N__21478\,
            I => \N__21475\
        );

    \I__3769\ : Span12Mux_h
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__3768\ : Odrv12
    port map (
            O => \N__21472\,
            I => \this_spr_ram.mem_out_bus0_0\
        );

    \I__3767\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21466\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__21466\,
            I => \N__21463\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__21463\,
            I => \N__21460\
        );

    \I__3764\ : Span4Mux_h
    port map (
            O => \N__21460\,
            I => \N__21457\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__21457\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__3762\ : CascadeMux
    port map (
            O => \N__21454\,
            I => \N__21449\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__21453\,
            I => \N__21444\
        );

    \I__3760\ : CascadeMux
    port map (
            O => \N__21452\,
            I => \N__21441\
        );

    \I__3759\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21436\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__21448\,
            I => \N__21433\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__21447\,
            I => \N__21430\
        );

    \I__3756\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21420\
        );

    \I__3755\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21417\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__21440\,
            I => \N__21414\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__21439\,
            I => \N__21411\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__21436\,
            I => \N__21406\
        );

    \I__3751\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21403\
        );

    \I__3750\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21400\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__21429\,
            I => \N__21397\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__21428\,
            I => \N__21394\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__21427\,
            I => \N__21391\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__21426\,
            I => \N__21388\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__21425\,
            I => \N__21385\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__21424\,
            I => \N__21382\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__21423\,
            I => \N__21379\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__21420\,
            I => \N__21376\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21373\
        );

    \I__3740\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21370\
        );

    \I__3739\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21367\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__21410\,
            I => \N__21364\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__21409\,
            I => \N__21361\
        );

    \I__3736\ : Sp12to4
    port map (
            O => \N__21406\,
            I => \N__21356\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__21403\,
            I => \N__21356\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__21400\,
            I => \N__21353\
        );

    \I__3733\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21350\
        );

    \I__3732\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21347\
        );

    \I__3731\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21344\
        );

    \I__3730\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21341\
        );

    \I__3729\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21338\
        );

    \I__3728\ : InMux
    port map (
            O => \N__21382\,
            I => \N__21335\
        );

    \I__3727\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21332\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__21376\,
            I => \N__21325\
        );

    \I__3725\ : Span4Mux_h
    port map (
            O => \N__21373\,
            I => \N__21325\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__21370\,
            I => \N__21325\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__21367\,
            I => \N__21322\
        );

    \I__3722\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21319\
        );

    \I__3721\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21316\
        );

    \I__3720\ : Span12Mux_s4_v
    port map (
            O => \N__21356\,
            I => \N__21311\
        );

    \I__3719\ : Span12Mux_s7_h
    port map (
            O => \N__21353\,
            I => \N__21311\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__21350\,
            I => \N__21300\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__21347\,
            I => \N__21300\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21300\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__21341\,
            I => \N__21300\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__21338\,
            I => \N__21300\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21297\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21294\
        );

    \I__3711\ : Span4Mux_v
    port map (
            O => \N__21325\,
            I => \N__21287\
        );

    \I__3710\ : Span4Mux_h
    port map (
            O => \N__21322\,
            I => \N__21287\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__21319\,
            I => \N__21287\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21284\
        );

    \I__3707\ : Span12Mux_h
    port map (
            O => \N__21311\,
            I => \N__21281\
        );

    \I__3706\ : Span12Mux_v
    port map (
            O => \N__21300\,
            I => \N__21274\
        );

    \I__3705\ : Span12Mux_v
    port map (
            O => \N__21297\,
            I => \N__21274\
        );

    \I__3704\ : Span12Mux_s7_h
    port map (
            O => \N__21294\,
            I => \N__21274\
        );

    \I__3703\ : Span4Mux_v
    port map (
            O => \N__21287\,
            I => \N__21269\
        );

    \I__3702\ : Span4Mux_h
    port map (
            O => \N__21284\,
            I => \N__21269\
        );

    \I__3701\ : Span12Mux_v
    port map (
            O => \N__21281\,
            I => \N__21264\
        );

    \I__3700\ : Span12Mux_h
    port map (
            O => \N__21274\,
            I => \N__21264\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__21269\,
            I => \N__21261\
        );

    \I__3698\ : Odrv12
    port map (
            O => \N__21264\,
            I => \M_this_ppu_spr_addr_8\
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__21261\,
            I => \M_this_ppu_spr_addr_8\
        );

    \I__3696\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21253\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__21253\,
            I => \N__21250\
        );

    \I__3694\ : Span12Mux_h
    port map (
            O => \N__21250\,
            I => \N__21247\
        );

    \I__3693\ : Odrv12
    port map (
            O => \N__21247\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__21244\,
            I => \N__21240\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__21243\,
            I => \N__21237\
        );

    \I__3690\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21232\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21229\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__21236\,
            I => \N__21226\
        );

    \I__3687\ : CascadeMux
    port map (
            O => \N__21235\,
            I => \N__21223\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21215\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21215\
        );

    \I__3684\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21212\
        );

    \I__3683\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21209\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__21222\,
            I => \N__21206\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__21221\,
            I => \N__21203\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__21220\,
            I => \N__21197\
        );

    \I__3679\ : Span4Mux_s3_v
    port map (
            O => \N__21215\,
            I => \N__21189\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__21212\,
            I => \N__21189\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__21209\,
            I => \N__21189\
        );

    \I__3676\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21186\
        );

    \I__3675\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21183\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__21202\,
            I => \N__21180\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__21201\,
            I => \N__21177\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__21200\,
            I => \N__21172\
        );

    \I__3671\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21168\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__21196\,
            I => \N__21165\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21159\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21159\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__21183\,
            I => \N__21156\
        );

    \I__3666\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21153\
        );

    \I__3665\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21150\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__21176\,
            I => \N__21147\
        );

    \I__3663\ : CascadeMux
    port map (
            O => \N__21175\,
            I => \N__21144\
        );

    \I__3662\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21141\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__21171\,
            I => \N__21138\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__21168\,
            I => \N__21135\
        );

    \I__3659\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21132\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__21164\,
            I => \N__21129\
        );

    \I__3657\ : Span4Mux_v
    port map (
            O => \N__21159\,
            I => \N__21119\
        );

    \I__3656\ : Span4Mux_v
    port map (
            O => \N__21156\,
            I => \N__21119\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__21153\,
            I => \N__21119\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__21150\,
            I => \N__21119\
        );

    \I__3653\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21116\
        );

    \I__3652\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21113\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__21141\,
            I => \N__21110\
        );

    \I__3650\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21107\
        );

    \I__3649\ : Span4Mux_h
    port map (
            O => \N__21135\,
            I => \N__21102\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__21132\,
            I => \N__21102\
        );

    \I__3647\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21099\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__21128\,
            I => \N__21096\
        );

    \I__3645\ : Span4Mux_v
    port map (
            O => \N__21119\,
            I => \N__21089\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__21116\,
            I => \N__21089\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__21113\,
            I => \N__21089\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__21110\,
            I => \N__21084\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__21107\,
            I => \N__21084\
        );

    \I__3640\ : Span4Mux_v
    port map (
            O => \N__21102\,
            I => \N__21079\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21079\
        );

    \I__3638\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21076\
        );

    \I__3637\ : Span4Mux_v
    port map (
            O => \N__21089\,
            I => \N__21073\
        );

    \I__3636\ : Span4Mux_v
    port map (
            O => \N__21084\,
            I => \N__21066\
        );

    \I__3635\ : Span4Mux_v
    port map (
            O => \N__21079\,
            I => \N__21066\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__21076\,
            I => \N__21066\
        );

    \I__3633\ : Span4Mux_h
    port map (
            O => \N__21073\,
            I => \N__21063\
        );

    \I__3632\ : Span4Mux_v
    port map (
            O => \N__21066\,
            I => \N__21060\
        );

    \I__3631\ : Span4Mux_h
    port map (
            O => \N__21063\,
            I => \N__21057\
        );

    \I__3630\ : Span4Mux_h
    port map (
            O => \N__21060\,
            I => \N__21054\
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__21057\,
            I => \M_this_ppu_spr_addr_7\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__21054\,
            I => \M_this_ppu_spr_addr_7\
        );

    \I__3627\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21046\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__21046\,
            I => \N__21043\
        );

    \I__3625\ : Span4Mux_h
    port map (
            O => \N__21043\,
            I => \N__21040\
        );

    \I__3624\ : Span4Mux_h
    port map (
            O => \N__21040\,
            I => \N__21037\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__21037\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__21034\,
            I => \N__21031\
        );

    \I__3621\ : InMux
    port map (
            O => \N__21031\,
            I => \N__21026\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__21030\,
            I => \N__21023\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__21029\,
            I => \N__21020\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21005\
        );

    \I__3617\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21002\
        );

    \I__3616\ : InMux
    port map (
            O => \N__21020\,
            I => \N__20999\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__21019\,
            I => \N__20996\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__21018\,
            I => \N__20993\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__21017\,
            I => \N__20989\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__21016\,
            I => \N__20986\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__21015\,
            I => \N__20983\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__21014\,
            I => \N__20980\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__21013\,
            I => \N__20977\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__21012\,
            I => \N__20974\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__21011\,
            I => \N__20971\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__21010\,
            I => \N__20968\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__21009\,
            I => \N__20965\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__21008\,
            I => \N__20962\
        );

    \I__3603\ : Span4Mux_v
    port map (
            O => \N__21005\,
            I => \N__20955\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__21002\,
            I => \N__20955\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20955\
        );

    \I__3600\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20952\
        );

    \I__3599\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20949\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__20992\,
            I => \N__20946\
        );

    \I__3597\ : InMux
    port map (
            O => \N__20989\,
            I => \N__20943\
        );

    \I__3596\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20940\
        );

    \I__3595\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20937\
        );

    \I__3594\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20934\
        );

    \I__3593\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20931\
        );

    \I__3592\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20928\
        );

    \I__3591\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20925\
        );

    \I__3590\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20922\
        );

    \I__3589\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20919\
        );

    \I__3588\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20916\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__20955\,
            I => \N__20909\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20909\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20909\
        );

    \I__3584\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20906\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20893\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__20940\,
            I => \N__20893\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__20937\,
            I => \N__20893\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__20934\,
            I => \N__20893\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__20931\,
            I => \N__20893\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__20928\,
            I => \N__20893\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20884\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__20922\,
            I => \N__20884\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__20919\,
            I => \N__20884\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20884\
        );

    \I__3573\ : Span4Mux_v
    port map (
            O => \N__20909\,
            I => \N__20879\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20879\
        );

    \I__3571\ : Span12Mux_s11_v
    port map (
            O => \N__20893\,
            I => \N__20876\
        );

    \I__3570\ : Span12Mux_v
    port map (
            O => \N__20884\,
            I => \N__20873\
        );

    \I__3569\ : Span4Mux_v
    port map (
            O => \N__20879\,
            I => \N__20870\
        );

    \I__3568\ : Span12Mux_h
    port map (
            O => \N__20876\,
            I => \N__20865\
        );

    \I__3567\ : Span12Mux_h
    port map (
            O => \N__20873\,
            I => \N__20865\
        );

    \I__3566\ : Span4Mux_h
    port map (
            O => \N__20870\,
            I => \N__20862\
        );

    \I__3565\ : Odrv12
    port map (
            O => \N__20865\,
            I => \M_this_ppu_spr_addr_9\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__20862\,
            I => \M_this_ppu_spr_addr_9\
        );

    \I__3563\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20854\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__20854\,
            I => \N__20851\
        );

    \I__3561\ : Span4Mux_h
    port map (
            O => \N__20851\,
            I => \N__20848\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__20848\,
            I => \N__20845\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__20845\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__20842\,
            I => \N__20828\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__20841\,
            I => \N__20825\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__20840\,
            I => \N__20822\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__20839\,
            I => \N__20819\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__20838\,
            I => \N__20816\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__20837\,
            I => \N__20812\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__20836\,
            I => \N__20809\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__20835\,
            I => \N__20806\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__20834\,
            I => \N__20802\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__20833\,
            I => \N__20799\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__20832\,
            I => \N__20796\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__20831\,
            I => \N__20793\
        );

    \I__3546\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20790\
        );

    \I__3545\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20787\
        );

    \I__3544\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20784\
        );

    \I__3543\ : InMux
    port map (
            O => \N__20819\,
            I => \N__20781\
        );

    \I__3542\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20776\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__20815\,
            I => \N__20773\
        );

    \I__3540\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20770\
        );

    \I__3539\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20767\
        );

    \I__3538\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20764\
        );

    \I__3537\ : CascadeMux
    port map (
            O => \N__20805\,
            I => \N__20761\
        );

    \I__3536\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20758\
        );

    \I__3535\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20755\
        );

    \I__3534\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20752\
        );

    \I__3533\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20749\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__20790\,
            I => \N__20744\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__20787\,
            I => \N__20744\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__20784\,
            I => \N__20739\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__20781\,
            I => \N__20739\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__20780\,
            I => \N__20736\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__20779\,
            I => \N__20733\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__20776\,
            I => \N__20730\
        );

    \I__3525\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20727\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__20770\,
            I => \N__20722\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__20767\,
            I => \N__20722\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20719\
        );

    \I__3521\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20716\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__20758\,
            I => \N__20711\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__20755\,
            I => \N__20711\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__20752\,
            I => \N__20708\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20705\
        );

    \I__3516\ : Span4Mux_v
    port map (
            O => \N__20744\,
            I => \N__20700\
        );

    \I__3515\ : Span4Mux_v
    port map (
            O => \N__20739\,
            I => \N__20700\
        );

    \I__3514\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20697\
        );

    \I__3513\ : InMux
    port map (
            O => \N__20733\,
            I => \N__20694\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__20730\,
            I => \N__20689\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__20727\,
            I => \N__20689\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__20722\,
            I => \N__20684\
        );

    \I__3509\ : Span4Mux_v
    port map (
            O => \N__20719\,
            I => \N__20684\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20679\
        );

    \I__3507\ : Span4Mux_v
    port map (
            O => \N__20711\,
            I => \N__20679\
        );

    \I__3506\ : Span4Mux_s1_v
    port map (
            O => \N__20708\,
            I => \N__20674\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__20705\,
            I => \N__20674\
        );

    \I__3504\ : Sp12to4
    port map (
            O => \N__20700\,
            I => \N__20671\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__20697\,
            I => \N__20664\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__20694\,
            I => \N__20664\
        );

    \I__3501\ : Sp12to4
    port map (
            O => \N__20689\,
            I => \N__20664\
        );

    \I__3500\ : Span4Mux_h
    port map (
            O => \N__20684\,
            I => \N__20659\
        );

    \I__3499\ : Span4Mux_v
    port map (
            O => \N__20679\,
            I => \N__20659\
        );

    \I__3498\ : Sp12to4
    port map (
            O => \N__20674\,
            I => \N__20656\
        );

    \I__3497\ : Span12Mux_h
    port map (
            O => \N__20671\,
            I => \N__20653\
        );

    \I__3496\ : Span12Mux_v
    port map (
            O => \N__20664\,
            I => \N__20650\
        );

    \I__3495\ : Span4Mux_h
    port map (
            O => \N__20659\,
            I => \N__20647\
        );

    \I__3494\ : Span12Mux_h
    port map (
            O => \N__20656\,
            I => \N__20644\
        );

    \I__3493\ : Span12Mux_v
    port map (
            O => \N__20653\,
            I => \N__20641\
        );

    \I__3492\ : Span12Mux_h
    port map (
            O => \N__20650\,
            I => \N__20634\
        );

    \I__3491\ : Sp12to4
    port map (
            O => \N__20647\,
            I => \N__20634\
        );

    \I__3490\ : Span12Mux_v
    port map (
            O => \N__20644\,
            I => \N__20634\
        );

    \I__3489\ : Odrv12
    port map (
            O => \N__20641\,
            I => \M_this_ppu_spr_addr_10\
        );

    \I__3488\ : Odrv12
    port map (
            O => \N__20634\,
            I => \M_this_ppu_spr_addr_10\
        );

    \I__3487\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20626\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__20626\,
            I => \N__20623\
        );

    \I__3485\ : Span12Mux_v
    port map (
            O => \N__20623\,
            I => \N__20620\
        );

    \I__3484\ : Span12Mux_h
    port map (
            O => \N__20620\,
            I => \N__20617\
        );

    \I__3483\ : Odrv12
    port map (
            O => \N__20617\,
            I => \this_ppu.oam_cache.mem_3\
        );

    \I__3482\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20611\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__20611\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_3\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__20608\,
            I => \N__20603\
        );

    \I__3479\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20599\
        );

    \I__3478\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20596\
        );

    \I__3477\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20593\
        );

    \I__3476\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20590\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__20599\,
            I => \this_vga_signals_M_lcounter_q_0\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__20596\,
            I => \this_vga_signals_M_lcounter_q_0\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__20593\,
            I => \this_vga_signals_M_lcounter_q_0\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__20590\,
            I => \this_vga_signals_M_lcounter_q_0\
        );

    \I__3471\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20577\
        );

    \I__3470\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20574\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20571\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20568\
        );

    \I__3467\ : Span4Mux_v
    port map (
            O => \N__20571\,
            I => \N__20565\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__20568\,
            I => \N__20562\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__20565\,
            I => \N__20557\
        );

    \I__3464\ : Span4Mux_v
    port map (
            O => \N__20562\,
            I => \N__20557\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__20557\,
            I => \this_ppu.N_759_0\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__20554\,
            I => \N__20548\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__20553\,
            I => \N__20545\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__20552\,
            I => \N__20542\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__20551\,
            I => \N__20539\
        );

    \I__3458\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20536\
        );

    \I__3457\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20533\
        );

    \I__3456\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20530\
        );

    \I__3455\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20527\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__20536\,
            I => \this_vga_signals_M_lcounter_q_1\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__20533\,
            I => \this_vga_signals_M_lcounter_q_1\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__20530\,
            I => \this_vga_signals_M_lcounter_q_1\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__20527\,
            I => \this_vga_signals_M_lcounter_q_1\
        );

    \I__3450\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20515\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20507\
        );

    \I__3448\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20504\
        );

    \I__3447\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20501\
        );

    \I__3446\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20498\
        );

    \I__3445\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20495\
        );

    \I__3444\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20492\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__20507\,
            I => \N__20485\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20485\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__20501\,
            I => \N__20485\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__20498\,
            I => \N__20480\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__20495\,
            I => \N__20475\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20470\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__20485\,
            I => \N__20467\
        );

    \I__3436\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20464\
        );

    \I__3435\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20461\
        );

    \I__3434\ : Span4Mux_h
    port map (
            O => \N__20480\,
            I => \N__20458\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__20479\,
            I => \N__20455\
        );

    \I__3432\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20452\
        );

    \I__3431\ : Span4Mux_h
    port map (
            O => \N__20475\,
            I => \N__20449\
        );

    \I__3430\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20444\
        );

    \I__3429\ : InMux
    port map (
            O => \N__20473\,
            I => \N__20444\
        );

    \I__3428\ : Span4Mux_v
    port map (
            O => \N__20470\,
            I => \N__20440\
        );

    \I__3427\ : Span4Mux_h
    port map (
            O => \N__20467\,
            I => \N__20437\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__20464\,
            I => \N__20430\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__20461\,
            I => \N__20430\
        );

    \I__3424\ : Span4Mux_h
    port map (
            O => \N__20458\,
            I => \N__20430\
        );

    \I__3423\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20427\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20420\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__20449\,
            I => \N__20420\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__20444\,
            I => \N__20420\
        );

    \I__3419\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20417\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__20440\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__20437\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__20430\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__20427\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__20420\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__20417\,
            I => \this_vga_signals_M_vcounter_q_9\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__20404\,
            I => \this_ppu.N_5_4_cascade_\
        );

    \I__3411\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20398\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__3408\ : Sp12to4
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__3407\ : Span12Mux_h
    port map (
            O => \N__20389\,
            I => \N__20386\
        );

    \I__3406\ : Odrv12
    port map (
            O => \N__20386\,
            I => \this_ppu.oam_cache.mem_0\
        );

    \I__3405\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__20380\,
            I => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\
        );

    \I__3403\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20371\
        );

    \I__3401\ : Span4Mux_h
    port map (
            O => \N__20371\,
            I => \N__20368\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__20368\,
            I => \M_this_map_ram_read_data_0\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__20365\,
            I => \N__20359\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__20364\,
            I => \N__20356\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__20363\,
            I => \N__20352\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__20362\,
            I => \N__20347\
        );

    \I__3395\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20343\
        );

    \I__3394\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20339\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__20355\,
            I => \N__20336\
        );

    \I__3392\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20332\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__20351\,
            I => \N__20329\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__20350\,
            I => \N__20326\
        );

    \I__3389\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20322\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__20346\,
            I => \N__20319\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__20343\,
            I => \N__20316\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__20342\,
            I => \N__20313\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__20339\,
            I => \N__20309\
        );

    \I__3384\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20306\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__20335\,
            I => \N__20303\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__20332\,
            I => \N__20299\
        );

    \I__3381\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20296\
        );

    \I__3380\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20293\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N__20290\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__20322\,
            I => \N__20287\
        );

    \I__3377\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20284\
        );

    \I__3376\ : Span4Mux_v
    port map (
            O => \N__20316\,
            I => \N__20281\
        );

    \I__3375\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20278\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__20312\,
            I => \N__20275\
        );

    \I__3373\ : Span4Mux_h
    port map (
            O => \N__20309\,
            I => \N__20269\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20269\
        );

    \I__3371\ : InMux
    port map (
            O => \N__20303\,
            I => \N__20266\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__20302\,
            I => \N__20263\
        );

    \I__3369\ : Span4Mux_h
    port map (
            O => \N__20299\,
            I => \N__20257\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__20296\,
            I => \N__20257\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__20293\,
            I => \N__20254\
        );

    \I__3366\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20251\
        );

    \I__3365\ : Span4Mux_v
    port map (
            O => \N__20287\,
            I => \N__20246\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__20284\,
            I => \N__20246\
        );

    \I__3363\ : Span4Mux_v
    port map (
            O => \N__20281\,
            I => \N__20241\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20241\
        );

    \I__3361\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20238\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N__20235\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__20269\,
            I => \N__20229\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__20266\,
            I => \N__20229\
        );

    \I__3357\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20226\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__20262\,
            I => \N__20223\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__20257\,
            I => \N__20218\
        );

    \I__3354\ : Span4Mux_h
    port map (
            O => \N__20254\,
            I => \N__20218\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__20251\,
            I => \N__20215\
        );

    \I__3352\ : Span4Mux_v
    port map (
            O => \N__20246\,
            I => \N__20208\
        );

    \I__3351\ : Span4Mux_h
    port map (
            O => \N__20241\,
            I => \N__20208\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__20238\,
            I => \N__20208\
        );

    \I__3349\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20205\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__20234\,
            I => \N__20202\
        );

    \I__3347\ : Span4Mux_h
    port map (
            O => \N__20229\,
            I => \N__20197\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__20226\,
            I => \N__20197\
        );

    \I__3345\ : InMux
    port map (
            O => \N__20223\,
            I => \N__20194\
        );

    \I__3344\ : Span4Mux_h
    port map (
            O => \N__20218\,
            I => \N__20191\
        );

    \I__3343\ : Span12Mux_s8_h
    port map (
            O => \N__20215\,
            I => \N__20188\
        );

    \I__3342\ : Span4Mux_v
    port map (
            O => \N__20208\,
            I => \N__20185\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__20205\,
            I => \N__20182\
        );

    \I__3340\ : InMux
    port map (
            O => \N__20202\,
            I => \N__20179\
        );

    \I__3339\ : Span4Mux_v
    port map (
            O => \N__20197\,
            I => \N__20174\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__20194\,
            I => \N__20174\
        );

    \I__3337\ : Span4Mux_h
    port map (
            O => \N__20191\,
            I => \N__20171\
        );

    \I__3336\ : Span12Mux_h
    port map (
            O => \N__20188\,
            I => \N__20168\
        );

    \I__3335\ : Sp12to4
    port map (
            O => \N__20185\,
            I => \N__20163\
        );

    \I__3334\ : Span12Mux_s8_h
    port map (
            O => \N__20182\,
            I => \N__20163\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__20179\,
            I => \N__20160\
        );

    \I__3332\ : Span4Mux_v
    port map (
            O => \N__20174\,
            I => \N__20157\
        );

    \I__3331\ : Span4Mux_h
    port map (
            O => \N__20171\,
            I => \N__20154\
        );

    \I__3330\ : Span12Mux_v
    port map (
            O => \N__20168\,
            I => \N__20147\
        );

    \I__3329\ : Span12Mux_h
    port map (
            O => \N__20163\,
            I => \N__20147\
        );

    \I__3328\ : Span12Mux_s11_h
    port map (
            O => \N__20160\,
            I => \N__20147\
        );

    \I__3327\ : Span4Mux_h
    port map (
            O => \N__20157\,
            I => \N__20144\
        );

    \I__3326\ : Odrv4
    port map (
            O => \N__20154\,
            I => \M_this_ppu_spr_addr_6\
        );

    \I__3325\ : Odrv12
    port map (
            O => \N__20147\,
            I => \M_this_ppu_spr_addr_6\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__20144\,
            I => \M_this_ppu_spr_addr_6\
        );

    \I__3323\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20134\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20131\
        );

    \I__3321\ : Span4Mux_v
    port map (
            O => \N__20131\,
            I => \N__20128\
        );

    \I__3320\ : Span4Mux_h
    port map (
            O => \N__20128\,
            I => \N__20125\
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__20125\,
            I => \this_spr_ram.mem_out_bus4_2\
        );

    \I__3318\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20119\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__20119\,
            I => \N__20116\
        );

    \I__3316\ : Span12Mux_v
    port map (
            O => \N__20116\,
            I => \N__20113\
        );

    \I__3315\ : Span12Mux_h
    port map (
            O => \N__20113\,
            I => \N__20110\
        );

    \I__3314\ : Odrv12
    port map (
            O => \N__20110\,
            I => \this_spr_ram.mem_out_bus0_2\
        );

    \I__3313\ : CEMux
    port map (
            O => \N__20107\,
            I => \N__20104\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20101\
        );

    \I__3311\ : Span4Mux_h
    port map (
            O => \N__20101\,
            I => \N__20098\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__20098\,
            I => \N__20095\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__20095\,
            I => \M_state_q_RNIQER3C_9\
        );

    \I__3308\ : InMux
    port map (
            O => \N__20092\,
            I => \N__20089\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__20089\,
            I => \N__20086\
        );

    \I__3306\ : Span4Mux_v
    port map (
            O => \N__20086\,
            I => \N__20083\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__20083\,
            I => \N__20080\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__20080\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__3303\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20058\
        );

    \I__3302\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20058\
        );

    \I__3301\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20048\
        );

    \I__3300\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20048\
        );

    \I__3299\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20048\
        );

    \I__3298\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20048\
        );

    \I__3297\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20043\
        );

    \I__3296\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20043\
        );

    \I__3295\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20038\
        );

    \I__3294\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20038\
        );

    \I__3293\ : InMux
    port map (
            O => \N__20067\,
            I => \N__20031\
        );

    \I__3292\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20031\
        );

    \I__3291\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20031\
        );

    \I__3290\ : InMux
    port map (
            O => \N__20064\,
            I => \N__20026\
        );

    \I__3289\ : CEMux
    port map (
            O => \N__20063\,
            I => \N__20021\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__20058\,
            I => \N__20018\
        );

    \I__3287\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20015\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__20048\,
            I => \N__20012\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__20007\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__20038\,
            I => \N__20007\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__20003\
        );

    \I__3282\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20000\
        );

    \I__3281\ : InMux
    port map (
            O => \N__20029\,
            I => \N__19997\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__20026\,
            I => \N__19994\
        );

    \I__3279\ : InMux
    port map (
            O => \N__20025\,
            I => \N__19991\
        );

    \I__3278\ : InMux
    port map (
            O => \N__20024\,
            I => \N__19988\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__19984\
        );

    \I__3276\ : Span4Mux_h
    port map (
            O => \N__20018\,
            I => \N__19981\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__19974\
        );

    \I__3274\ : Span4Mux_v
    port map (
            O => \N__20012\,
            I => \N__19974\
        );

    \I__3273\ : Span4Mux_h
    port map (
            O => \N__20007\,
            I => \N__19974\
        );

    \I__3272\ : InMux
    port map (
            O => \N__20006\,
            I => \N__19971\
        );

    \I__3271\ : Span4Mux_v
    port map (
            O => \N__20003\,
            I => \N__19966\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__20000\,
            I => \N__19966\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__19997\,
            I => \N__19959\
        );

    \I__3268\ : Span4Mux_v
    port map (
            O => \N__19994\,
            I => \N__19959\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__19991\,
            I => \N__19959\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19956\
        );

    \I__3265\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19952\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__19984\,
            I => \N__19947\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__19981\,
            I => \N__19947\
        );

    \I__3262\ : Span4Mux_v
    port map (
            O => \N__19974\,
            I => \N__19944\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__19971\,
            I => \N__19941\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__19966\,
            I => \N__19938\
        );

    \I__3259\ : Span4Mux_h
    port map (
            O => \N__19959\,
            I => \N__19935\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__19956\,
            I => \N__19932\
        );

    \I__3257\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19929\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19926\
        );

    \I__3255\ : Span4Mux_v
    port map (
            O => \N__19947\,
            I => \N__19923\
        );

    \I__3254\ : Span4Mux_h
    port map (
            O => \N__19944\,
            I => \N__19920\
        );

    \I__3253\ : Span12Mux_v
    port map (
            O => \N__19941\,
            I => \N__19917\
        );

    \I__3252\ : Span4Mux_v
    port map (
            O => \N__19938\,
            I => \N__19912\
        );

    \I__3251\ : Span4Mux_h
    port map (
            O => \N__19935\,
            I => \N__19912\
        );

    \I__3250\ : Span4Mux_v
    port map (
            O => \N__19932\,
            I => \N__19909\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__19929\,
            I => \this_vga_signals.GZ0Z_406\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__19926\,
            I => \this_vga_signals.GZ0Z_406\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__19923\,
            I => \this_vga_signals.GZ0Z_406\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__19920\,
            I => \this_vga_signals.GZ0Z_406\
        );

    \I__3245\ : Odrv12
    port map (
            O => \N__19917\,
            I => \this_vga_signals.GZ0Z_406\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__19912\,
            I => \this_vga_signals.GZ0Z_406\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__19909\,
            I => \this_vga_signals.GZ0Z_406\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__19894\,
            I => \N__19887\
        );

    \I__3241\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19882\
        );

    \I__3240\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19882\
        );

    \I__3239\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19877\
        );

    \I__3238\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19874\
        );

    \I__3237\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19871\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__19882\,
            I => \N__19867\
        );

    \I__3235\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19864\
        );

    \I__3234\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19861\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19858\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__19874\,
            I => \N__19853\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__19871\,
            I => \N__19853\
        );

    \I__3230\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19850\
        );

    \I__3229\ : Span4Mux_h
    port map (
            O => \N__19867\,
            I => \N__19843\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__19864\,
            I => \N__19843\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__19861\,
            I => \N__19840\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__19858\,
            I => \N__19836\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__19853\,
            I => \N__19833\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__19850\,
            I => \N__19830\
        );

    \I__3223\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19827\
        );

    \I__3222\ : InMux
    port map (
            O => \N__19848\,
            I => \N__19824\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__19843\,
            I => \N__19821\
        );

    \I__3220\ : Span4Mux_v
    port map (
            O => \N__19840\,
            I => \N__19818\
        );

    \I__3219\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19815\
        );

    \I__3218\ : Span4Mux_h
    port map (
            O => \N__19836\,
            I => \N__19808\
        );

    \I__3217\ : Span4Mux_h
    port map (
            O => \N__19833\,
            I => \N__19808\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__19830\,
            I => \N__19808\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__19827\,
            I => \this_vga_signals.N_83_1\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__19824\,
            I => \this_vga_signals.N_83_1\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__19821\,
            I => \this_vga_signals.N_83_1\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__19818\,
            I => \this_vga_signals.N_83_1\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__19815\,
            I => \this_vga_signals.N_83_1\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__19808\,
            I => \this_vga_signals.N_83_1\
        );

    \I__3209\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19790\
        );

    \I__3208\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19785\
        );

    \I__3207\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19785\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__19790\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__19785\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__3204\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__19777\,
            I => \N__19774\
        );

    \I__3202\ : Span4Mux_v
    port map (
            O => \N__19774\,
            I => \N__19771\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__19771\,
            I => \M_this_map_ram_write_data_1\
        );

    \I__3200\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__19765\,
            I => \N__19762\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__19762\,
            I => \M_this_map_ram_write_data_2\
        );

    \I__3197\ : InMux
    port map (
            O => \N__19759\,
            I => \N__19756\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__19756\,
            I => \N__19753\
        );

    \I__3195\ : Span4Mux_h
    port map (
            O => \N__19753\,
            I => \N__19750\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__19750\,
            I => \M_this_map_ram_write_data_7\
        );

    \I__3193\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19744\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__3191\ : Span4Mux_h
    port map (
            O => \N__19741\,
            I => \N__19738\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__19738\,
            I => \M_this_map_ram_write_data_5\
        );

    \I__3189\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19732\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__19729\,
            I => \N__19726\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__19726\,
            I => \N__19723\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__19723\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__3184\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19715\
        );

    \I__3183\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19712\
        );

    \I__3182\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19707\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19704\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19701\
        );

    \I__3179\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19698\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__19710\,
            I => \N__19695\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__19707\,
            I => \N__19692\
        );

    \I__3176\ : Span4Mux_v
    port map (
            O => \N__19704\,
            I => \N__19689\
        );

    \I__3175\ : Span4Mux_v
    port map (
            O => \N__19701\,
            I => \N__19684\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19684\
        );

    \I__3173\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19681\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__19692\,
            I => \N__19678\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__19689\,
            I => \N__19671\
        );

    \I__3170\ : Span4Mux_v
    port map (
            O => \N__19684\,
            I => \N__19671\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19671\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__19678\,
            I => \N_825_0\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__19671\,
            I => \N_825_0\
        );

    \I__3166\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19660\
        );

    \I__3165\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19660\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__19660\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__3163\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19654\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__19654\,
            I => \N__19651\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__19651\,
            I => \N__19648\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__19648\,
            I => \M_this_map_ram_write_data_0\
        );

    \I__3159\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19642\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__19642\,
            I => \N__19639\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__19639\,
            I => \M_this_map_ram_write_data_3\
        );

    \I__3156\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19633\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__19633\,
            I => \N__19630\
        );

    \I__3154\ : Span4Mux_h
    port map (
            O => \N__19630\,
            I => \N__19627\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__19627\,
            I => \M_this_map_ram_write_data_4\
        );

    \I__3152\ : IoInMux
    port map (
            O => \N__19624\,
            I => \N__19621\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19616\
        );

    \I__3150\ : IoInMux
    port map (
            O => \N__19620\,
            I => \N__19613\
        );

    \I__3149\ : IoInMux
    port map (
            O => \N__19619\,
            I => \N__19610\
        );

    \I__3148\ : IoSpan4Mux
    port map (
            O => \N__19616\,
            I => \N__19600\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__19613\,
            I => \N__19600\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19600\
        );

    \I__3145\ : IoInMux
    port map (
            O => \N__19609\,
            I => \N__19597\
        );

    \I__3144\ : IoInMux
    port map (
            O => \N__19608\,
            I => \N__19594\
        );

    \I__3143\ : IoInMux
    port map (
            O => \N__19607\,
            I => \N__19590\
        );

    \I__3142\ : IoSpan4Mux
    port map (
            O => \N__19600\,
            I => \N__19580\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__19597\,
            I => \N__19580\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19577\
        );

    \I__3139\ : IoInMux
    port map (
            O => \N__19593\,
            I => \N__19574\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__19590\,
            I => \N__19571\
        );

    \I__3137\ : IoInMux
    port map (
            O => \N__19589\,
            I => \N__19568\
        );

    \I__3136\ : IoInMux
    port map (
            O => \N__19588\,
            I => \N__19565\
        );

    \I__3135\ : IoInMux
    port map (
            O => \N__19587\,
            I => \N__19561\
        );

    \I__3134\ : IoInMux
    port map (
            O => \N__19586\,
            I => \N__19558\
        );

    \I__3133\ : IoInMux
    port map (
            O => \N__19585\,
            I => \N__19555\
        );

    \I__3132\ : IoSpan4Mux
    port map (
            O => \N__19580\,
            I => \N__19547\
        );

    \I__3131\ : IoSpan4Mux
    port map (
            O => \N__19577\,
            I => \N__19547\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__19574\,
            I => \N__19547\
        );

    \I__3129\ : IoSpan4Mux
    port map (
            O => \N__19571\,
            I => \N__19540\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19540\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__19565\,
            I => \N__19540\
        );

    \I__3126\ : IoInMux
    port map (
            O => \N__19564\,
            I => \N__19537\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__19561\,
            I => \N__19531\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19531\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__19555\,
            I => \N__19528\
        );

    \I__3122\ : IoInMux
    port map (
            O => \N__19554\,
            I => \N__19525\
        );

    \I__3121\ : IoSpan4Mux
    port map (
            O => \N__19547\,
            I => \N__19522\
        );

    \I__3120\ : IoSpan4Mux
    port map (
            O => \N__19540\,
            I => \N__19516\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__19537\,
            I => \N__19516\
        );

    \I__3118\ : IoInMux
    port map (
            O => \N__19536\,
            I => \N__19513\
        );

    \I__3117\ : IoSpan4Mux
    port map (
            O => \N__19531\,
            I => \N__19510\
        );

    \I__3116\ : IoSpan4Mux
    port map (
            O => \N__19528\,
            I => \N__19505\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__19525\,
            I => \N__19505\
        );

    \I__3114\ : Span4Mux_s3_v
    port map (
            O => \N__19522\,
            I => \N__19502\
        );

    \I__3113\ : IoInMux
    port map (
            O => \N__19521\,
            I => \N__19499\
        );

    \I__3112\ : Sp12to4
    port map (
            O => \N__19516\,
            I => \N__19494\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19494\
        );

    \I__3110\ : IoSpan4Mux
    port map (
            O => \N__19510\,
            I => \N__19489\
        );

    \I__3109\ : IoSpan4Mux
    port map (
            O => \N__19505\,
            I => \N__19489\
        );

    \I__3108\ : Sp12to4
    port map (
            O => \N__19502\,
            I => \N__19483\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__19499\,
            I => \N__19483\
        );

    \I__3106\ : Span12Mux_s9_h
    port map (
            O => \N__19494\,
            I => \N__19480\
        );

    \I__3105\ : Sp12to4
    port map (
            O => \N__19489\,
            I => \N__19477\
        );

    \I__3104\ : IoInMux
    port map (
            O => \N__19488\,
            I => \N__19474\
        );

    \I__3103\ : Span12Mux_s10_v
    port map (
            O => \N__19483\,
            I => \N__19471\
        );

    \I__3102\ : Span12Mux_v
    port map (
            O => \N__19480\,
            I => \N__19466\
        );

    \I__3101\ : Span12Mux_s9_h
    port map (
            O => \N__19477\,
            I => \N__19466\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19463\
        );

    \I__3099\ : Span12Mux_v
    port map (
            O => \N__19471\,
            I => \N__19460\
        );

    \I__3098\ : Span12Mux_h
    port map (
            O => \N__19466\,
            I => \N__19455\
        );

    \I__3097\ : Span12Mux_s10_h
    port map (
            O => \N__19463\,
            I => \N__19455\
        );

    \I__3096\ : Odrv12
    port map (
            O => \N__19460\,
            I => dma_0_i
        );

    \I__3095\ : Odrv12
    port map (
            O => \N__19455\,
            I => dma_0_i
        );

    \I__3094\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19446\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__19449\,
            I => \N__19442\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__19446\,
            I => \N__19439\
        );

    \I__3091\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19436\
        );

    \I__3090\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19433\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__19439\,
            I => \N__19428\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__19436\,
            I => \N__19428\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__19433\,
            I => \N__19425\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__19428\,
            I => \N__19420\
        );

    \I__3085\ : Span4Mux_v
    port map (
            O => \N__19425\,
            I => \N__19420\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__19420\,
            I => \this_vga_signals.N_819_0\
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__19417\,
            I => \this_vga_signals.N_827_0_cascade_\
        );

    \I__3082\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__19411\,
            I => \this_vga_signals.N_826_0\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__19408\,
            I => \N__19405\
        );

    \I__3079\ : CascadeBuf
    port map (
            O => \N__19405\,
            I => \N__19402\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__3077\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19395\
        );

    \I__3076\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19392\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__19395\,
            I => \N__19389\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__19392\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__19389\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__3072\ : InMux
    port map (
            O => \N__19384\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__19381\,
            I => \N__19378\
        );

    \I__3070\ : CascadeBuf
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__19375\,
            I => \N__19372\
        );

    \I__3068\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19369\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19365\
        );

    \I__3066\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19362\
        );

    \I__3065\ : Span4Mux_h
    port map (
            O => \N__19365\,
            I => \N__19359\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__19362\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__19359\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__3062\ : InMux
    port map (
            O => \N__19354\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__19351\,
            I => \N__19348\
        );

    \I__3060\ : CascadeBuf
    port map (
            O => \N__19348\,
            I => \N__19345\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__19345\,
            I => \N__19342\
        );

    \I__3058\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19338\
        );

    \I__3057\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19335\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__19338\,
            I => \N__19332\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__19335\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__19332\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__3053\ : InMux
    port map (
            O => \N__19327\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__3051\ : CascadeBuf
    port map (
            O => \N__19321\,
            I => \N__19318\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__19318\,
            I => \N__19315\
        );

    \I__3049\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19311\
        );

    \I__3048\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19308\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__19311\,
            I => \N__19305\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__19308\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__19305\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__3044\ : InMux
    port map (
            O => \N__19300\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__19297\,
            I => \N__19294\
        );

    \I__3042\ : CascadeBuf
    port map (
            O => \N__19294\,
            I => \N__19291\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__19291\,
            I => \N__19288\
        );

    \I__3040\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19285\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__19285\,
            I => \N__19281\
        );

    \I__3038\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19278\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__19281\,
            I => \N__19275\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__19278\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__19275\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__3034\ : InMux
    port map (
            O => \N__19270\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__3032\ : CascadeBuf
    port map (
            O => \N__19264\,
            I => \N__19261\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__19261\,
            I => \N__19258\
        );

    \I__3030\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19255\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__19255\,
            I => \N__19251\
        );

    \I__3028\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19248\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__19251\,
            I => \N__19245\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__19248\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__19245\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__3024\ : InMux
    port map (
            O => \N__19240\,
            I => \bfn_9_22_0_\
        );

    \I__3023\ : InMux
    port map (
            O => \N__19237\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__19234\,
            I => \N__19231\
        );

    \I__3021\ : CascadeBuf
    port map (
            O => \N__19231\,
            I => \N__19228\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__19228\,
            I => \N__19225\
        );

    \I__3019\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19221\
        );

    \I__3018\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19218\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__19221\,
            I => \N__19215\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__19218\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__19215\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__3014\ : IoInMux
    port map (
            O => \N__19210\,
            I => \N__19207\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19204\
        );

    \I__3012\ : IoSpan4Mux
    port map (
            O => \N__19204\,
            I => \N__19201\
        );

    \I__3011\ : IoSpan4Mux
    port map (
            O => \N__19201\,
            I => \N__19198\
        );

    \I__3010\ : Span4Mux_s3_v
    port map (
            O => \N__19198\,
            I => \N__19195\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__19195\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__3007\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19186\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__19186\,
            I => \this_vga_signals.M_lcounter_q_3_i_o2_0_1\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__19183\,
            I => \N__19180\
        );

    \I__3004\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19175\
        );

    \I__3003\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19172\
        );

    \I__3002\ : InMux
    port map (
            O => \N__19178\,
            I => \N__19169\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__19175\,
            I => \this_vga_signals.pixel_clk_i\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__19172\,
            I => \this_vga_signals.pixel_clk_i\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__19169\,
            I => \this_vga_signals.pixel_clk_i\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__19162\,
            I => \this_vga_signals.N_83_1_cascade_\
        );

    \I__2997\ : InMux
    port map (
            O => \N__19159\,
            I => \N__19153\
        );

    \I__2996\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19153\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__19153\,
            I => \this_vga_signals.N_2_0\
        );

    \I__2994\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19147\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__19147\,
            I => \N__19143\
        );

    \I__2992\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19140\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__19143\,
            I => \this_vga_signals.M_pcounter_q_i_2_1\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__19140\,
            I => \this_vga_signals.M_pcounter_q_i_2_1\
        );

    \I__2989\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19129\
        );

    \I__2988\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19126\
        );

    \I__2987\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19123\
        );

    \I__2986\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19120\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__19129\,
            I => \N__19117\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__19126\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__19123\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__19120\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__19117\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2980\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__19102\,
            I => \this_vga_signals.M_pcounter_q_0Z0Z_1\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__19099\,
            I => \N__19093\
        );

    \I__2976\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19088\
        );

    \I__2975\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19085\
        );

    \I__2974\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19082\
        );

    \I__2973\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19079\
        );

    \I__2972\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19076\
        );

    \I__2971\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19073\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__19088\,
            I => \N__19070\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__19085\,
            I => \N__19066\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__19082\,
            I => \N__19063\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__19079\,
            I => \N__19056\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19056\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__19073\,
            I => \N__19056\
        );

    \I__2964\ : Span4Mux_v
    port map (
            O => \N__19070\,
            I => \N__19050\
        );

    \I__2963\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19047\
        );

    \I__2962\ : Span4Mux_h
    port map (
            O => \N__19066\,
            I => \N__19044\
        );

    \I__2961\ : Span4Mux_h
    port map (
            O => \N__19063\,
            I => \N__19039\
        );

    \I__2960\ : Span4Mux_v
    port map (
            O => \N__19056\,
            I => \N__19039\
        );

    \I__2959\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19036\
        );

    \I__2958\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19033\
        );

    \I__2957\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19030\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__19050\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__19047\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__19044\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__19039\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__19036\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__19033\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__19030\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__2949\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19010\
        );

    \I__2948\ : InMux
    port map (
            O => \N__19014\,
            I => \N__19005\
        );

    \I__2947\ : InMux
    port map (
            O => \N__19013\,
            I => \N__19002\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__19010\,
            I => \N__18998\
        );

    \I__2945\ : InMux
    port map (
            O => \N__19009\,
            I => \N__18992\
        );

    \I__2944\ : InMux
    port map (
            O => \N__19008\,
            I => \N__18992\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__19005\,
            I => \N__18983\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__19002\,
            I => \N__18980\
        );

    \I__2941\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18977\
        );

    \I__2940\ : Span4Mux_h
    port map (
            O => \N__18998\,
            I => \N__18974\
        );

    \I__2939\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18971\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__18992\,
            I => \N__18968\
        );

    \I__2937\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18965\
        );

    \I__2936\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18954\
        );

    \I__2935\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18954\
        );

    \I__2934\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18954\
        );

    \I__2933\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18954\
        );

    \I__2932\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18954\
        );

    \I__2931\ : Odrv12
    port map (
            O => \N__18983\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2930\ : Odrv4
    port map (
            O => \N__18980\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__18977\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__18974\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__18971\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__18968\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__18965\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__18954\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__2923\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18933\
        );

    \I__2922\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18929\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__18933\,
            I => \N__18925\
        );

    \I__2920\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18921\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__18929\,
            I => \N__18914\
        );

    \I__2918\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18911\
        );

    \I__2917\ : Span4Mux_v
    port map (
            O => \N__18925\,
            I => \N__18908\
        );

    \I__2916\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18905\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18902\
        );

    \I__2914\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18899\
        );

    \I__2913\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18896\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__18918\,
            I => \N__18893\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__18917\,
            I => \N__18890\
        );

    \I__2910\ : Span4Mux_v
    port map (
            O => \N__18914\,
            I => \N__18887\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__18911\,
            I => \N__18884\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__18908\,
            I => \N__18873\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__18905\,
            I => \N__18873\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__18902\,
            I => \N__18873\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__18899\,
            I => \N__18873\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__18896\,
            I => \N__18873\
        );

    \I__2903\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18870\
        );

    \I__2902\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18867\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__18887\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2900\ : Odrv12
    port map (
            O => \N__18884\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__18873\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__18870\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__18867\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__18856\,
            I => \this_vga_signals.N_809_0_cascade_\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__18853\,
            I => \N__18850\
        );

    \I__2894\ : InMux
    port map (
            O => \N__18850\,
            I => \N__18844\
        );

    \I__2893\ : InMux
    port map (
            O => \N__18849\,
            I => \N__18841\
        );

    \I__2892\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18836\
        );

    \I__2891\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18833\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__18844\,
            I => \N__18828\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__18841\,
            I => \N__18828\
        );

    \I__2888\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18823\
        );

    \I__2887\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18823\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__18836\,
            I => \N__18820\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18816\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__18828\,
            I => \N__18810\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18810\
        );

    \I__2882\ : Span4Mux_v
    port map (
            O => \N__18820\,
            I => \N__18806\
        );

    \I__2881\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18803\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__18816\,
            I => \N__18800\
        );

    \I__2879\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18797\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__18810\,
            I => \N__18794\
        );

    \I__2877\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18791\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__18806\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__18803\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__18800\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__18797\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__18794\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__18791\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__2869\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18772\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__18772\,
            I => \N__18769\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__18769\,
            I => \N__18766\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__18766\,
            I => \N__18763\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__18763\,
            I => \N_34_0\
        );

    \I__2864\ : IoInMux
    port map (
            O => \N__18760\,
            I => \N__18757\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__18757\,
            I => \N__18754\
        );

    \I__2862\ : Span4Mux_s2_h
    port map (
            O => \N__18754\,
            I => \N__18751\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__18751\,
            I => \N__18748\
        );

    \I__2860\ : Span4Mux_h
    port map (
            O => \N__18748\,
            I => \N__18745\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__18745\,
            I => port_nmib_1_i
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__18742\,
            I => \N__18739\
        );

    \I__2857\ : CascadeBuf
    port map (
            O => \N__18739\,
            I => \N__18736\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__18736\,
            I => \N__18733\
        );

    \I__2855\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18730\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__18730\,
            I => \N__18726\
        );

    \I__2853\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18723\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__18726\,
            I => \N__18720\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__18723\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__18720\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__18715\,
            I => \N__18712\
        );

    \I__2848\ : CascadeBuf
    port map (
            O => \N__18712\,
            I => \N__18709\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__18709\,
            I => \N__18706\
        );

    \I__2846\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__18703\,
            I => \N__18699\
        );

    \I__2844\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18696\
        );

    \I__2843\ : Span4Mux_v
    port map (
            O => \N__18699\,
            I => \N__18693\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__18696\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__18693\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__2840\ : InMux
    port map (
            O => \N__18688\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__2838\ : CascadeBuf
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__18679\,
            I => \N__18676\
        );

    \I__2836\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18673\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__18673\,
            I => \N__18669\
        );

    \I__2834\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18666\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__18669\,
            I => \N__18663\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__18666\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__18663\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__2830\ : InMux
    port map (
            O => \N__18658\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__18655\,
            I => \N__18651\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__18654\,
            I => \N__18647\
        );

    \I__2827\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18641\
        );

    \I__2826\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18637\
        );

    \I__2825\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18632\
        );

    \I__2824\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18632\
        );

    \I__2823\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18629\
        );

    \I__2822\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18626\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18619\
        );

    \I__2820\ : InMux
    port map (
            O => \N__18640\,
            I => \N__18616\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18613\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__18632\,
            I => \N__18608\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__18629\,
            I => \N__18608\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__18626\,
            I => \N__18604\
        );

    \I__2815\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18599\
        );

    \I__2814\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18599\
        );

    \I__2813\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18594\
        );

    \I__2812\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18594\
        );

    \I__2811\ : Span4Mux_v
    port map (
            O => \N__18619\,
            I => \N__18585\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__18616\,
            I => \N__18585\
        );

    \I__2809\ : Span4Mux_v
    port map (
            O => \N__18613\,
            I => \N__18585\
        );

    \I__2808\ : Span4Mux_v
    port map (
            O => \N__18608\,
            I => \N__18585\
        );

    \I__2807\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18582\
        );

    \I__2806\ : Odrv12
    port map (
            O => \N__18604\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__18599\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__18594\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2803\ : Odrv4
    port map (
            O => \N__18585\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__18582\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2801\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18567\
        );

    \I__2800\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18564\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__18567\,
            I => \N__18560\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__18564\,
            I => \N__18557\
        );

    \I__2797\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18554\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__18560\,
            I => \this_vga_signals.mult1_un68_sum_axbxc1\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__18557\,
            I => \this_vga_signals.mult1_un68_sum_axbxc1\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__18554\,
            I => \this_vga_signals.mult1_un68_sum_axbxc1\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__18547\,
            I => \N__18543\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__18546\,
            I => \N__18539\
        );

    \I__2791\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18536\
        );

    \I__2790\ : InMux
    port map (
            O => \N__18542\,
            I => \N__18529\
        );

    \I__2789\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18529\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18520\
        );

    \I__2787\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18517\
        );

    \I__2786\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18514\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__18529\,
            I => \N__18511\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__18528\,
            I => \N__18508\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__18527\,
            I => \N__18504\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__18526\,
            I => \N__18501\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__18525\,
            I => \N__18497\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__18524\,
            I => \N__18494\
        );

    \I__2779\ : InMux
    port map (
            O => \N__18523\,
            I => \N__18491\
        );

    \I__2778\ : Span12Mux_h
    port map (
            O => \N__18520\,
            I => \N__18488\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__18517\,
            I => \N__18481\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__18514\,
            I => \N__18481\
        );

    \I__2775\ : Span4Mux_h
    port map (
            O => \N__18511\,
            I => \N__18481\
        );

    \I__2774\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18478\
        );

    \I__2773\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18473\
        );

    \I__2772\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18473\
        );

    \I__2771\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18470\
        );

    \I__2770\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18463\
        );

    \I__2769\ : InMux
    port map (
            O => \N__18497\,
            I => \N__18463\
        );

    \I__2768\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18463\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__18491\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__18488\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__18481\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__18478\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__18473\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__18470\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__18463\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2760\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18445\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__18445\,
            I => \N__18438\
        );

    \I__2758\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18435\
        );

    \I__2757\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18430\
        );

    \I__2756\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18430\
        );

    \I__2755\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18424\
        );

    \I__2754\ : Span4Mux_v
    port map (
            O => \N__18438\,
            I => \N__18417\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__18435\,
            I => \N__18417\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__18430\,
            I => \N__18417\
        );

    \I__2751\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18412\
        );

    \I__2750\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18412\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18409\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__18424\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__18417\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__18412\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18409\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__2744\ : InMux
    port map (
            O => \N__18400\,
            I => \N__18394\
        );

    \I__2743\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18390\
        );

    \I__2742\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18385\
        );

    \I__2741\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18385\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__18394\,
            I => \N__18380\
        );

    \I__2739\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18377\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__18390\,
            I => \N__18370\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__18385\,
            I => \N__18370\
        );

    \I__2736\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18365\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18365\
        );

    \I__2734\ : Span4Mux_h
    port map (
            O => \N__18380\,
            I => \N__18359\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__18377\,
            I => \N__18359\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18356\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18353\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__18370\,
            I => \N__18348\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__18365\,
            I => \N__18348\
        );

    \I__2728\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18345\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__18359\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18356\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__18353\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__18348\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__18345\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__18334\,
            I => \this_vga_signals.if_N_8_i_cascade_\
        );

    \I__2721\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18326\
        );

    \I__2720\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18321\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__18329\,
            I => \N__18318\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__18326\,
            I => \N__18314\
        );

    \I__2717\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18309\
        );

    \I__2716\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18309\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__18321\,
            I => \N__18306\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18301\
        );

    \I__2713\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18301\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__18314\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__18309\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2710\ : Odrv12
    port map (
            O => \N__18306\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__18301\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2708\ : InMux
    port map (
            O => \N__18292\,
            I => \N__18289\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__18289\,
            I => \this_vga_signals.if_N_9_1\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__18286\,
            I => \this_vga_signals.M_pcounter_q_3_1_cascade_\
        );

    \I__2705\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18278\
        );

    \I__2704\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18273\
        );

    \I__2703\ : InMux
    port map (
            O => \N__18281\,
            I => \N__18273\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__18278\,
            I => \this_vga_signals.N_3_0\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__18273\,
            I => \this_vga_signals.N_3_0\
        );

    \I__2700\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18264\
        );

    \I__2699\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18261\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__18264\,
            I => \N__18255\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__18261\,
            I => \N__18255\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__18260\,
            I => \N__18252\
        );

    \I__2695\ : Span4Mux_v
    port map (
            O => \N__18255\,
            I => \N__18248\
        );

    \I__2694\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18243\
        );

    \I__2693\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18243\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__18248\,
            I => \this_vga_signals.SUM_3_i_0_0\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__18243\,
            I => \this_vga_signals.SUM_3_i_0_0\
        );

    \I__2690\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18235\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__18235\,
            I => \N__18230\
        );

    \I__2688\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18225\
        );

    \I__2687\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18225\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__18230\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__18225\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\
        );

    \I__2684\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18214\
        );

    \I__2682\ : Odrv12
    port map (
            O => \N__18214\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__18211\,
            I => \N__18205\
        );

    \I__2680\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18201\
        );

    \I__2679\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18198\
        );

    \I__2678\ : InMux
    port map (
            O => \N__18208\,
            I => \N__18191\
        );

    \I__2677\ : InMux
    port map (
            O => \N__18205\,
            I => \N__18191\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__18204\,
            I => \N__18188\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__18201\,
            I => \N__18182\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__18198\,
            I => \N__18179\
        );

    \I__2673\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18176\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18173\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__18191\,
            I => \N__18170\
        );

    \I__2670\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18167\
        );

    \I__2669\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18160\
        );

    \I__2668\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18160\
        );

    \I__2667\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18160\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__18182\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__18179\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__18176\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__18173\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__18170\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__18167\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__18160\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__18145\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\
        );

    \I__2658\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18137\
        );

    \I__2657\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18134\
        );

    \I__2656\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18130\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__18137\,
            I => \N__18124\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__18134\,
            I => \N__18121\
        );

    \I__2653\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18118\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__18130\,
            I => \N__18109\
        );

    \I__2651\ : InMux
    port map (
            O => \N__18129\,
            I => \N__18106\
        );

    \I__2650\ : InMux
    port map (
            O => \N__18128\,
            I => \N__18103\
        );

    \I__2649\ : InMux
    port map (
            O => \N__18127\,
            I => \N__18100\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__18124\,
            I => \N__18093\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__18121\,
            I => \N__18093\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__18118\,
            I => \N__18093\
        );

    \I__2645\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18086\
        );

    \I__2644\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18086\
        );

    \I__2643\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18086\
        );

    \I__2642\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18079\
        );

    \I__2641\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18079\
        );

    \I__2640\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18079\
        );

    \I__2639\ : Odrv12
    port map (
            O => \N__18109\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__18106\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__18103\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__18100\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__18093\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__18086\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__18079\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__2632\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18061\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__18061\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_1_0\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__18058\,
            I => \N__18053\
        );

    \I__2629\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18040\
        );

    \I__2628\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18040\
        );

    \I__2627\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18040\
        );

    \I__2626\ : InMux
    port map (
            O => \N__18052\,
            I => \N__18040\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18037\
        );

    \I__2624\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18034\
        );

    \I__2623\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18031\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__18040\,
            I => \N__18024\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__18037\,
            I => \N__18024\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__18034\,
            I => \N__18024\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__18031\,
            I => \N_28_0\
        );

    \I__2618\ : Odrv12
    port map (
            O => \N__18024\,
            I => \N_28_0\
        );

    \I__2617\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18016\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__18016\,
            I => \this_vga_signals.M_hcounter_d7lt7_0\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__18013\,
            I => \N__18010\
        );

    \I__2614\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18007\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__18007\,
            I => \N__18004\
        );

    \I__2612\ : Span4Mux_s2_v
    port map (
            O => \N__18004\,
            I => \N__18001\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__18001\,
            I => \M_this_vga_signals_address_5\
        );

    \I__2610\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17987\
        );

    \I__2609\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17987\
        );

    \I__2608\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17987\
        );

    \I__2607\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17984\
        );

    \I__2606\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17981\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__17987\,
            I => \N__17978\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__17984\,
            I => \N__17973\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__17981\,
            I => \N__17973\
        );

    \I__2602\ : Span4Mux_h
    port map (
            O => \N__17978\,
            I => \N__17970\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__17973\,
            I => \N__17967\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__17970\,
            I => \M_this_vram_read_data_2\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__17967\,
            I => \M_this_vram_read_data_2\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__17962\,
            I => \N__17957\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__17961\,
            I => \N__17953\
        );

    \I__2596\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17949\
        );

    \I__2595\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17944\
        );

    \I__2594\ : InMux
    port map (
            O => \N__17956\,
            I => \N__17944\
        );

    \I__2593\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17940\
        );

    \I__2592\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17937\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__17949\,
            I => \N__17934\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__17944\,
            I => \N__17931\
        );

    \I__2589\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17928\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__17940\,
            I => \N__17925\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__17937\,
            I => \N__17922\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__17934\,
            I => \N__17919\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__17931\,
            I => \N__17912\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__17928\,
            I => \N__17912\
        );

    \I__2583\ : Span4Mux_h
    port map (
            O => \N__17925\,
            I => \N__17912\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__17922\,
            I => \N__17909\
        );

    \I__2581\ : Odrv4
    port map (
            O => \N__17919\,
            I => \M_this_vram_read_data_1\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__17912\,
            I => \M_this_vram_read_data_1\
        );

    \I__2579\ : Odrv4
    port map (
            O => \N__17909\,
            I => \M_this_vram_read_data_1\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__17902\,
            I => \N__17898\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__17901\,
            I => \N__17894\
        );

    \I__2576\ : InMux
    port map (
            O => \N__17898\,
            I => \N__17888\
        );

    \I__2575\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17885\
        );

    \I__2574\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17882\
        );

    \I__2573\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17875\
        );

    \I__2572\ : InMux
    port map (
            O => \N__17892\,
            I => \N__17875\
        );

    \I__2571\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17875\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__17888\,
            I => \N__17866\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__17885\,
            I => \N__17866\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__17882\,
            I => \N__17866\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__17875\,
            I => \N__17866\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__17866\,
            I => \N__17863\
        );

    \I__2565\ : Span4Mux_h
    port map (
            O => \N__17863\,
            I => \N__17860\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__17860\,
            I => \M_this_vram_read_data_0\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__17857\,
            I => \N__17854\
        );

    \I__2562\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17847\
        );

    \I__2561\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17847\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__17852\,
            I => \N__17843\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17838\
        );

    \I__2558\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17835\
        );

    \I__2557\ : InMux
    port map (
            O => \N__17843\,
            I => \N__17832\
        );

    \I__2556\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17829\
        );

    \I__2555\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17826\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__17838\,
            I => \N__17823\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__17835\,
            I => \N__17814\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__17832\,
            I => \N__17814\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__17829\,
            I => \N__17814\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__17826\,
            I => \N__17814\
        );

    \I__2549\ : Span4Mux_h
    port map (
            O => \N__17823\,
            I => \N__17809\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__17814\,
            I => \N__17809\
        );

    \I__2547\ : Sp12to4
    port map (
            O => \N__17809\,
            I => \N__17806\
        );

    \I__2546\ : Odrv12
    port map (
            O => \N__17806\,
            I => \M_this_vram_read_data_3\
        );

    \I__2545\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17800\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__17800\,
            I => \N__17797\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__17797\,
            I => \N__17794\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__17794\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__17791\,
            I => \this_vga_signals.N_2_8_0_cascade_\
        );

    \I__2540\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17785\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__17785\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_2_am\
        );

    \I__2538\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17779\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__17779\,
            I => \N__17776\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__17776\,
            I => \this_vga_signals.haddress_1Z0Z_0\
        );

    \I__2535\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17767\
        );

    \I__2534\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17767\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__17767\,
            I => \N__17762\
        );

    \I__2532\ : InMux
    port map (
            O => \N__17766\,
            I => \N__17757\
        );

    \I__2531\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17757\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__17762\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__17757\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__2528\ : InMux
    port map (
            O => \N__17752\,
            I => \N__17749\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__17749\,
            I => \N__17746\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__17746\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__17743\,
            I => \N__17740\
        );

    \I__2524\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17734\
        );

    \I__2523\ : InMux
    port map (
            O => \N__17739\,
            I => \N__17734\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__17734\,
            I => \N__17730\
        );

    \I__2521\ : InMux
    port map (
            O => \N__17733\,
            I => \N__17727\
        );

    \I__2520\ : Span4Mux_h
    port map (
            O => \N__17730\,
            I => \N__17724\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__17727\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__17724\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0\
        );

    \I__2517\ : InMux
    port map (
            O => \N__17719\,
            I => \N__17716\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__17716\,
            I => \N__17712\
        );

    \I__2515\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17709\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__17712\,
            I => \N__17699\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__17709\,
            I => \N__17699\
        );

    \I__2512\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17692\
        );

    \I__2511\ : InMux
    port map (
            O => \N__17707\,
            I => \N__17692\
        );

    \I__2510\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17692\
        );

    \I__2509\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17687\
        );

    \I__2508\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17687\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__17699\,
            I => \N__17682\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17682\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__17687\,
            I => \this_vga_signals.mult1_un61_sum_0_3\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__17682\,
            I => \this_vga_signals.mult1_un61_sum_0_3\
        );

    \I__2503\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17674\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__17674\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_2_bm\
        );

    \I__2501\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17667\
        );

    \I__2500\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17664\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__17667\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__17664\,
            I => \this_vga_signals.mult1_un75_sum_c2_0\
        );

    \I__2497\ : InMux
    port map (
            O => \N__17659\,
            I => \N__17656\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__17656\,
            I => \N__17653\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__17653\,
            I => \this_vga_ramdac.i2_mux\
        );

    \I__2494\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17647\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17639\
        );

    \I__2492\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17634\
        );

    \I__2491\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17634\
        );

    \I__2490\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17627\
        );

    \I__2489\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17627\
        );

    \I__2488\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17627\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__17639\,
            I => \M_pcounter_q_ret_1_RNI4VLK7\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__17634\,
            I => \M_pcounter_q_ret_1_RNI4VLK7\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__17627\,
            I => \M_pcounter_q_ret_1_RNI4VLK7\
        );

    \I__2484\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17613\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__17616\,
            I => \N__17610\
        );

    \I__2481\ : Span12Mux_v
    port map (
            O => \N__17613\,
            I => \N__17607\
        );

    \I__2480\ : InMux
    port map (
            O => \N__17610\,
            I => \N__17604\
        );

    \I__2479\ : Odrv12
    port map (
            O => \N__17607\,
            I => \this_vga_ramdac.N_2688_reto\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__17604\,
            I => \this_vga_ramdac.N_2688_reto\
        );

    \I__2477\ : InMux
    port map (
            O => \N__17599\,
            I => \N__17591\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__17598\,
            I => \N__17587\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__17597\,
            I => \N__17580\
        );

    \I__2474\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17577\
        );

    \I__2473\ : InMux
    port map (
            O => \N__17595\,
            I => \N__17573\
        );

    \I__2472\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17560\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__17591\,
            I => \N__17557\
        );

    \I__2470\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17554\
        );

    \I__2469\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17551\
        );

    \I__2468\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17546\
        );

    \I__2467\ : InMux
    port map (
            O => \N__17585\,
            I => \N__17546\
        );

    \I__2466\ : InMux
    port map (
            O => \N__17584\,
            I => \N__17543\
        );

    \I__2465\ : InMux
    port map (
            O => \N__17583\,
            I => \N__17540\
        );

    \I__2464\ : InMux
    port map (
            O => \N__17580\,
            I => \N__17537\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__17577\,
            I => \N__17534\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__17576\,
            I => \N__17531\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__17573\,
            I => \N__17526\
        );

    \I__2460\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17521\
        );

    \I__2459\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17521\
        );

    \I__2458\ : InMux
    port map (
            O => \N__17570\,
            I => \N__17517\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__17569\,
            I => \N__17513\
        );

    \I__2456\ : InMux
    port map (
            O => \N__17568\,
            I => \N__17503\
        );

    \I__2455\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17503\
        );

    \I__2454\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17503\
        );

    \I__2453\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17503\
        );

    \I__2452\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17498\
        );

    \I__2451\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17498\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__17560\,
            I => \N__17495\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__17557\,
            I => \N__17492\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__17554\,
            I => \N__17485\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__17551\,
            I => \N__17485\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__17546\,
            I => \N__17485\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__17543\,
            I => \N__17482\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__17540\,
            I => \N__17479\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17476\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__17534\,
            I => \N__17472\
        );

    \I__2441\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17467\
        );

    \I__2440\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17467\
        );

    \I__2439\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17464\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__17526\,
            I => \N__17459\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__17521\,
            I => \N__17459\
        );

    \I__2436\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17456\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__17517\,
            I => \N__17453\
        );

    \I__2434\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17446\
        );

    \I__2433\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17446\
        );

    \I__2432\ : InMux
    port map (
            O => \N__17512\,
            I => \N__17446\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__17503\,
            I => \N__17437\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__17498\,
            I => \N__17437\
        );

    \I__2429\ : Span4Mux_h
    port map (
            O => \N__17495\,
            I => \N__17437\
        );

    \I__2428\ : Span4Mux_h
    port map (
            O => \N__17492\,
            I => \N__17437\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__17485\,
            I => \N__17428\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__17482\,
            I => \N__17428\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__17479\,
            I => \N__17428\
        );

    \I__2424\ : Span4Mux_v
    port map (
            O => \N__17476\,
            I => \N__17428\
        );

    \I__2423\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17425\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__17472\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__17467\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__17464\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__17459\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__17456\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__17453\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__17446\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__17437\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__17428\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__17425\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2412\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17400\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__17403\,
            I => \N__17396\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__17400\,
            I => \N__17386\
        );

    \I__2409\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17381\
        );

    \I__2408\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17381\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__17395\,
            I => \N__17376\
        );

    \I__2406\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17372\
        );

    \I__2405\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17369\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17365\
        );

    \I__2403\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17362\
        );

    \I__2402\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17359\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17356\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__17386\,
            I => \N__17351\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17381\,
            I => \N__17351\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__17380\,
            I => \N__17347\
        );

    \I__2397\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17340\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17335\
        );

    \I__2395\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17335\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17330\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__17369\,
            I => \N__17330\
        );

    \I__2392\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17327\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__17365\,
            I => \N__17322\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__17362\,
            I => \N__17319\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17314\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17314\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__17351\,
            I => \N__17311\
        );

    \I__2386\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17306\
        );

    \I__2385\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17306\
        );

    \I__2384\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17301\
        );

    \I__2383\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17301\
        );

    \I__2382\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17298\
        );

    \I__2381\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17295\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17292\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__17335\,
            I => \N__17289\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__17330\,
            I => \N__17284\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__17327\,
            I => \N__17284\
        );

    \I__2376\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17279\
        );

    \I__2375\ : InMux
    port map (
            O => \N__17325\,
            I => \N__17279\
        );

    \I__2374\ : Span4Mux_s1_h
    port map (
            O => \N__17322\,
            I => \N__17270\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__17319\,
            I => \N__17270\
        );

    \I__2372\ : Span4Mux_v
    port map (
            O => \N__17314\,
            I => \N__17270\
        );

    \I__2371\ : Span4Mux_s1_h
    port map (
            O => \N__17311\,
            I => \N__17270\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__17306\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__17301\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__17298\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__17295\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__17292\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__17289\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__17284\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__17279\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__17270\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__17251\,
            I => \N__17248\
        );

    \I__2360\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17245\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17242\
        );

    \I__2358\ : Span4Mux_h
    port map (
            O => \N__17242\,
            I => \N__17239\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__17239\,
            I => \this_vga_signals.g0_6_0_0\
        );

    \I__2356\ : IoInMux
    port map (
            O => \N__17236\,
            I => \N__17233\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__17233\,
            I => \N__17230\
        );

    \I__2354\ : Span4Mux_s3_v
    port map (
            O => \N__17230\,
            I => \N__17227\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__17227\,
            I => \N__17224\
        );

    \I__2352\ : Sp12to4
    port map (
            O => \N__17224\,
            I => \N__17221\
        );

    \I__2351\ : Span12Mux_s5_h
    port map (
            O => \N__17221\,
            I => \N__17218\
        );

    \I__2350\ : Odrv12
    port map (
            O => \N__17218\,
            I => \M_hcounter_q_esr_RNIU8TO_9\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__17215\,
            I => \N__17212\
        );

    \I__2348\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17209\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__17209\,
            I => \M_this_vga_signals_address_2\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__17206\,
            I => \N__17203\
        );

    \I__2345\ : InMux
    port map (
            O => \N__17203\,
            I => \N__17200\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__17200\,
            I => \M_this_vga_signals_address_0\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__17197\,
            I => \N__17194\
        );

    \I__2342\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17191\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__17191\,
            I => \M_this_vga_signals_address_3\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__17188\,
            I => \N__17185\
        );

    \I__2339\ : InMux
    port map (
            O => \N__17185\,
            I => \N__17182\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__17182\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2337\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__2336\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17173\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__17173\,
            I => \N__17170\
        );

    \I__2334\ : Span4Mux_h
    port map (
            O => \N__17170\,
            I => \N__17167\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__17167\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_0\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__17164\,
            I => \N__17161\
        );

    \I__2331\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17158\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__17158\,
            I => \N__17155\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__17155\,
            I => \M_this_vga_signals_address_1\
        );

    \I__2328\ : InMux
    port map (
            O => \N__17152\,
            I => \N__17149\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__17149\,
            I => \this_vga_signals.M_hcounter_d7lt4\
        );

    \I__2326\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17143\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__2324\ : Span4Mux_v
    port map (
            O => \N__17140\,
            I => \N__17136\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__17139\,
            I => \N__17133\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__17136\,
            I => \N__17130\
        );

    \I__2321\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17127\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__17130\,
            I => \this_vga_ramdac.N_2691_reto\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__17127\,
            I => \this_vga_ramdac.N_2691_reto\
        );

    \I__2318\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17119\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__17116\,
            I => \this_vga_ramdac.m16\
        );

    \I__2315\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17110\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__17107\,
            I => \N__17103\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__2311\ : Span4Mux_v
    port map (
            O => \N__17103\,
            I => \N__17097\
        );

    \I__2310\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17094\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__17097\,
            I => \this_vga_ramdac.N_2689_reto\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__17094\,
            I => \this_vga_ramdac.N_2689_reto\
        );

    \I__2307\ : InMux
    port map (
            O => \N__17089\,
            I => \N__17086\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__17086\,
            I => \N__17083\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__17083\,
            I => \this_vga_signals.N_822_0\
        );

    \I__2304\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__17077\,
            I => \N__17074\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__17074\,
            I => \this_vga_signals.M_lcounter_q_3_i_o2_2_1_1\
        );

    \I__2301\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17068\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__17068\,
            I => \N__17065\
        );

    \I__2299\ : Odrv12
    port map (
            O => \N__17065\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__17062\,
            I => \M_pcounter_q_ret_1_RNI4VLK7_cascade_\
        );

    \I__2297\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__17056\,
            I => \N__17053\
        );

    \I__2295\ : Span4Mux_h
    port map (
            O => \N__17053\,
            I => \N__17049\
        );

    \I__2294\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17046\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__17049\,
            I => \this_vga_ramdac.N_2686_reto\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__17046\,
            I => \this_vga_ramdac.N_2686_reto\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__17041\,
            I => \N__17038\
        );

    \I__2290\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17035\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__17035\,
            I => \this_vga_signals.mult1_un82_sum_c3\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__17032\,
            I => \this_vga_signals.d_N_11_cascade_\
        );

    \I__2287\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17026\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__17026\,
            I => \N__17023\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__17023\,
            I => \this_vga_ramdac.m6\
        );

    \I__2284\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17016\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__17019\,
            I => \N__17013\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__17016\,
            I => \N__17010\
        );

    \I__2281\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17007\
        );

    \I__2280\ : Odrv12
    port map (
            O => \N__17010\,
            I => \this_vga_ramdac.N_2687_reto\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__17007\,
            I => \this_vga_ramdac.N_2687_reto\
        );

    \I__2278\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16998\
        );

    \I__2277\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16994\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__16998\,
            I => \N__16989\
        );

    \I__2275\ : InMux
    port map (
            O => \N__16997\,
            I => \N__16986\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__16994\,
            I => \N__16983\
        );

    \I__2273\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16980\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__16992\,
            I => \N__16977\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__16989\,
            I => \N__16973\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__16986\,
            I => \N__16970\
        );

    \I__2269\ : Span4Mux_v
    port map (
            O => \N__16983\,
            I => \N__16965\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__16980\,
            I => \N__16965\
        );

    \I__2267\ : InMux
    port map (
            O => \N__16977\,
            I => \N__16960\
        );

    \I__2266\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16960\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__16973\,
            I => \N__16954\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__16970\,
            I => \N__16954\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__16965\,
            I => \N__16951\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__16960\,
            I => \N__16948\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__16959\,
            I => \N__16945\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__16954\,
            I => \N__16942\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__16951\,
            I => \N__16939\
        );

    \I__2258\ : Span12Mux_s8_v
    port map (
            O => \N__16948\,
            I => \N__16936\
        );

    \I__2257\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16933\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__16942\,
            I => \this_vga_ramdac.N_28_i_reto\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__16939\,
            I => \this_vga_ramdac.N_28_i_reto\
        );

    \I__2254\ : Odrv12
    port map (
            O => \N__16936\,
            I => \this_vga_ramdac.N_28_i_reto\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__16933\,
            I => \this_vga_ramdac.N_28_i_reto\
        );

    \I__2252\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16921\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__16921\,
            I => \N__16918\
        );

    \I__2250\ : Odrv12
    port map (
            O => \N__16918\,
            I => \this_vga_ramdac.m19\
        );

    \I__2249\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16912\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__16912\,
            I => \N__16909\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__16909\,
            I => \N__16905\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__16908\,
            I => \N__16902\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__16905\,
            I => \N__16899\
        );

    \I__2244\ : InMux
    port map (
            O => \N__16902\,
            I => \N__16896\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__16899\,
            I => \this_vga_ramdac.N_2690_reto\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__16896\,
            I => \this_vga_ramdac.N_2690_reto\
        );

    \I__2241\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16886\
        );

    \I__2240\ : InMux
    port map (
            O => \N__16890\,
            I => \N__16881\
        );

    \I__2239\ : InMux
    port map (
            O => \N__16889\,
            I => \N__16881\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__16886\,
            I => \N__16878\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__16881\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__16878\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__16873\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_cascade_\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__16870\,
            I => \N__16866\
        );

    \I__2233\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16861\
        );

    \I__2232\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16861\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__16861\,
            I => \N__16850\
        );

    \I__2230\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16847\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__16859\,
            I => \N__16843\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__16858\,
            I => \N__16837\
        );

    \I__2227\ : InMux
    port map (
            O => \N__16857\,
            I => \N__16833\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__16856\,
            I => \N__16830\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__16855\,
            I => \N__16827\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__16854\,
            I => \N__16824\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__16853\,
            I => \N__16819\
        );

    \I__2222\ : Span4Mux_v
    port map (
            O => \N__16850\,
            I => \N__16815\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__16847\,
            I => \N__16812\
        );

    \I__2220\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16809\
        );

    \I__2219\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16804\
        );

    \I__2218\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16804\
        );

    \I__2217\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16795\
        );

    \I__2216\ : InMux
    port map (
            O => \N__16840\,
            I => \N__16795\
        );

    \I__2215\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16795\
        );

    \I__2214\ : InMux
    port map (
            O => \N__16836\,
            I => \N__16795\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__16833\,
            I => \N__16792\
        );

    \I__2212\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16789\
        );

    \I__2211\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16786\
        );

    \I__2210\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16781\
        );

    \I__2209\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16781\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__16822\,
            I => \N__16775\
        );

    \I__2207\ : InMux
    port map (
            O => \N__16819\,
            I => \N__16771\
        );

    \I__2206\ : InMux
    port map (
            O => \N__16818\,
            I => \N__16768\
        );

    \I__2205\ : Span4Mux_h
    port map (
            O => \N__16815\,
            I => \N__16765\
        );

    \I__2204\ : Span4Mux_h
    port map (
            O => \N__16812\,
            I => \N__16756\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__16809\,
            I => \N__16756\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__16804\,
            I => \N__16756\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__16795\,
            I => \N__16756\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__16792\,
            I => \N__16753\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__16789\,
            I => \N__16746\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__16786\,
            I => \N__16746\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__16781\,
            I => \N__16746\
        );

    \I__2196\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16743\
        );

    \I__2195\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16738\
        );

    \I__2194\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16738\
        );

    \I__2193\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16733\
        );

    \I__2192\ : InMux
    port map (
            O => \N__16774\,
            I => \N__16733\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__16771\,
            I => \N__16728\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__16768\,
            I => \N__16728\
        );

    \I__2189\ : Span4Mux_s0_h
    port map (
            O => \N__16765\,
            I => \N__16723\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__16756\,
            I => \N__16723\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__16753\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__16746\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__16743\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__16738\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__16733\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2182\ : Odrv12
    port map (
            O => \N__16728\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__16723\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2180\ : InMux
    port map (
            O => \N__16708\,
            I => \N__16699\
        );

    \I__2179\ : InMux
    port map (
            O => \N__16707\,
            I => \N__16695\
        );

    \I__2178\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16692\
        );

    \I__2177\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16689\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__16704\,
            I => \N__16683\
        );

    \I__2175\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16675\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16675\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__16699\,
            I => \N__16672\
        );

    \I__2172\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16669\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__16695\,
            I => \N__16666\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__16692\,
            I => \N__16663\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__16689\,
            I => \N__16660\
        );

    \I__2168\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16657\
        );

    \I__2167\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16654\
        );

    \I__2166\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16651\
        );

    \I__2165\ : InMux
    port map (
            O => \N__16683\,
            I => \N__16646\
        );

    \I__2164\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16646\
        );

    \I__2163\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16643\
        );

    \I__2162\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16640\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__16675\,
            I => \N__16633\
        );

    \I__2160\ : Span4Mux_h
    port map (
            O => \N__16672\,
            I => \N__16633\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__16669\,
            I => \N__16633\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__16666\,
            I => \N__16624\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__16663\,
            I => \N__16624\
        );

    \I__2156\ : Span4Mux_v
    port map (
            O => \N__16660\,
            I => \N__16624\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__16657\,
            I => \N__16624\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__16654\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__16651\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__16646\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__16643\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__16640\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__16633\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__16624\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__2147\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16606\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__16606\,
            I => \this_vga_signals.g0_0_2\
        );

    \I__2145\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16598\
        );

    \I__2144\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16595\
        );

    \I__2143\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16587\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__16598\,
            I => \N__16584\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__16595\,
            I => \N__16581\
        );

    \I__2140\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16575\
        );

    \I__2139\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16575\
        );

    \I__2138\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16568\
        );

    \I__2137\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16568\
        );

    \I__2136\ : InMux
    port map (
            O => \N__16590\,
            I => \N__16568\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__16587\,
            I => \N__16558\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__16584\,
            I => \N__16558\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__16581\,
            I => \N__16558\
        );

    \I__2132\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16555\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__16575\,
            I => \N__16550\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__16568\,
            I => \N__16550\
        );

    \I__2129\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16547\
        );

    \I__2128\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16542\
        );

    \I__2127\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16542\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__16558\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__16555\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__16550\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__16547\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__16542\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__16531\,
            I => \N__16528\
        );

    \I__2120\ : InMux
    port map (
            O => \N__16528\,
            I => \N__16525\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__16525\,
            I => \N__16522\
        );

    \I__2118\ : Span4Mux_s2_h
    port map (
            O => \N__16522\,
            I => \N__16519\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__16519\,
            I => \this_vga_signals.g0_0_3_0\
        );

    \I__2116\ : SRMux
    port map (
            O => \N__16516\,
            I => \N__16511\
        );

    \I__2115\ : SRMux
    port map (
            O => \N__16515\,
            I => \N__16508\
        );

    \I__2114\ : SRMux
    port map (
            O => \N__16514\,
            I => \N__16505\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__16511\,
            I => \N__16502\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__16508\,
            I => \N__16499\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16496\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__16502\,
            I => \N__16492\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__16499\,
            I => \N__16487\
        );

    \I__2108\ : Span4Mux_h
    port map (
            O => \N__16496\,
            I => \N__16487\
        );

    \I__2107\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16484\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__16492\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__16487\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__16484\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9\
        );

    \I__2103\ : CEMux
    port map (
            O => \N__16477\,
            I => \N__16474\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__16474\,
            I => \N__16471\
        );

    \I__2101\ : Span4Mux_h
    port map (
            O => \N__16471\,
            I => \N__16468\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__16468\,
            I => \N__16465\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__16465\,
            I => \this_vga_signals.N_935_1\
        );

    \I__2098\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16459\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__16459\,
            I => \N__16456\
        );

    \I__2096\ : Span4Mux_h
    port map (
            O => \N__16456\,
            I => \N__16453\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__16453\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__16450\,
            I => \N__16447\
        );

    \I__2093\ : InMux
    port map (
            O => \N__16447\,
            I => \N__16444\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__16444\,
            I => \this_vga_signals.g0_0_0\
        );

    \I__2091\ : IoInMux
    port map (
            O => \N__16441\,
            I => \N__16438\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__16438\,
            I => \N__16435\
        );

    \I__2089\ : Span12Mux_s9_v
    port map (
            O => \N__16435\,
            I => \N__16432\
        );

    \I__2088\ : Odrv12
    port map (
            O => \N__16432\,
            I => \M_vcounter_q_esr_RNIQJSA2_0_9\
        );

    \I__2087\ : InMux
    port map (
            O => \N__16429\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__2086\ : InMux
    port map (
            O => \N__16426\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__2085\ : InMux
    port map (
            O => \N__16423\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__2084\ : InMux
    port map (
            O => \N__16420\,
            I => \bfn_5_10_0_\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__16417\,
            I => \this_vga_signals.un4_hsynclto3_0_cascade_\
        );

    \I__2082\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16411\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__16411\,
            I => this_vga_signals_un4_lvisibility_1
        );

    \I__2080\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16404\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__16407\,
            I => \N__16401\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__16404\,
            I => \N__16394\
        );

    \I__2077\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16391\
        );

    \I__2076\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16388\
        );

    \I__2075\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16382\
        );

    \I__2074\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16382\
        );

    \I__2073\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16373\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__16394\,
            I => \N__16368\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__16391\,
            I => \N__16368\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__16388\,
            I => \N__16365\
        );

    \I__2069\ : InMux
    port map (
            O => \N__16387\,
            I => \N__16362\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__16382\,
            I => \N__16359\
        );

    \I__2067\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16356\
        );

    \I__2066\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16351\
        );

    \I__2065\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16351\
        );

    \I__2064\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16346\
        );

    \I__2063\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16346\
        );

    \I__2062\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16343\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__16373\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__16368\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__16365\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__16362\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__16359\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__16356\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__16351\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__16346\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__16343\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__2052\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16321\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__16321\,
            I => \N__16317\
        );

    \I__2050\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16314\
        );

    \I__2049\ : Span4Mux_h
    port map (
            O => \N__16317\,
            I => \N__16308\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__16314\,
            I => \N__16308\
        );

    \I__2047\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16305\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__16308\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__16305\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2044\ : CEMux
    port map (
            O => \N__16300\,
            I => \N__16273\
        );

    \I__2043\ : CEMux
    port map (
            O => \N__16299\,
            I => \N__16273\
        );

    \I__2042\ : CEMux
    port map (
            O => \N__16298\,
            I => \N__16273\
        );

    \I__2041\ : CEMux
    port map (
            O => \N__16297\,
            I => \N__16273\
        );

    \I__2040\ : CEMux
    port map (
            O => \N__16296\,
            I => \N__16273\
        );

    \I__2039\ : CEMux
    port map (
            O => \N__16295\,
            I => \N__16273\
        );

    \I__2038\ : CEMux
    port map (
            O => \N__16294\,
            I => \N__16273\
        );

    \I__2037\ : CEMux
    port map (
            O => \N__16293\,
            I => \N__16273\
        );

    \I__2036\ : CEMux
    port map (
            O => \N__16292\,
            I => \N__16273\
        );

    \I__2035\ : GlobalMux
    port map (
            O => \N__16273\,
            I => \N__16270\
        );

    \I__2034\ : gio2CtrlBuf
    port map (
            O => \N__16270\,
            I => \this_vga_signals.N_935_0_g\
        );

    \I__2033\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16264\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__16264\,
            I => \N__16251\
        );

    \I__2031\ : SRMux
    port map (
            O => \N__16263\,
            I => \N__16228\
        );

    \I__2030\ : SRMux
    port map (
            O => \N__16262\,
            I => \N__16228\
        );

    \I__2029\ : SRMux
    port map (
            O => \N__16261\,
            I => \N__16228\
        );

    \I__2028\ : SRMux
    port map (
            O => \N__16260\,
            I => \N__16228\
        );

    \I__2027\ : SRMux
    port map (
            O => \N__16259\,
            I => \N__16228\
        );

    \I__2026\ : SRMux
    port map (
            O => \N__16258\,
            I => \N__16228\
        );

    \I__2025\ : SRMux
    port map (
            O => \N__16257\,
            I => \N__16228\
        );

    \I__2024\ : SRMux
    port map (
            O => \N__16256\,
            I => \N__16228\
        );

    \I__2023\ : SRMux
    port map (
            O => \N__16255\,
            I => \N__16228\
        );

    \I__2022\ : SRMux
    port map (
            O => \N__16254\,
            I => \N__16228\
        );

    \I__2021\ : Glb2LocalMux
    port map (
            O => \N__16251\,
            I => \N__16228\
        );

    \I__2020\ : GlobalMux
    port map (
            O => \N__16228\,
            I => \N__16225\
        );

    \I__2019\ : gio2CtrlBuf
    port map (
            O => \N__16225\,
            I => \this_vga_signals.N_1212_g\
        );

    \I__2018\ : InMux
    port map (
            O => \N__16222\,
            I => \N__16219\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__16216\,
            I => \this_vga_signals.un4_hsynclto7_0\
        );

    \I__2015\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16207\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__16204\,
            I => \this_vga_signals.un4_hsynclt9\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__16201\,
            I => \this_vga_signals.if_N_8_i_0_cascade_\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__16198\,
            I => \this_vga_signals.if_N_9_0_0_cascade_\
        );

    \I__2009\ : InMux
    port map (
            O => \N__16195\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__2008\ : InMux
    port map (
            O => \N__16192\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__2007\ : InMux
    port map (
            O => \N__16189\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__2006\ : InMux
    port map (
            O => \N__16186\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__16183\,
            I => \this_vga_signals.r_N_4_mux_cascade_\
        );

    \I__2004\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16176\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__16176\,
            I => \this_vga_signals.N_24_0\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__16173\,
            I => \this_vga_signals.N_24_0\
        );

    \I__2000\ : InMux
    port map (
            O => \N__16168\,
            I => \N__16165\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__16165\,
            I => \this_vga_signals.r_N_4_mux\
        );

    \I__1998\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16157\
        );

    \I__1997\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16151\
        );

    \I__1996\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16148\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16145\
        );

    \I__1994\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16140\
        );

    \I__1993\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16140\
        );

    \I__1992\ : InMux
    port map (
            O => \N__16154\,
            I => \N__16137\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__16151\,
            I => \N__16134\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__16148\,
            I => \N__16130\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__16145\,
            I => \N__16123\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__16140\,
            I => \N__16123\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__16137\,
            I => \N__16123\
        );

    \I__1986\ : Span4Mux_v
    port map (
            O => \N__16134\,
            I => \N__16120\
        );

    \I__1985\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16117\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__16130\,
            I => \N__16114\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__16123\,
            I => \N__16111\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__16120\,
            I => \this_vga_signals.N_32_0\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__16117\,
            I => \this_vga_signals.N_32_0\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__16114\,
            I => \this_vga_signals.N_32_0\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__16111\,
            I => \this_vga_signals.N_32_0\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__16102\,
            I => \this_vga_signals.N_24_0_2_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16093\
        );

    \I__1976\ : InMux
    port map (
            O => \N__16098\,
            I => \N__16090\
        );

    \I__1975\ : InMux
    port map (
            O => \N__16097\,
            I => \N__16087\
        );

    \I__1974\ : InMux
    port map (
            O => \N__16096\,
            I => \N__16084\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__16093\,
            I => \this_vga_signals.mult1_un40_sum_c2_0\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__16090\,
            I => \this_vga_signals.mult1_un40_sum_c2_0\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__16087\,
            I => \this_vga_signals.mult1_un40_sum_c2_0\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__16084\,
            I => \this_vga_signals.mult1_un40_sum_c2_0\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16072\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__16072\,
            I => \N__16068\
        );

    \I__1967\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16065\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__16068\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__16065\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__16057\,
            I => \N__16052\
        );

    \I__1962\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16047\
        );

    \I__1961\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16047\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__16052\,
            I => \N__16041\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__16047\,
            I => \N__16041\
        );

    \I__1958\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16038\
        );

    \I__1957\ : Span4Mux_h
    port map (
            O => \N__16041\,
            I => \N__16035\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__16038\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_0_0\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__16035\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_0_0\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__16030\,
            I => \this_vga_signals.g0_23_cascade_\
        );

    \I__1953\ : InMux
    port map (
            O => \N__16027\,
            I => \N__16020\
        );

    \I__1952\ : InMux
    port map (
            O => \N__16026\,
            I => \N__16015\
        );

    \I__1951\ : InMux
    port map (
            O => \N__16025\,
            I => \N__16015\
        );

    \I__1950\ : InMux
    port map (
            O => \N__16024\,
            I => \N__16010\
        );

    \I__1949\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16010\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__16020\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__16015\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__16010\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__16003\,
            I => \N__16000\
        );

    \I__1944\ : InMux
    port map (
            O => \N__16000\,
            I => \N__15997\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__15997\,
            I => \this_vga_signals.g0_1_0_0\
        );

    \I__1942\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15991\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__15991\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__1940\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15985\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__15985\,
            I => \this_vga_signals.g0_0_2_0\
        );

    \I__1938\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15979\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__15979\,
            I => \N__15976\
        );

    \I__1936\ : Odrv12
    port map (
            O => \N__15976\,
            I => \this_vga_signals.un2_hsynclt7\
        );

    \I__1935\ : IoInMux
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__15970\,
            I => \N__15967\
        );

    \I__1933\ : IoSpan4Mux
    port map (
            O => \N__15967\,
            I => \N__15964\
        );

    \I__1932\ : Sp12to4
    port map (
            O => \N__15964\,
            I => \N__15961\
        );

    \I__1931\ : Span12Mux_s6_v
    port map (
            O => \N__15961\,
            I => \N__15958\
        );

    \I__1930\ : Odrv12
    port map (
            O => \N__15958\,
            I => this_vga_signals_hsync_1_i
        );

    \I__1929\ : IoInMux
    port map (
            O => \N__15955\,
            I => \N__15952\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__15952\,
            I => \N__15949\
        );

    \I__1927\ : Span4Mux_s3_h
    port map (
            O => \N__15949\,
            I => \N__15946\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__15946\,
            I => \N__15943\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__15943\,
            I => \N__15940\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__15940\,
            I => rgb_c_5
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__15937\,
            I => \this_vga_signals.r_N_4_mux_1_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__15934\,
            I => \N__15931\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__15931\,
            I => \N__15928\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__15928\,
            I => \this_vga_signals.N_24_0_1\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__15925\,
            I => \this_vga_signals.un2_hsynclt6_0_cascade_\
        );

    \I__1918\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15919\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__15919\,
            I => \N__15914\
        );

    \I__1916\ : InMux
    port map (
            O => \N__15918\,
            I => \N__15911\
        );

    \I__1915\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15908\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__15914\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__15911\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__15908\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__1911\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15898\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__15898\,
            I => \N__15895\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__15895\,
            I => \this_vga_signals.r_N_4_mux_0\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__15892\,
            I => \this_vga_signals.N_24_0_0_cascade_\
        );

    \I__1907\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15883\
        );

    \I__1906\ : InMux
    port map (
            O => \N__15888\,
            I => \N__15883\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__15883\,
            I => \this_vga_signals.N_4_2_0\
        );

    \I__1904\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15877\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__15877\,
            I => \N__15873\
        );

    \I__1902\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15870\
        );

    \I__1901\ : Span4Mux_v
    port map (
            O => \N__15873\,
            I => \N__15864\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__15870\,
            I => \N__15864\
        );

    \I__1899\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15861\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__15864\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__15861\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1896\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15853\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__15853\,
            I => \N__15850\
        );

    \I__1894\ : Span4Mux_s3_h
    port map (
            O => \N__15850\,
            I => \N__15847\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__15847\,
            I => \this_vga_signals.g0_0_i_a5_1_0\
        );

    \I__1892\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15841\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__15841\,
            I => \N__15834\
        );

    \I__1890\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15831\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__15839\,
            I => \N__15828\
        );

    \I__1888\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15825\
        );

    \I__1887\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15818\
        );

    \I__1886\ : Span4Mux_h
    port map (
            O => \N__15834\,
            I => \N__15815\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__15831\,
            I => \N__15812\
        );

    \I__1884\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15809\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__15825\,
            I => \N__15806\
        );

    \I__1882\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15797\
        );

    \I__1881\ : InMux
    port map (
            O => \N__15823\,
            I => \N__15797\
        );

    \I__1880\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15797\
        );

    \I__1879\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15797\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__15818\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__15815\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1876\ : Odrv12
    port map (
            O => \N__15812\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__15809\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__15806\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__15797\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__1872\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15779\
        );

    \I__1871\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15774\
        );

    \I__1870\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15774\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__15779\,
            I => \N__15769\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__15774\,
            I => \N__15766\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__15773\,
            I => \N__15758\
        );

    \I__1866\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15754\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__15769\,
            I => \N__15751\
        );

    \I__1864\ : Span4Mux_h
    port map (
            O => \N__15766\,
            I => \N__15748\
        );

    \I__1863\ : InMux
    port map (
            O => \N__15765\,
            I => \N__15745\
        );

    \I__1862\ : InMux
    port map (
            O => \N__15764\,
            I => \N__15732\
        );

    \I__1861\ : InMux
    port map (
            O => \N__15763\,
            I => \N__15732\
        );

    \I__1860\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15732\
        );

    \I__1859\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15732\
        );

    \I__1858\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15732\
        );

    \I__1857\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15732\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__15754\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__15751\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__15748\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__15745\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__15732\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__1851\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15718\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__15718\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__15715\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_\
        );

    \I__1848\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15709\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__15709\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0_0\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__15706\,
            I => \this_vga_signals.vvisibility_i_o2_1_cascade_\
        );

    \I__1845\ : InMux
    port map (
            O => \N__15703\,
            I => \N__15700\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__15700\,
            I => \N__15696\
        );

    \I__1843\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15693\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__15696\,
            I => \this_vga_signals.vaddress_m2_e_1\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__15693\,
            I => \this_vga_signals.vaddress_m2_e_1\
        );

    \I__1840\ : InMux
    port map (
            O => \N__15688\,
            I => \N__15684\
        );

    \I__1839\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15681\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__15684\,
            I => \N__15674\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__15681\,
            I => \N__15674\
        );

    \I__1836\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15667\
        );

    \I__1835\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15667\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__15674\,
            I => \N__15664\
        );

    \I__1833\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15661\
        );

    \I__1832\ : InMux
    port map (
            O => \N__15672\,
            I => \N__15657\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__15667\,
            I => \N__15654\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__15664\,
            I => \N__15649\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__15661\,
            I => \N__15649\
        );

    \I__1828\ : InMux
    port map (
            O => \N__15660\,
            I => \N__15646\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__15657\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1826\ : Odrv12
    port map (
            O => \N__15654\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__15649\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__15646\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__1823\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15634\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15628\
        );

    \I__1821\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15622\
        );

    \I__1820\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15622\
        );

    \I__1819\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15617\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__15628\,
            I => \N__15614\
        );

    \I__1817\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15611\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15606\
        );

    \I__1815\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15603\
        );

    \I__1814\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15600\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__15617\,
            I => \N__15594\
        );

    \I__1812\ : IoSpan4Mux
    port map (
            O => \N__15614\,
            I => \N__15591\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__15611\,
            I => \N__15588\
        );

    \I__1810\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15583\
        );

    \I__1809\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15583\
        );

    \I__1808\ : Span4Mux_s2_h
    port map (
            O => \N__15606\,
            I => \N__15580\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__15603\,
            I => \N__15577\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__15600\,
            I => \N__15573\
        );

    \I__1805\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15570\
        );

    \I__1804\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15565\
        );

    \I__1803\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15565\
        );

    \I__1802\ : Span4Mux_v
    port map (
            O => \N__15594\,
            I => \N__15558\
        );

    \I__1801\ : Span4Mux_s2_h
    port map (
            O => \N__15591\,
            I => \N__15558\
        );

    \I__1800\ : Span4Mux_s2_h
    port map (
            O => \N__15588\,
            I => \N__15558\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__15583\,
            I => \N__15551\
        );

    \I__1798\ : Span4Mux_h
    port map (
            O => \N__15580\,
            I => \N__15551\
        );

    \I__1797\ : Span4Mux_s2_h
    port map (
            O => \N__15577\,
            I => \N__15551\
        );

    \I__1796\ : InMux
    port map (
            O => \N__15576\,
            I => \N__15547\
        );

    \I__1795\ : Span4Mux_s2_h
    port map (
            O => \N__15573\,
            I => \N__15544\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__15570\,
            I => \N__15541\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__15565\,
            I => \N__15534\
        );

    \I__1792\ : Sp12to4
    port map (
            O => \N__15558\,
            I => \N__15534\
        );

    \I__1791\ : Sp12to4
    port map (
            O => \N__15551\,
            I => \N__15534\
        );

    \I__1790\ : InMux
    port map (
            O => \N__15550\,
            I => \N__15531\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__15547\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__15544\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__15541\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__15534\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__15531\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__15520\,
            I => \N__15509\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__15519\,
            I => \N__15506\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__15518\,
            I => \N__15502\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__15517\,
            I => \N__15499\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \N__15495\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__15515\,
            I => \N__15492\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__15514\,
            I => \N__15487\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__15513\,
            I => \N__15484\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__15512\,
            I => \N__15481\
        );

    \I__1775\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15477\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15506\,
            I => \N__15473\
        );

    \I__1773\ : InMux
    port map (
            O => \N__15505\,
            I => \N__15470\
        );

    \I__1772\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15467\
        );

    \I__1771\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15458\
        );

    \I__1770\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15458\
        );

    \I__1769\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15458\
        );

    \I__1768\ : InMux
    port map (
            O => \N__15492\,
            I => \N__15458\
        );

    \I__1767\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15455\
        );

    \I__1766\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15452\
        );

    \I__1765\ : InMux
    port map (
            O => \N__15487\,
            I => \N__15449\
        );

    \I__1764\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15444\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15444\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15441\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15477\,
            I => \N__15438\
        );

    \I__1760\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15435\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__15473\,
            I => \N__15430\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__15470\,
            I => \N__15430\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__15467\,
            I => \N__15425\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__15458\,
            I => \N__15425\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__15455\,
            I => \N__15417\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__15452\,
            I => \N__15417\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__15449\,
            I => \N__15412\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__15444\,
            I => \N__15412\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__15441\,
            I => \N__15401\
        );

    \I__1750\ : Span4Mux_s1_h
    port map (
            O => \N__15438\,
            I => \N__15401\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__15435\,
            I => \N__15401\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__15430\,
            I => \N__15401\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__15425\,
            I => \N__15401\
        );

    \I__1746\ : InMux
    port map (
            O => \N__15424\,
            I => \N__15396\
        );

    \I__1745\ : InMux
    port map (
            O => \N__15423\,
            I => \N__15393\
        );

    \I__1744\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15390\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__15417\,
            I => \N__15387\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__15412\,
            I => \N__15384\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__15401\,
            I => \N__15381\
        );

    \I__1740\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15377\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__15399\,
            I => \N__15374\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__15396\,
            I => \N__15369\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__15393\,
            I => \N__15369\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__15390\,
            I => \N__15360\
        );

    \I__1735\ : Span4Mux_s1_h
    port map (
            O => \N__15387\,
            I => \N__15360\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__15384\,
            I => \N__15360\
        );

    \I__1733\ : Span4Mux_s1_h
    port map (
            O => \N__15381\,
            I => \N__15360\
        );

    \I__1732\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15357\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__15377\,
            I => \N__15354\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15351\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__15369\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__15360\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__15357\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__15354\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__15351\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__1724\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15336\
        );

    \I__1723\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15332\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__15336\,
            I => \N__15329\
        );

    \I__1721\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15326\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__15332\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1719\ : Odrv12
    port map (
            O => \N__15329\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__15326\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__15319\,
            I => \this_vga_signals.N_822_0_cascade_\
        );

    \I__1716\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15308\
        );

    \I__1715\ : InMux
    port map (
            O => \N__15315\,
            I => \N__15308\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__15314\,
            I => \N__15302\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__15313\,
            I => \N__15299\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__15308\,
            I => \N__15296\
        );

    \I__1711\ : InMux
    port map (
            O => \N__15307\,
            I => \N__15293\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15290\
        );

    \I__1709\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15285\
        );

    \I__1708\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15285\
        );

    \I__1707\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15282\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__15296\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__15293\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__15290\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__15285\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__15282\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__1701\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15265\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__15270\,
            I => \N__15257\
        );

    \I__1699\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15248\
        );

    \I__1698\ : InMux
    port map (
            O => \N__15268\,
            I => \N__15248\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__15265\,
            I => \N__15245\
        );

    \I__1696\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15242\
        );

    \I__1695\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15235\
        );

    \I__1694\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15235\
        );

    \I__1693\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15235\
        );

    \I__1692\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15232\
        );

    \I__1691\ : InMux
    port map (
            O => \N__15257\,
            I => \N__15225\
        );

    \I__1690\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15225\
        );

    \I__1689\ : InMux
    port map (
            O => \N__15255\,
            I => \N__15225\
        );

    \I__1688\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15220\
        );

    \I__1687\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15220\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__15248\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__15245\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__15242\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__15235\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__15232\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__15225\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__15220\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__1679\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15202\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__15202\,
            I => \N__15195\
        );

    \I__1677\ : InMux
    port map (
            O => \N__15201\,
            I => \N__15192\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__15200\,
            I => \N__15189\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__15199\,
            I => \N__15186\
        );

    \I__1674\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15180\
        );

    \I__1673\ : Span4Mux_s3_h
    port map (
            O => \N__15195\,
            I => \N__15177\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__15192\,
            I => \N__15174\
        );

    \I__1671\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15171\
        );

    \I__1670\ : InMux
    port map (
            O => \N__15186\,
            I => \N__15168\
        );

    \I__1669\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15165\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15162\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15159\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__15180\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__15177\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__15174\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__15171\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__15168\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__15165\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__15162\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__15159\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__1658\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15133\
        );

    \I__1657\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15128\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15128\
        );

    \I__1655\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15125\
        );

    \I__1654\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15118\
        );

    \I__1653\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15118\
        );

    \I__1652\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15118\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__15133\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__15128\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__15125\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__15118\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__15109\,
            I => \N__15106\
        );

    \I__1646\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15103\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15100\
        );

    \I__1644\ : Span4Mux_s3_h
    port map (
            O => \N__15100\,
            I => \N__15097\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__15097\,
            I => \this_vga_signals.mult1_un40_sum_ac0_0_0\
        );

    \I__1642\ : IoInMux
    port map (
            O => \N__15094\,
            I => \N__15091\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__15091\,
            I => \N__15088\
        );

    \I__1640\ : Span4Mux_s2_h
    port map (
            O => \N__15088\,
            I => \N__15085\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__15085\,
            I => rgb_c_2
        );

    \I__1638\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15079\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__15079\,
            I => \N__15076\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__15076\,
            I => \this_vga_signals.vsync_1_0_a2_3\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__15073\,
            I => \N__15070\
        );

    \I__1634\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15067\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__15067\,
            I => \this_vga_signals.vsync_1_0_a2_4\
        );

    \I__1632\ : IoInMux
    port map (
            O => \N__15064\,
            I => \N__15061\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__15061\,
            I => \N__15058\
        );

    \I__1630\ : Span12Mux_s11_v
    port map (
            O => \N__15058\,
            I => \N__15055\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__15055\,
            I => this_vga_signals_vsync_1_i
        );

    \I__1628\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15049\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__15049\,
            I => \N__15046\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__15046\,
            I => \this_vga_signals.if_N_6_0\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__15043\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__15040\,
            I => \N__15037\
        );

    \I__1623\ : InMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__15034\,
            I => \this_vga_signals.mult1_un75_sum_axb2_0\
        );

    \I__1621\ : IoInMux
    port map (
            O => \N__15031\,
            I => \N__15028\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__15028\,
            I => \N__15025\
        );

    \I__1619\ : Span4Mux_s2_h
    port map (
            O => \N__15025\,
            I => \N__15022\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__15022\,
            I => \N__15019\
        );

    \I__1617\ : Span4Mux_v
    port map (
            O => \N__15019\,
            I => \N__15016\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__15016\,
            I => rgb_c_3
        );

    \I__1615\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15009\
        );

    \I__1614\ : InMux
    port map (
            O => \N__15012\,
            I => \N__15003\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__15009\,
            I => \N__15000\
        );

    \I__1612\ : InMux
    port map (
            O => \N__15008\,
            I => \N__14995\
        );

    \I__1611\ : InMux
    port map (
            O => \N__15007\,
            I => \N__14995\
        );

    \I__1610\ : InMux
    port map (
            O => \N__15006\,
            I => \N__14992\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__15003\,
            I => \N__14989\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__15000\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_1\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__14995\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_1\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__14992\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_1\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__14989\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1_1\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__14980\,
            I => \N__14975\
        );

    \I__1603\ : InMux
    port map (
            O => \N__14979\,
            I => \N__14970\
        );

    \I__1602\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14966\
        );

    \I__1601\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14963\
        );

    \I__1600\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14955\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__14973\,
            I => \N__14947\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__14970\,
            I => \N__14944\
        );

    \I__1597\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14941\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__14966\,
            I => \N__14938\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__14963\,
            I => \N__14935\
        );

    \I__1594\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14930\
        );

    \I__1593\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14930\
        );

    \I__1592\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14927\
        );

    \I__1591\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14922\
        );

    \I__1590\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14922\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__14955\,
            I => \N__14919\
        );

    \I__1588\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14916\
        );

    \I__1587\ : InMux
    port map (
            O => \N__14953\,
            I => \N__14911\
        );

    \I__1586\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14911\
        );

    \I__1585\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14904\
        );

    \I__1584\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14904\
        );

    \I__1583\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14904\
        );

    \I__1582\ : Span4Mux_v
    port map (
            O => \N__14944\,
            I => \N__14891\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__14941\,
            I => \N__14891\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__14938\,
            I => \N__14891\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__14935\,
            I => \N__14891\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__14930\,
            I => \N__14891\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14891\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14922\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__14919\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__14916\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__14911\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__14904\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__14891\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__1570\ : InMux
    port map (
            O => \N__14878\,
            I => \N__14875\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__14875\,
            I => \this_vga_signals.g3_0_1\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__14872\,
            I => \N__14869\
        );

    \I__1567\ : InMux
    port map (
            O => \N__14869\,
            I => \N__14866\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__14866\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_c_0\
        );

    \I__1565\ : InMux
    port map (
            O => \N__14863\,
            I => \N__14860\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__14860\,
            I => \N__14857\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__14857\,
            I => \this_vga_signals.mult1_un75_sum_ac0_3_d\
        );

    \I__1562\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14851\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__14851\,
            I => \this_vga_signals.M_vcounter_q_RNI0FQEQVZ0Z_2\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__14848\,
            I => \this_vga_signals.mult1_un75_sum_c3_0_0_0_cascade_\
        );

    \I__1559\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14842\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__14842\,
            I => \this_vga_signals.vaddress_m6_0\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__14839\,
            I => \N__14836\
        );

    \I__1556\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14833\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__14833\,
            I => \N__14830\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__14830\,
            I => \N__14827\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__14827\,
            I => \N__14824\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__14824\,
            I => \N__14821\
        );

    \I__1551\ : Span4Mux_v
    port map (
            O => \N__14821\,
            I => \N__14818\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__14818\,
            I => \M_this_vga_signals_address_7\
        );

    \I__1549\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14809\
        );

    \I__1548\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14806\
        );

    \I__1547\ : InMux
    port map (
            O => \N__14813\,
            I => \N__14803\
        );

    \I__1546\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14800\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__14809\,
            I => \this_vga_signals.mult1_un61_sum_ac0_4\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__14806\,
            I => \this_vga_signals.mult1_un61_sum_ac0_4\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__14803\,
            I => \this_vga_signals.mult1_un61_sum_ac0_4\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__14800\,
            I => \this_vga_signals.mult1_un61_sum_ac0_4\
        );

    \I__1541\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14788\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__14788\,
            I => \N__14785\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__14785\,
            I => \this_vga_signals.g0_0\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__14782\,
            I => \N__14779\
        );

    \I__1537\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14776\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__14776\,
            I => \this_vga_signals.g0_0_0_0\
        );

    \I__1535\ : InMux
    port map (
            O => \N__14773\,
            I => \N__14770\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__14770\,
            I => \this_vga_signals.g3\
        );

    \I__1533\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14764\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__14764\,
            I => \N__14761\
        );

    \I__1531\ : Odrv12
    port map (
            O => \N__14761\,
            I => \this_vga_signals.g0_0_0_a2_2_0\
        );

    \I__1530\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14755\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__14755\,
            I => \this_vga_signals.g0_6_0_a2_3\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__14752\,
            I => \this_vga_signals.N_12_0_0_cascade_\
        );

    \I__1527\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14745\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__14748\,
            I => \N__14741\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__14745\,
            I => \N__14735\
        );

    \I__1524\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14732\
        );

    \I__1523\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14729\
        );

    \I__1522\ : InMux
    port map (
            O => \N__14740\,
            I => \N__14722\
        );

    \I__1521\ : InMux
    port map (
            O => \N__14739\,
            I => \N__14722\
        );

    \I__1520\ : InMux
    port map (
            O => \N__14738\,
            I => \N__14722\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__14735\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__14732\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__14729\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__14722\,
            I => \this_vga_signals.mult1_un68_sum_c3\
        );

    \I__1515\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14710\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__14710\,
            I => \this_vga_signals.g0_1_1\
        );

    \I__1513\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14700\
        );

    \I__1512\ : InMux
    port map (
            O => \N__14706\,
            I => \N__14700\
        );

    \I__1511\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14697\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__14700\,
            I => \N__14687\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__14697\,
            I => \N__14684\
        );

    \I__1508\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14681\
        );

    \I__1507\ : InMux
    port map (
            O => \N__14695\,
            I => \N__14678\
        );

    \I__1506\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14675\
        );

    \I__1505\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14672\
        );

    \I__1504\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14667\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14667\
        );

    \I__1502\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14664\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__14687\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1500\ : Odrv4
    port map (
            O => \N__14684\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__14681\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__14678\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__14675\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__14672\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__14667\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__14664\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__1493\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14644\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__14644\,
            I => \this_vga_signals.g0_0_i_a5_1\
        );

    \I__1491\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14638\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__14638\,
            I => \N__14635\
        );

    \I__1489\ : Span4Mux_v
    port map (
            O => \N__14635\,
            I => \N__14632\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__14632\,
            I => \this_vga_signals.N_8\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__14629\,
            I => \this_vga_signals.N_6_0_cascade_\
        );

    \I__1486\ : InMux
    port map (
            O => \N__14626\,
            I => \N__14623\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__14623\,
            I => \this_vga_signals.g0_1\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14617\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__14617\,
            I => \this_vga_signals.g3_0_0\
        );

    \I__1482\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14611\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__14611\,
            I => \this_vga_signals.g3_1_0\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__14608\,
            I => \N__14605\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14605\,
            I => \N__14602\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__14602\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_0\
        );

    \I__1477\ : InMux
    port map (
            O => \N__14599\,
            I => \N__14596\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__14596\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_0_2\
        );

    \I__1475\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14587\
        );

    \I__1474\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14584\
        );

    \I__1473\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14577\
        );

    \I__1472\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14577\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14574\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__14584\,
            I => \N__14571\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14562\
        );

    \I__1468\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14559\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__14577\,
            I => \N__14552\
        );

    \I__1466\ : Span4Mux_v
    port map (
            O => \N__14574\,
            I => \N__14552\
        );

    \I__1465\ : Span4Mux_s2_h
    port map (
            O => \N__14571\,
            I => \N__14552\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14549\
        );

    \I__1463\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14544\
        );

    \I__1462\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14544\
        );

    \I__1461\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14537\
        );

    \I__1460\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14537\
        );

    \I__1459\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14537\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__14562\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__14559\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__14552\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__14549\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__14544\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__14537\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__1452\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__14521\,
            I => \N__14518\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__14518\,
            I => \this_vga_signals.g0_15\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__14515\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1_cascade_\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__14512\,
            I => \this_vga_signals.N_1_4_1_cascade_\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__14509\,
            I => \this_vga_signals.mult1_un40_sum_c2_1_cascade_\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__14506\,
            I => \this_vga_signals.mult1_un40_sum_c2_0_cascade_\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__14503\,
            I => \this_vga_signals.mult1_un40_sum_c2_2_1_0_cascade_\
        );

    \I__1444\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14497\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__14497\,
            I => \this_vga_signals.mult1_un40_sum_c2_2\
        );

    \I__1442\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14491\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__14491\,
            I => \N__14488\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__14488\,
            I => \this_vga_signals.N_4_3\
        );

    \I__1439\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14482\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__14482\,
            I => \this_vga_signals.g1_1_1\
        );

    \I__1437\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14476\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__14476\,
            I => \this_vga_signals.mult1_un40_sum_ac0_2\
        );

    \I__1435\ : InMux
    port map (
            O => \N__14473\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__14470\,
            I => \N__14467\
        );

    \I__1433\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14464\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__14464\,
            I => \N__14461\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__14461\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2_2_N_2L1\
        );

    \I__1430\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14455\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__14455\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2_2\
        );

    \I__1428\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14447\
        );

    \I__1427\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14444\
        );

    \I__1426\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14441\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__14447\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__14444\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__14441\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__1422\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14431\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__14431\,
            I => \N__14427\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14424\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__14427\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__14424\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__1417\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14416\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__14416\,
            I => \N__14410\
        );

    \I__1415\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14405\
        );

    \I__1414\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14405\
        );

    \I__1413\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14402\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__14410\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__14405\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__14402\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14395\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__1408\ : InMux
    port map (
            O => \N__14392\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__1407\ : InMux
    port map (
            O => \N__14389\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__1406\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14383\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__14383\,
            I => \N__14379\
        );

    \I__1404\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14376\
        );

    \I__1403\ : Span4Mux_s2_h
    port map (
            O => \N__14379\,
            I => \N__14372\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__14376\,
            I => \N__14369\
        );

    \I__1401\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14366\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__14372\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__14369\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__14366\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1397\ : InMux
    port map (
            O => \N__14359\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__1396\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14350\
        );

    \I__1395\ : InMux
    port map (
            O => \N__14355\,
            I => \N__14350\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__14350\,
            I => \N__14347\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__14347\,
            I => \N__14343\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14340\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__14343\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14340\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1389\ : InMux
    port map (
            O => \N__14335\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__1388\ : InMux
    port map (
            O => \N__14332\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__1387\ : InMux
    port map (
            O => \N__14329\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__1386\ : InMux
    port map (
            O => \N__14326\,
            I => \bfn_3_10_0_\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__14323\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_cascade_\
        );

    \I__1384\ : InMux
    port map (
            O => \N__14320\,
            I => \N__14317\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__14317\,
            I => \this_vga_signals.g0_2\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__14314\,
            I => \this_vga_signals.mult1_un68_sum_0_3_cascade_\
        );

    \I__1381\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14308\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__14308\,
            I => \this_vga_signals.mult1_un75_sum_ac0_1\
        );

    \I__1379\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14294\
        );

    \I__1378\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14294\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14294\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__14302\,
            I => \N__14289\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__14301\,
            I => \N__14286\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__14294\,
            I => \N__14278\
        );

    \I__1373\ : InMux
    port map (
            O => \N__14293\,
            I => \N__14273\
        );

    \I__1372\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14273\
        );

    \I__1371\ : InMux
    port map (
            O => \N__14289\,
            I => \N__14270\
        );

    \I__1370\ : InMux
    port map (
            O => \N__14286\,
            I => \N__14267\
        );

    \I__1369\ : InMux
    port map (
            O => \N__14285\,
            I => \N__14259\
        );

    \I__1368\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14259\
        );

    \I__1367\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14252\
        );

    \I__1366\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14252\
        );

    \I__1365\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14252\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__14278\,
            I => \N__14243\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__14273\,
            I => \N__14243\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__14270\,
            I => \N__14243\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__14267\,
            I => \N__14243\
        );

    \I__1360\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14236\
        );

    \I__1359\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14236\
        );

    \I__1358\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14236\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__14259\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__14252\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__14243\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__14236\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1353\ : InMux
    port map (
            O => \N__14227\,
            I => \N__14224\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14220\
        );

    \I__1351\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14214\
        );

    \I__1350\ : Span4Mux_h
    port map (
            O => \N__14220\,
            I => \N__14211\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14204\
        );

    \I__1348\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14204\
        );

    \I__1347\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14204\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__14214\,
            I => \N__14201\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__14211\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__14204\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__14201\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__14194\,
            I => \this_vga_signals.g3_0_a2_2_cascade_\
        );

    \I__1341\ : InMux
    port map (
            O => \N__14191\,
            I => \N__14184\
        );

    \I__1340\ : InMux
    port map (
            O => \N__14190\,
            I => \N__14184\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14189\,
            I => \N__14181\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__14184\,
            I => \this_vga_signals.mult1_un75_sum_axb2\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__14181\,
            I => \this_vga_signals.mult1_un75_sum_axb2\
        );

    \I__1336\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14173\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__14173\,
            I => \this_vga_signals.g0_1_0\
        );

    \I__1334\ : InMux
    port map (
            O => \N__14170\,
            I => \N__14166\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14169\,
            I => \N__14163\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__14166\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__14163\,
            I => \this_vga_signals.mult1_un61_sum_c3_0\
        );

    \I__1330\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__14155\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0\
        );

    \I__1328\ : InMux
    port map (
            O => \N__14152\,
            I => \N__14149\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__14149\,
            I => \this_vga_signals.if_i4_mux_0\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__14146\,
            I => \this_vga_signals.vaddress_N_3_i_0_0_cascade_\
        );

    \I__1325\ : InMux
    port map (
            O => \N__14143\,
            I => \N__14140\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__14140\,
            I => \N__14137\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__14137\,
            I => \this_vga_signals.g2_4_0\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__14134\,
            I => \N__14131\
        );

    \I__1321\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14128\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__14128\,
            I => \this_vga_signals.g2_0_0\
        );

    \I__1319\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14122\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__14122\,
            I => \this_vga_signals.g0_4_0\
        );

    \I__1317\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14115\
        );

    \I__1316\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14112\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__14115\,
            I => \N__14109\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__14112\,
            I => \N__14106\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__14109\,
            I => \N__14103\
        );

    \I__1312\ : Odrv12
    port map (
            O => \N__14106\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__14103\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0\
        );

    \I__1310\ : InMux
    port map (
            O => \N__14098\,
            I => \N__14095\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__14095\,
            I => \N__14092\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__14092\,
            I => \this_vga_signals.g0_0_6\
        );

    \I__1307\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14086\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__14086\,
            I => \this_vga_signals.g1_0_0_0_0\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__14083\,
            I => \N__14079\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__14082\,
            I => \N__14076\
        );

    \I__1303\ : InMux
    port map (
            O => \N__14079\,
            I => \N__14072\
        );

    \I__1302\ : InMux
    port map (
            O => \N__14076\,
            I => \N__14069\
        );

    \I__1301\ : InMux
    port map (
            O => \N__14075\,
            I => \N__14066\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__14072\,
            I => \N__14056\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__14069\,
            I => \N__14056\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__14066\,
            I => \N__14053\
        );

    \I__1297\ : InMux
    port map (
            O => \N__14065\,
            I => \N__14046\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14046\
        );

    \I__1295\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14046\
        );

    \I__1294\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14041\
        );

    \I__1293\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14041\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__14056\,
            I => \this_vga_signals.mult1_un54_sum_ac0_4\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__14053\,
            I => \this_vga_signals.mult1_un54_sum_ac0_4\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__14046\,
            I => \this_vga_signals.mult1_un54_sum_ac0_4\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__14041\,
            I => \this_vga_signals.mult1_un54_sum_ac0_4\
        );

    \I__1288\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14029\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__14029\,
            I => \N__14026\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__14026\,
            I => \N__14023\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__14023\,
            I => \this_vga_signals.g3_0\
        );

    \I__1284\ : InMux
    port map (
            O => \N__14020\,
            I => \N__14017\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__14017\,
            I => \this_vga_signals.N_3_2\
        );

    \I__1282\ : InMux
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__1281\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14005\
        );

    \I__1280\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14000\
        );

    \I__1279\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14000\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__14008\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__14005\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__14000\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__1274\ : InMux
    port map (
            O => \N__13992\,
            I => \N__13977\
        );

    \I__1273\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13977\
        );

    \I__1272\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13977\
        );

    \I__1271\ : InMux
    port map (
            O => \N__13987\,
            I => \N__13964\
        );

    \I__1270\ : InMux
    port map (
            O => \N__13986\,
            I => \N__13961\
        );

    \I__1269\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13956\
        );

    \I__1268\ : InMux
    port map (
            O => \N__13984\,
            I => \N__13956\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__13977\,
            I => \N__13953\
        );

    \I__1266\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13944\
        );

    \I__1265\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13944\
        );

    \I__1264\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13944\
        );

    \I__1263\ : InMux
    port map (
            O => \N__13973\,
            I => \N__13944\
        );

    \I__1262\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13935\
        );

    \I__1261\ : InMux
    port map (
            O => \N__13971\,
            I => \N__13935\
        );

    \I__1260\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13935\
        );

    \I__1259\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13935\
        );

    \I__1258\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13930\
        );

    \I__1257\ : InMux
    port map (
            O => \N__13967\,
            I => \N__13930\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__13964\,
            I => \N__13927\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__13961\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__13956\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__13953\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__13944\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__13935\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__13930\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1249\ : Odrv12
    port map (
            O => \N__13927\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1248\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13909\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__13909\,
            I => \this_vga_signals.g2_0_0_0\
        );

    \I__1246\ : InMux
    port map (
            O => \N__13906\,
            I => \N__13903\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__13903\,
            I => \this_vga_signals.g3_x0\
        );

    \I__1244\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13893\
        );

    \I__1243\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13893\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__13898\,
            I => \N__13888\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__13893\,
            I => \N__13882\
        );

    \I__1240\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13877\
        );

    \I__1239\ : InMux
    port map (
            O => \N__13891\,
            I => \N__13877\
        );

    \I__1238\ : InMux
    port map (
            O => \N__13888\,
            I => \N__13868\
        );

    \I__1237\ : InMux
    port map (
            O => \N__13887\,
            I => \N__13868\
        );

    \I__1236\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13868\
        );

    \I__1235\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13868\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__13882\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__13877\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__13868\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1231\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13858\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__13858\,
            I => \this_vga_signals.g3_x1\
        );

    \I__1229\ : InMux
    port map (
            O => \N__13855\,
            I => \N__13846\
        );

    \I__1228\ : InMux
    port map (
            O => \N__13854\,
            I => \N__13846\
        );

    \I__1227\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13843\
        );

    \I__1226\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13840\
        );

    \I__1225\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13837\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__13846\,
            I => \N__13834\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__13843\,
            I => \N__13831\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__13840\,
            I => \this_vga_signals.mult1_un61_sum_axb2_i\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__13837\,
            I => \this_vga_signals.mult1_un61_sum_axb2_i\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__13834\,
            I => \this_vga_signals.mult1_un61_sum_axb2_i\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__13831\,
            I => \this_vga_signals.mult1_un61_sum_axb2_i\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__13822\,
            I => \N__13819\
        );

    \I__1217\ : InMux
    port map (
            O => \N__13819\,
            I => \N__13816\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__13816\,
            I => \this_vga_signals.mult1_un61_sum_ac0_1\
        );

    \I__1215\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13810\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__13810\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_3\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__13807\,
            I => \this_vga_signals.g1_0_0_2_cascade_\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__13804\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13798\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__13798\,
            I => \this_vga_signals.g0_0_0_1_0\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__13795\,
            I => \N__13788\
        );

    \I__1208\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13783\
        );

    \I__1207\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13783\
        );

    \I__1206\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13780\
        );

    \I__1205\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13777\
        );

    \I__1204\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13774\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__13783\,
            I => \N__13771\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__13780\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__13777\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__13774\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__13771\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__1198\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13759\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__13759\,
            I => \N__13756\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__13756\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__13753\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13741\
        );

    \I__1193\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13741\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__13748\,
            I => \N__13738\
        );

    \I__1191\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13735\
        );

    \I__1190\ : InMux
    port map (
            O => \N__13746\,
            I => \N__13732\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__13741\,
            I => \N__13729\
        );

    \I__1188\ : InMux
    port map (
            O => \N__13738\,
            I => \N__13726\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__13735\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__13732\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__13729\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__13726\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__13717\,
            I => \N__13712\
        );

    \I__1182\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13698\
        );

    \I__1181\ : InMux
    port map (
            O => \N__13715\,
            I => \N__13698\
        );

    \I__1180\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13693\
        );

    \I__1179\ : InMux
    port map (
            O => \N__13711\,
            I => \N__13693\
        );

    \I__1178\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13688\
        );

    \I__1177\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13688\
        );

    \I__1176\ : InMux
    port map (
            O => \N__13708\,
            I => \N__13679\
        );

    \I__1175\ : InMux
    port map (
            O => \N__13707\,
            I => \N__13679\
        );

    \I__1174\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13679\
        );

    \I__1173\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13679\
        );

    \I__1172\ : InMux
    port map (
            O => \N__13704\,
            I => \N__13674\
        );

    \I__1171\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13674\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__13698\,
            I => \N__13669\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__13693\,
            I => \N__13669\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__13688\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__13679\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__13674\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__13669\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__13660\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_4_cascade_\
        );

    \I__1163\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13654\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__13654\,
            I => \N__13650\
        );

    \I__1161\ : InMux
    port map (
            O => \N__13653\,
            I => \N__13647\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__13650\,
            I => \N__13644\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__13647\,
            I => \this_vga_signals.g2_1_0\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__13644\,
            I => \this_vga_signals.g2_1_0\
        );

    \I__1157\ : InMux
    port map (
            O => \N__13639\,
            I => \N__13636\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__13636\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2_mb_sn\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__13633\,
            I => \N__13629\
        );

    \I__1154\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13625\
        );

    \I__1153\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13620\
        );

    \I__1152\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13620\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__13625\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1_0\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__13620\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1_0\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__13615\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_\
        );

    \I__1148\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13609\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__13609\,
            I => \N__13606\
        );

    \I__1146\ : Span4Mux_v
    port map (
            O => \N__13606\,
            I => \N__13603\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__13603\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_1\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__13600\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x1_cascade_\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__13597\,
            I => \N__13593\
        );

    \I__1142\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13590\
        );

    \I__1141\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13587\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13584\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__13587\,
            I => \this_vga_signals.SUM_2_i_i_1_1_3\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__13584\,
            I => \this_vga_signals.SUM_2_i_i_1_1_3\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__13579\,
            I => \N__13576\
        );

    \I__1136\ : InMux
    port map (
            O => \N__13576\,
            I => \N__13573\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__13573\,
            I => \this_vga_signals.mult1_un40_sum_axb1_x0\
        );

    \I__1134\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13567\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__13567\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x0\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__13564\,
            I => \N__13560\
        );

    \I__1131\ : InMux
    port map (
            O => \N__13563\,
            I => \N__13557\
        );

    \I__1130\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13554\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__13557\,
            I => \this_vga_signals.SUM_2_i_i_1_0_3\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__13554\,
            I => \this_vga_signals.SUM_2_i_i_1_0_3\
        );

    \I__1127\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13546\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__13546\,
            I => \this_vga_signals.mult1_un40_sum_axb1_x1\
        );

    \I__1125\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13538\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__13542\,
            I => \N__13535\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__13541\,
            I => \N__13531\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__13538\,
            I => \N__13528\
        );

    \I__1121\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13525\
        );

    \I__1120\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13520\
        );

    \I__1119\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13520\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__13528\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__13525\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__13520\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__13513\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_x1_cascade_\
        );

    \I__1114\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13507\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__13507\,
            I => \N__13501\
        );

    \I__1112\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13498\
        );

    \I__1111\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13493\
        );

    \I__1110\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13493\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__13501\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__13498\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__13493\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__1106\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13483\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__13483\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_ns\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__13480\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_ns_cascade_\
        );

    \I__1103\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13474\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__13474\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__13471\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__13468\,
            I => \N__13464\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__13467\,
            I => \N__13461\
        );

    \I__1098\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13458\
        );

    \I__1097\ : InMux
    port map (
            O => \N__13461\,
            I => \N__13455\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__13458\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__13455\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__13450\,
            I => \this_vga_signals.SUM_2_i_i_1_0_3_cascade_\
        );

    \I__1093\ : InMux
    port map (
            O => \N__13447\,
            I => \N__13442\
        );

    \I__1092\ : InMux
    port map (
            O => \N__13446\,
            I => \N__13437\
        );

    \I__1091\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13437\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__13442\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__13437\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__13432\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2_x1_cascade_\
        );

    \I__1087\ : InMux
    port map (
            O => \N__13429\,
            I => \N__13426\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__13426\,
            I => \this_vga_signals.g1_0_0_1\
        );

    \I__1085\ : IoInMux
    port map (
            O => \N__13423\,
            I => \N__13420\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__13420\,
            I => \N__13417\
        );

    \I__1083\ : Span4Mux_s2_h
    port map (
            O => \N__13417\,
            I => \N__13414\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__13414\,
            I => \N__13411\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__13411\,
            I => port_data_rw_0_i
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__13408\,
            I => \N__13405\
        );

    \I__1079\ : InMux
    port map (
            O => \N__13405\,
            I => \N__13402\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__13402\,
            I => \this_vga_signals.g2_2_0\
        );

    \I__1077\ : IoInMux
    port map (
            O => \N__13399\,
            I => \N__13396\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__13396\,
            I => \N__13393\
        );

    \I__1075\ : Span4Mux_s2_h
    port map (
            O => \N__13393\,
            I => \N__13390\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__13390\,
            I => rgb_c_0
        );

    \I__1073\ : IoInMux
    port map (
            O => \N__13387\,
            I => \N__13384\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__13384\,
            I => \N__13381\
        );

    \I__1071\ : Span4Mux_s1_h
    port map (
            O => \N__13381\,
            I => \N__13378\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__13378\,
            I => \N__13375\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__13375\,
            I => \N__13372\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__13372\,
            I => rgb_c_1
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__13369\,
            I => \N__13366\
        );

    \I__1066\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13363\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__13363\,
            I => \N__13360\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__13360\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_2\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__13357\,
            I => \N__13354\
        );

    \I__1062\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13351\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__13351\,
            I => \N__13348\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__13348\,
            I => \this_vga_signals.g1_1_0\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__13345\,
            I => \this_vga_signals.g1_4_cascade_\
        );

    \I__1058\ : IoInMux
    port map (
            O => \N__13342\,
            I => \N__13339\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__13339\,
            I => \N__13336\
        );

    \I__1056\ : Span12Mux_s0_h
    port map (
            O => \N__13336\,
            I => \N__13333\
        );

    \I__1055\ : Span12Mux_v
    port map (
            O => \N__13333\,
            I => \N__13330\
        );

    \I__1054\ : Odrv12
    port map (
            O => \N__13330\,
            I => rgb_c_4
        );

    \I__1053\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13322\
        );

    \I__1052\ : InMux
    port map (
            O => \N__13326\,
            I => \N__13317\
        );

    \I__1051\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13317\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__13322\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__13317\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_1\
        );

    \I__1048\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13309\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13306\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__13306\,
            I => \this_vga_signals.vaddress_m2_2\
        );

    \I__1045\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13300\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__13300\,
            I => \N__13297\
        );

    \I__1043\ : IoSpan4Mux
    port map (
            O => \N__13297\,
            I => \N__13294\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__13294\,
            I => port_clk_c
        );

    \I__1041\ : InMux
    port map (
            O => \N__13291\,
            I => \N__13288\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__13288\,
            I => \N__13285\
        );

    \I__1039\ : Odrv12
    port map (
            O => \N__13285\,
            I => \this_vga_signals.g2\
        );

    \I__1038\ : InMux
    port map (
            O => \N__13282\,
            I => \N__13279\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__13279\,
            I => \N__13275\
        );

    \I__1036\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13272\
        );

    \I__1035\ : Span4Mux_v
    port map (
            O => \N__13275\,
            I => \N__13267\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__13272\,
            I => \N__13267\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__13267\,
            I => \this_vga_signals.g1\
        );

    \I__1032\ : IoInMux
    port map (
            O => \N__13264\,
            I => \N__13261\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__13261\,
            I => \this_vga_signals.N_935_0\
        );

    \I__1030\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13255\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__13255\,
            I => \N__13252\
        );

    \I__1028\ : Odrv12
    port map (
            O => \N__13252\,
            I => \this_vga_signals.g3_2\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__13249\,
            I => \this_vga_signals.mult1_un75_sum_axb1_3_cascade_\
        );

    \I__1026\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13243\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N__13240\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__13240\,
            I => \N__13237\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__13237\,
            I => \this_vga_signals.vaddress_m2_1\
        );

    \I__1022\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__13228\,
            I => \this_vga_signals.if_N_9_i\
        );

    \I__1019\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13222\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__13222\,
            I => \this_vga_signals.if_m1_0\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__13219\,
            I => \this_vga_signals.mult1_un68_sum_c3_cascade_\
        );

    \I__1016\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13213\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__13213\,
            I => \N__13210\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__13210\,
            I => \this_vga_signals.mult1_un61_sum_axb2_i_0\
        );

    \I__1013\ : InMux
    port map (
            O => \N__13207\,
            I => \N__13204\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__13204\,
            I => \this_vga_signals.g2_3\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__13201\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0_0_0_cascade_\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__13198\,
            I => \this_vga_signals.mult1_un75_sum_axb1_3_1_1_cascade_\
        );

    \I__1009\ : InMux
    port map (
            O => \N__13195\,
            I => \N__13191\
        );

    \I__1008\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13188\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__13191\,
            I => \this_vga_signals.mult1_un75_sum_axb1_3_1\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__13188\,
            I => \this_vga_signals.mult1_un75_sum_axb1_3_1\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__13183\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_cascade_\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__13180\,
            I => \this_vga_signals.g1_0_0_0_cascade_\
        );

    \I__1003\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13174\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__13174\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__1001\ : InMux
    port map (
            O => \N__13171\,
            I => \N__13168\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__13168\,
            I => \N__13165\
        );

    \I__999\ : Odrv12
    port map (
            O => \N__13165\,
            I => \this_vga_signals.g2_1\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__13162\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_cascade_\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__13159\,
            I => \this_vga_signals.g2_1_0_cascade_\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__13156\,
            I => \this_vga_signals.g2_0_cascade_\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__13153\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1_cascade_\
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__13150\,
            I => \N__13147\
        );

    \I__993\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13144\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__13144\,
            I => \N__13141\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__13141\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0\
        );

    \I__990\ : InMux
    port map (
            O => \N__13138\,
            I => \N__13135\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__13135\,
            I => \N__13132\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__13132\,
            I => \this_vga_signals.g1_0\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__13126\,
            I => \this_vga_signals.g3_1_cascade_\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__13123\,
            I => \this_vga_signals.mult1_un54_sum_ac0_2_mb_rn_0_cascade_\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__13120\,
            I => \this_vga_signals.mult1_un54_sum_axb1_cascade_\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__13117\,
            I => \this_vga_signals.g1_1_cascade_\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__13114\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1_0_cascade_\
        );

    \IN_MUX_bfv_24_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_21_0_\
        );

    \IN_MUX_bfv_24_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_ext_address_q_cry_7\,
            carryinitout => \bfn_24_22_0_\
        );

    \IN_MUX_bfv_21_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_20_0_\
        );

    \IN_MUX_bfv_21_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_oam_data_1_cry_7\,
            carryinitout => \bfn_21_21_0_\
        );

    \IN_MUX_bfv_21_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_23_0_\
        );

    \IN_MUX_bfv_21_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_voffset_d_cry_7\,
            carryinitout => \bfn_21_24_0_\
        );

    \IN_MUX_bfv_20_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_24_0_\
        );

    \IN_MUX_bfv_22_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_21_0_\
        );

    \IN_MUX_bfv_22_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_oam_cache_read_data_3_cry_7\,
            carryinitout => \bfn_22_22_0_\
        );

    \IN_MUX_bfv_20_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_19_0_\
        );

    \IN_MUX_bfv_20_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_oam_cache_read_data_2_cry_7\,
            carryinitout => \bfn_20_20_0_\
        );

    \IN_MUX_bfv_22_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_18_0_\
        );

    \IN_MUX_bfv_22_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_hoffset_q_cry_7\,
            carryinitout => \bfn_22_19_0_\
        );

    \IN_MUX_bfv_19_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_17_0_\
        );

    \IN_MUX_bfv_19_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_hoffset_d_cry_7\,
            carryinitout => \bfn_19_18_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_21_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_22_0_\
        );

    \IN_MUX_bfv_22_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_24_0_\
        );

    \IN_MUX_bfv_22_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_voffset_q_cry_7\,
            carryinitout => \bfn_22_25_0_\
        );

    \IN_MUX_bfv_21_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_18_0_\
        );

    \IN_MUX_bfv_21_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_hoffset_q_2_cry_7\,
            carryinitout => \bfn_21_19_0_\
        );

    \IN_MUX_bfv_21_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_17_0_\
        );

    \IN_MUX_bfv_19_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_13_0_\
        );

    \IN_MUX_bfv_19_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_spr_address_q_cry_7\,
            carryinitout => \bfn_19_14_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_9_22_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR1G77_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__13264\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_935_0_g\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19210\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_1212_g\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23974\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22600\,
            GLOBALBUFFEROUTPUT => \N_504_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI93SL3_6_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001101001"
        )
    port map (
            in0 => \N__17404\,
            in1 => \N__16133\,
            in2 => \N__13408\,
            in3 => \N__16603\,
            lcout => \this_vga_signals.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIDHDA1_1_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__15673\,
            in1 => \N__15400\,
            in2 => \_gnd_net_\,
            in3 => \N__15599\,
            lcout => \this_vga_signals.vaddress_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_RNI0SND1_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111100000000"
        )
    port map (
            in0 => \N__15205\,
            in1 => \N__16580\,
            in2 => \N__13597\,
            in3 => \N__13563\,
            lcout => \this_vga_signals.N_32_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_a5_1_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__15856\,
            in1 => \N__14695\,
            in2 => \N__16858\,
            in3 => \N__14582\,
            lcout => \this_vga_signals.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011101101101"
        )
    port map (
            in0 => \N__13709\,
            in1 => \N__16841\,
            in2 => \N__17576\,
            in3 => \N__14285\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110110000100"
        )
    port map (
            in0 => \N__14959\,
            in1 => \N__15490\,
            in2 => \N__13117\,
            in3 => \N__15620\,
            lcout => \this_vga_signals.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17475\,
            in2 => \_gnd_net_\,
            in3 => \N__16836\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_20_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17530\,
            in1 => \N__16840\,
            in2 => \_gnd_net_\,
            in3 => \N__14284\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100011"
        )
    port map (
            in0 => \N__14958\,
            in1 => \N__14075\,
            in2 => \N__13114\,
            in3 => \N__13710\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_2_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111011"
        )
    port map (
            in0 => \N__13429\,
            in1 => \N__15480\,
            in2 => \N__13129\,
            in3 => \N__13853\,
            lcout => \this_vga_signals.g3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010110111"
        )
    port map (
            in0 => \N__16846\,
            in1 => \N__17390\,
            in2 => \N__17569\,
            in3 => \N__14692\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101101"
        )
    port map (
            in0 => \N__14282\,
            in1 => \N__17516\,
            in2 => \N__16859\,
            in3 => \N__13704\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__14953\,
            in1 => \N__13138\,
            in2 => \N__13126\,
            in3 => \N__14283\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_rn_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100110010000"
        )
    port map (
            in0 => \N__15765\,
            in1 => \N__15838\,
            in2 => \N__13795\,
            in3 => \N__14570\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_2_mb_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_mb_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14691\,
            in2 => \N__13123\,
            in3 => \N__13639\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14386\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40414\,
            ce => \N__16293\,
            sr => \N__16261\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17512\,
            in1 => \N__16842\,
            in2 => \_gnd_net_\,
            in3 => \N__14281\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010011"
        )
    port map (
            in0 => \N__17520\,
            in1 => \N__14952\,
            in2 => \N__13120\,
            in3 => \N__13703\,
            lcout => \this_vga_signals.if_N_9_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_i_o2_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16778\,
            lcout => \this_vga_signals.g2_1_0\,
            ltout => \this_vga_signals.g2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101111"
        )
    port map (
            in0 => \N__14950\,
            in1 => \N__17590\,
            in2 => \N__13159\,
            in3 => \N__13708\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110011010"
        )
    port map (
            in0 => \N__13653\,
            in1 => \N__14065\,
            in2 => \N__13156\,
            in3 => \N__13986\,
            lcout => \this_vga_signals.mult1_un61_sum_axb2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__15837\,
            in1 => \N__15772\,
            in2 => \_gnd_net_\,
            in3 => \N__14264\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_1\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_12_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001101"
        )
    port map (
            in0 => \N__13706\,
            in1 => \N__14951\,
            in2 => \N__13153\,
            in3 => \N__14064\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_0_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110001"
        )
    port map (
            in0 => \N__16779\,
            in1 => \N__13705\,
            in2 => \N__17598\,
            in3 => \N__14266\,
            lcout => \this_vga_signals.g3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_0_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111101111"
        )
    port map (
            in0 => \N__17389\,
            in1 => \N__14696\,
            in2 => \N__13150\,
            in3 => \N__14583\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010001"
        )
    port map (
            in0 => \N__14063\,
            in1 => \N__13707\,
            in2 => \N__14973\,
            in3 => \N__13746\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__17392\,
            in1 => \N__17563\,
            in2 => \N__16822\,
            in3 => \N__14705\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14302\,
            in3 => \N__16774\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__13970\,
            in1 => \_gnd_net_\,
            in2 => \N__13183\,
            in3 => \N__15627\,
            lcout => \this_vga_signals.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_0_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13969\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => \this_vga_signals.g1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_x0_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110111"
        )
    port map (
            in0 => \N__13971\,
            in1 => \N__15476\,
            in2 => \N__13180\,
            in3 => \N__14011\,
            lcout => \this_vga_signals.g3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14356\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40428\,
            ce => \N__16292\,
            sr => \N__16263\
        );

    \this_vga_signals.un5_vaddress_g3_x1_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111111111"
        )
    port map (
            in0 => \N__13972\,
            in1 => \N__14012\,
            in2 => \N__15520\,
            in3 => \N__13177\,
            lcout => \this_vga_signals.g3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14355\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40428\,
            ce => \N__16292\,
            sr => \N__16263\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__17567\,
            in1 => \N__13887\,
            in2 => \N__15513\,
            in3 => \N__13976\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI1NB793_6_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13171\,
            in1 => \N__14118\,
            in2 => \N__13162\,
            in3 => \N__13278\,
            lcout => \this_vga_signals.g2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__17566\,
            in1 => \N__13886\,
            in2 => \N__15512\,
            in3 => \N__13974\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13852\,
            in1 => \N__13327\,
            in2 => \N__14748\,
            in3 => \N__13195\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axb1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__15688\,
            in1 => \N__13258\,
            in2 => \N__13249\,
            in3 => \N__13801\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBN8KM1_4_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13975\,
            in1 => \N__13246\,
            in2 => \N__13898\,
            in3 => \N__17568\,
            lcout => \this_vga_signals.vaddress_m2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m1_0_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17565\,
            in1 => \N__13973\,
            in2 => \_gnd_net_\,
            in3 => \N__13885\,
            lcout => \this_vga_signals.if_m1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000001111"
        )
    port map (
            in0 => \N__15632\,
            in1 => \N__13234\,
            in2 => \N__15516\,
            in3 => \N__13225\,
            lcout => \this_vga_signals.mult1_un68_sum_c3\,
            ltout => \this_vga_signals.mult1_un68_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_3_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15008\,
            in1 => \N__13912\,
            in2 => \N__13219\,
            in3 => \N__13194\,
            lcout => \this_vga_signals.g2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__13216\,
            in1 => \N__14125\,
            in2 => \N__15517\,
            in3 => \N__14020\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000000000"
        )
    port map (
            in0 => \N__13207\,
            in1 => \N__15687\,
            in2 => \N__13201\,
            in3 => \N__14189\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_3_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_1_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101101001"
        )
    port map (
            in0 => \N__17585\,
            in1 => \N__15621\,
            in2 => \N__15515\,
            in3 => \N__13990\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axb1_3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001111000"
        )
    port map (
            in0 => \N__15505\,
            in1 => \N__17586\,
            in2 => \N__13198\,
            in3 => \N__13900\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13899\,
            in1 => \N__15007\,
            in2 => \N__14980\,
            in3 => \N__13991\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_14_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13992\,
            in1 => \N__15498\,
            in2 => \N__13369\,
            in3 => \N__15633\,
            lcout => \this_vga_signals.g0_0_0_a2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_4_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13612\,
            in1 => \N__14223\,
            in2 => \N__13357\,
            in3 => \N__13325\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__15052\,
            in1 => \N__14744\,
            in2 => \N__13345\,
            in3 => \N__14169\,
            lcout => \this_vga_signals.if_i4_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__16915\,
            in1 => \N__17002\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNILB7N84_2_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010011101011"
        )
    port map (
            in0 => \N__13326\,
            in1 => \N__15637\,
            in2 => \N__15519\,
            in3 => \N__13312\,
            lcout => \this_vga_signals.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13303\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110101001110"
        )
    port map (
            in0 => \N__14098\,
            in1 => \N__13291\,
            in2 => \N__15518\,
            in3 => \N__13282\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20064\,
            in2 => \_gnd_net_\,
            in3 => \N__16267\,
            lcout => \this_vga_signals.N_935_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.port_data_rw_0_i_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__29223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32217\,
            lcout => port_data_rw_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUQPR1_7_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010001001011"
        )
    port map (
            in0 => \N__17570\,
            in1 => \N__16860\,
            in2 => \N__14134\,
            in3 => \N__16708\,
            lcout => \this_vga_signals.g2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16976\,
            in2 => \_gnd_net_\,
            in3 => \N__17059\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__17020\,
            in1 => \_gnd_net_\,
            in2 => \N__16992\,
            in3 => \_gnd_net_\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_0_9_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000010001"
        )
    port map (
            in0 => \N__13447\,
            in1 => \N__14415\,
            in2 => \N__13468\,
            in3 => \N__15139\,
            lcout => \this_vga_signals.SUM_2_i_i_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_9_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40385\,
            ce => \N__16298\,
            sr => \N__16255\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16313\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40385\,
            ce => \N__16298\,
            sr => \N__16255\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15869\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40385\,
            ce => \N__16298\,
            sr => \N__16255\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_N_2L1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__14430\,
            in1 => \N__13506\,
            in2 => \N__13542\,
            in3 => \N__14414\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_2_2_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14375\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40385\,
            ce => \N__16298\,
            sr => \N__16255\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14452\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40385\,
            ce => \N__16298\,
            sr => \N__16255\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14346\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40385\,
            ce => \N__16298\,
            sr => \N__16255\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_9_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011110101111"
        )
    port map (
            in0 => \N__15136\,
            in1 => \N__13445\,
            in2 => \N__13467\,
            in3 => \N__14413\,
            lcout => \this_vga_signals.SUM_2_i_i_1_0_3\,
            ltout => \this_vga_signals.SUM_2_i_i_1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__15184\,
            in1 => \N__15255\,
            in2 => \N__13450\,
            in3 => \N__16565\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13541\,
            in3 => \N__13504\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_x1_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__13446\,
            in1 => \N__15256\,
            in2 => \N__15314\,
            in3 => \N__15137\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_2_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_ns_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__16566\,
            in1 => \_gnd_net_\,
            in2 => \N__13432\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_2_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13993\,
            in3 => \N__17529\,
            lcout => \this_vga_signals.g1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__15138\,
            in1 => \N__13505\,
            in2 => \N__15270\,
            in3 => \N__15305\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_ns_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__13570\,
            in1 => \_gnd_net_\,
            in2 => \N__13600\,
            in3 => \N__13534\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_ns_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13596\,
            in2 => \N__13579\,
            in3 => \N__13549\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x0_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__15253\,
            in1 => \N__15140\,
            in2 => \N__15313\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000110010100"
        )
    port map (
            in0 => \N__14569\,
            in1 => \N__13794\,
            in2 => \N__13633\,
            in3 => \N__14693\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x1_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000111001"
        )
    port map (
            in0 => \N__15183\,
            in1 => \N__15260\,
            in2 => \N__13564\,
            in3 => \N__16567\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_x1_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15141\,
            in1 => \N__13543\,
            in2 => \N__15200\,
            in3 => \N__15254\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_ns_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13513\,
            in3 => \N__13510\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__13486\,
            in1 => \N__14458\,
            in2 => \N__13480\,
            in3 => \N__13477\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101010101"
        )
    port map (
            in0 => \N__13793\,
            in1 => \N__13628\,
            in2 => \N__13471\,
            in3 => \N__14568\,
            lcout => \this_vga_signals.mult1_un47_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_sn_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000100000000"
        )
    port map (
            in0 => \N__15763\,
            in1 => \N__13632\,
            in2 => \N__15839\,
            in3 => \N__14565\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_2_mb_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__15821\,
            in1 => \N__15757\,
            in2 => \_gnd_net_\,
            in3 => \N__15263\,
            lcout => \this_vga_signals.r_N_4_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14382\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40419\,
            ce => \N__16294\,
            sr => \N__16262\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001110111"
        )
    port map (
            in0 => \N__15823\,
            in1 => \N__15761\,
            in2 => \_gnd_net_\,
            in3 => \N__15261\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011010"
        )
    port map (
            in0 => \N__15262\,
            in1 => \_gnd_net_\,
            in2 => \N__15773\,
            in3 => \N__15822\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc1_0\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010100"
        )
    port map (
            in0 => \N__14566\,
            in1 => \N__14694\,
            in2 => \N__13615\,
            in3 => \N__13792\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_0_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010011111"
        )
    port map (
            in0 => \N__15762\,
            in1 => \N__15824\,
            in2 => \N__17403\,
            in3 => \N__14690\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_a5_1_3_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14567\,
            in1 => \N__17399\,
            in2 => \_gnd_net_\,
            in3 => \N__15764\,
            lcout => \this_vga_signals.g0_0_i_a5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001101"
        )
    port map (
            in0 => \N__13747\,
            in1 => \N__14974\,
            in2 => \N__13717\,
            in3 => \N__14062\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_3_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13968\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17572\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_3_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111101"
        )
    port map (
            in0 => \N__15491\,
            in1 => \N__13813\,
            in2 => \N__13807\,
            in3 => \N__13851\,
            lcout => \this_vga_signals.g3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000101"
        )
    port map (
            in0 => \N__14061\,
            in1 => \N__14960\,
            in2 => \N__13748\,
            in3 => \N__13711\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14013\,
            in2 => \N__13804\,
            in3 => \N__13967\,
            lcout => \this_vga_signals.mult1_un61_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_0_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16046\,
            in1 => \N__14485\,
            in2 => \_gnd_net_\,
            in3 => \N__14813\,
            lcout => \this_vga_signals.g0_0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14592\,
            in1 => \N__13791\,
            in2 => \N__14301\,
            in3 => \N__13762\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_1_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13753\,
            in3 => \N__17571\,
            lcout => \this_vga_signals.g1_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_1_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__13715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13749\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001101"
        )
    port map (
            in0 => \N__13750\,
            in1 => \N__14961\,
            in2 => \N__14082\,
            in3 => \N__13716\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_0_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__13985\,
            in1 => \N__14626\,
            in2 => \N__13660\,
            in3 => \N__13657\,
            lcout => \this_vga_signals.g0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_6_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14293\,
            in1 => \N__14119\,
            in2 => \N__16531\,
            in3 => \N__16161\,
            lcout => \this_vga_signals.g0_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100110"
        )
    port map (
            in0 => \N__14089\,
            in1 => \N__14969\,
            in2 => \N__14083\,
            in3 => \N__14032\,
            lcout => \this_vga_signals.N_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_4_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__14014\,
            in1 => \N__13891\,
            in2 => \_gnd_net_\,
            in3 => \N__13984\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_0_0_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14962\,
            in1 => \N__16780\,
            in2 => \_gnd_net_\,
            in3 => \N__14292\,
            lcout => \this_vga_signals.g2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_ns_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13906\,
            in1 => \N__13892\,
            in2 => \_gnd_net_\,
            in3 => \N__13861\,
            lcout => \this_vga_signals.g3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13855\,
            in1 => \N__14217\,
            in2 => \N__15040\,
            in3 => \N__14738\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14979\,
            in1 => \N__15013\,
            in2 => \N__16855\,
            in3 => \N__14304\,
            lcout => \this_vga_signals.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001100"
        )
    port map (
            in0 => \N__13854\,
            in1 => \N__14599\,
            in2 => \N__13822\,
            in3 => \N__14812\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14740\,
            in1 => \N__14227\,
            in2 => \N__14323\,
            in3 => \N__14320\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7RTI411_2_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110011010"
        )
    port map (
            in0 => \N__14191\,
            in1 => \N__15610\,
            in2 => \N__14314\,
            in3 => \N__14311\,
            lcout => \this_vga_signals.vaddress_m6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_0_a2_3_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14218\,
            in1 => \N__16823\,
            in2 => \_gnd_net_\,
            in3 => \N__14303\,
            lcout => \this_vga_signals.g0_6_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_0_a2_2_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14305\,
            in1 => \N__14219\,
            in2 => \N__16854\,
            in3 => \N__14739\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__15609\,
            in1 => \N__14614\,
            in2 => \N__14194\,
            in3 => \N__14190\,
            lcout => \this_vga_signals.mult1_un75_sum_ac0_3_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20510\,
            in1 => \N__17595\,
            in2 => \N__16856\,
            in3 => \N__16408\,
            lcout => \this_vga_signals.vsync_1_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIGAFCKA_2_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011000110"
        )
    port map (
            in0 => \N__15631\,
            in1 => \N__14176\,
            in2 => \N__15514\,
            in3 => \N__14170\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_N_3_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI0FQEQV_2_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000111"
        )
    port map (
            in0 => \N__14158\,
            in1 => \N__14152\,
            in2 => \N__14146\,
            in3 => \N__14143\,
            lcout => \this_vga_signals.M_vcounter_q_RNI0FQEQVZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICSHP_6_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15380\,
            in2 => \_gnd_net_\,
            in3 => \N__17393\,
            lcout => \this_vga_signals.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20068\,
            in1 => \N__15339\,
            in2 => \N__19894\,
            in3 => \N__19890\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__40378\,
            ce => 'H',
            sr => \N__16254\
        );

    \this_vga_signals.M_vcounter_q_1_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20070\,
            in1 => \N__15672\,
            in2 => \_gnd_net_\,
            in3 => \N__14395\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__40378\,
            ce => 'H',
            sr => \N__16254\
        );

    \this_vga_signals.M_vcounter_q_2_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20069\,
            in1 => \N__15576\,
            in2 => \_gnd_net_\,
            in3 => \N__14392\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__40378\,
            ce => 'H',
            sr => \N__16254\
        );

    \this_vga_signals.M_vcounter_q_3_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20071\,
            in1 => \N__15422\,
            in2 => \_gnd_net_\,
            in3 => \N__14389\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__40378\,
            ce => 'H',
            sr => \N__16254\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17596\,
            in2 => \_gnd_net_\,
            in3 => \N__14359\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16857\,
            in2 => \_gnd_net_\,
            in3 => \N__14335\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17394\,
            in2 => \_gnd_net_\,
            in3 => \N__14332\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16706\,
            in2 => \_gnd_net_\,
            in3 => \N__14329\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16397\,
            in2 => \_gnd_net_\,
            in3 => \N__14326\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20484\,
            in2 => \_gnd_net_\,
            in3 => \N__14473\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15917\,
            lcout => \this_vga_signals.M_vcounter_q_9_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40386\,
            ce => \N__16299\,
            sr => \N__16256\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14450\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40386\,
            ce => \N__16299\,
            sr => \N__16256\
        );

    \this_vga_signals.un5_vaddress_g0_0_3_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14954\,
            in2 => \_gnd_net_\,
            in3 => \N__15012\,
            lcout => \this_vga_signals.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101111001101"
        )
    port map (
            in0 => \N__16376\,
            in1 => \N__15185\,
            in2 => \N__14470\,
            in3 => \N__15306\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16320\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40398\,
            ce => \N__16296\,
            sr => \N__16258\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14451\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals_M_vcounter_q_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40398\,
            ce => \N__16296\,
            sr => \N__16258\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15876\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40398\,
            ce => \N__16296\,
            sr => \N__16258\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_1_a0_1_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14434\,
            in2 => \_gnd_net_\,
            in3 => \N__14419\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_1_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011111101111"
        )
    port map (
            in0 => \N__15316\,
            in1 => \N__16688\,
            in2 => \N__14512\,
            in3 => \N__15699\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_c2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__16594\,
            in1 => \N__14479\,
            in2 => \N__14509\,
            in3 => \N__14500\,
            lcout => \this_vga_signals.mult1_un40_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_18_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__15934\,
            in1 => \_gnd_net_\,
            in2 => \N__14506\,
            in3 => \N__16156\,
            lcout => \this_vga_signals.N_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIOKSG_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16378\,
            in2 => \_gnd_net_\,
            in3 => \N__15268\,
            lcout => \this_vga_signals.vaddress_m2_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_15_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16179\,
            in1 => \N__16155\,
            in2 => \_gnd_net_\,
            in3 => \N__16097\,
            lcout => \this_vga_signals.g0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_1_0_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011011101"
        )
    port map (
            in0 => \N__15198\,
            in1 => \N__16377\,
            in2 => \_gnd_net_\,
            in3 => \N__15315\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_c2_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__15269\,
            in1 => \_gnd_net_\,
            in2 => \N__14503\,
            in3 => \N__16593\,
            lcout => \this_vga_signals.mult1_un40_sum_c2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_5_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010111101111"
        )
    port map (
            in0 => \N__14494\,
            in1 => \N__14591\,
            in2 => \N__17251\,
            in3 => \N__16024\,
            lcout => \this_vga_signals.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001100000"
        )
    port map (
            in0 => \N__15201\,
            in1 => \N__16590\,
            in2 => \N__15109\,
            in3 => \N__15271\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16591\,
            in1 => \N__14590\,
            in2 => \N__17380\,
            in3 => \N__14706\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_a5_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__14707\,
            in1 => \N__14647\,
            in2 => \N__16853\,
            in3 => \N__15888\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_2_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__15889\,
            in1 => \N__14641\,
            in2 => \N__14629\,
            in3 => \N__16023\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_8_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101111110"
        )
    port map (
            in0 => \N__16705\,
            in1 => \N__16592\,
            in2 => \N__16407\,
            in3 => \N__17350\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__16180\,
            in1 => \N__16160\,
            in2 => \_gnd_net_\,
            in3 => \N__16099\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_1_0_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__14814\,
            in1 => \N__14878\,
            in2 => \N__16003\,
            in3 => \N__14620\,
            lcout => \this_vga_signals.g3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000101010"
        )
    port map (
            in0 => \N__16056\,
            in1 => \N__16071\,
            in2 => \N__14608\,
            in3 => \N__16026\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_1_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17594\,
            in1 => \N__17345\,
            in2 => \_gnd_net_\,
            in3 => \N__14593\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__16055\,
            in1 => \N__14524\,
            in2 => \N__14515\,
            in3 => \N__16025\,
            lcout => \this_vga_signals.g0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_0_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__15423\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15597\,
            lcout => \this_vga_signals.mult1_un75_sum_axb2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17113\,
            in2 => \_gnd_net_\,
            in3 => \N__16993\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI87V41_7_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16707\,
            in1 => \N__17346\,
            in2 => \_gnd_net_\,
            in3 => \N__15598\,
            lcout => \this_vga_signals.vsync_1_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g3_0_1_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15006\,
            in2 => \_gnd_net_\,
            in3 => \N__14978\,
            lcout => \this_vga_signals.g3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_9_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14713\,
            in2 => \N__14872\,
            in3 => \N__14863\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_c3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIU4E93J3_8_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__15988\,
            in1 => \N__14854\,
            in2 => \N__14848\,
            in3 => \N__14845\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_13_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__14815\,
            in1 => \N__14791\,
            in2 => \N__14782\,
            in3 => \N__14773\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_12_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011110111101"
        )
    port map (
            in0 => \N__14767\,
            in1 => \N__14758\,
            in2 => \N__14752\,
            in3 => \N__14749\,
            lcout => \this_vga_signals.g0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17001\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__15680\,
            in1 => \N__15082\,
            in2 => \N__15073\,
            in3 => \N__15424\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_8_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15679\,
            in2 => \_gnd_net_\,
            in3 => \N__15340\,
            lcout => \this_vga_signals.if_N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__20077\,
            in1 => \N__18324\,
            in2 => \_gnd_net_\,
            in3 => \N__18376\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40353\,
            ce => 'H',
            sr => \N__16515\
        );

    \this_vga_signals.M_hcounter_q_0_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20076\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40353\,
            ce => 'H',
            sr => \N__16515\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__18987\,
            in1 => \N__18185\,
            in2 => \_gnd_net_\,
            in3 => \N__18112\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000010011"
        )
    port map (
            in0 => \N__18990\,
            in1 => \N__18187\,
            in2 => \N__18260\,
            in3 => \N__18234\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__18815\,
            in1 => \N__19055\,
            in2 => \N__18918\,
            in3 => \N__18986\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011100000"
        )
    port map (
            in0 => \N__18988\,
            in1 => \N__18186\,
            in2 => \N__15043\,
            in3 => \N__18113\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001011110"
        )
    port map (
            in0 => \N__18989\,
            in1 => \N__18114\,
            in2 => \N__18204\,
            in3 => \N__18233\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010001"
        )
    port map (
            in0 => \N__15721\,
            in1 => \N__18251\,
            in2 => \N__15715\,
            in3 => \N__15712\,
            lcout => \this_vga_signals.mult1_un61_sum_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010111010111"
        )
    port map (
            in0 => \N__18809\,
            in1 => \N__19054\,
            in2 => \N__18917\,
            in3 => \N__18991\,
            lcout => \this_vga_signals.SUM_3_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_0_8_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001111111"
        )
    port map (
            in0 => \N__16702\,
            in1 => \N__16380\,
            in2 => \N__17395\,
            in3 => \N__16601\,
            lcout => OPEN,
            ltout => \this_vga_signals.vvisibility_i_o2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_9_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000101010001"
        )
    port map (
            in0 => \N__20483\,
            in1 => \N__16703\,
            in2 => \N__15706\,
            in3 => \N__15703\,
            lcout => \N_825_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17375\,
            in1 => \N__16698\,
            in2 => \N__16870\,
            in3 => \N__16379\,
            lcout => \this_vga_signals.M_lcounter_q_3_i_o2_2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__15660\,
            in1 => \N__15550\,
            in2 => \N__15399\,
            in3 => \N__15335\,
            lcout => \this_vga_signals.N_822_0\,
            ltout => \this_vga_signals.N_822_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__16869\,
            in1 => \N__17379\,
            in2 => \N__15319\,
            in3 => \N__17583\,
            lcout => this_vga_signals_un4_lvisibility_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__15307\,
            in1 => \N__15264\,
            in2 => \N__15199\,
            in3 => \N__15142\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__17368\,
            in1 => \N__15844\,
            in2 => \_gnd_net_\,
            in3 => \N__15784\,
            lcout => OPEN,
            ltout => \this_vga_signals.r_N_4_mux_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI767P1_1_9_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011011110011"
        )
    port map (
            in0 => \N__20443\,
            in1 => \N__16680\,
            in2 => \N__15937\,
            in3 => \N__16381\,
            lcout => \this_vga_signals.N_24_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18393\,
            in1 => \N__18535\,
            in2 => \N__18655\,
            in3 => \N__18331\,
            lcout => OPEN,
            ltout => \this_vga_signals.un2_hsynclt6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18142\,
            in1 => \N__18210\,
            in2 => \N__15925\,
            in3 => \N__19013\,
            lcout => \this_vga_signals.un2_hsynclt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15922\,
            lcout => \this_vga_signals_M_vcounter_q_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40399\,
            ce => \N__16297\,
            sr => \N__16259\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI539J1_9_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001011011101"
        )
    port map (
            in0 => \N__16686\,
            in1 => \N__15901\,
            in2 => \N__20479\,
            in3 => \N__16387\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_24_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_27_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16154\,
            in2 => \N__15892\,
            in3 => \N__16096\,
            lcout => \this_vga_signals.N_4_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15880\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40408\,
            ce => \N__16295\,
            sr => \N__16260\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_a5_1_0_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17325\,
            lcout => \this_vga_signals.g0_0_i_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__17326\,
            in1 => \N__15840\,
            in2 => \_gnd_net_\,
            in3 => \N__15782\,
            lcout => \this_vga_signals.r_N_4_mux\,
            ltout => \this_vga_signals.r_N_4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI767P1_9_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011011110011"
        )
    port map (
            in0 => \N__20473\,
            in1 => \N__16682\,
            in2 => \N__16183\,
            in3 => \N__16398\,
            lcout => \this_vga_signals.N_24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI767P1_0_9_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011101100101"
        )
    port map (
            in0 => \N__16399\,
            in1 => \N__16168\,
            in2 => \N__16704\,
            in3 => \N__20474\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_24_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16162\,
            in2 => \N__16102\,
            in3 => \N__16098\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_1_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011000100"
        )
    port map (
            in0 => \N__16075\,
            in1 => \N__16060\,
            in2 => \N__16030\,
            in3 => \N__16027\,
            lcout => \this_vga_signals.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3SF72_8_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__18849\,
            in1 => \N__15994\,
            in2 => \N__16450\,
            in3 => \N__19091\,
            lcout => \this_vga_signals.g0_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20025\,
            in2 => \_gnd_net_\,
            in3 => \N__19880\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__16213\,
            in1 => \N__15982\,
            in2 => \N__19099\,
            in3 => \N__18937\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17146\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16997\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101001011001"
        )
    port map (
            in0 => \N__16889\,
            in1 => \N__18127\,
            in2 => \N__18526\,
            in3 => \N__17704\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_8_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18622\,
            in2 => \N__16201\,
            in3 => \N__18375\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_9_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100011101"
        )
    port map (
            in0 => \N__18623\,
            in1 => \N__18507\,
            in2 => \N__16198\,
            in3 => \N__18441\,
            lcout => \this_vga_signals.mult1_un82_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100110010011"
        )
    port map (
            in0 => \N__17705\,
            in1 => \N__16890\,
            in2 => \N__18527\,
            in3 => \N__18128\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__18317\,
            in1 => \N__18364\,
            in2 => \N__18329\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_d7lt4\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20072\,
            in1 => \N__18640\,
            in2 => \_gnd_net_\,
            in3 => \N__16195\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__40354\,
            ce => 'H',
            sr => \N__16516\
        );

    \this_vga_signals.M_hcounter_q_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20065\,
            in1 => \N__18523\,
            in2 => \_gnd_net_\,
            in3 => \N__16192\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__40354\,
            ce => 'H',
            sr => \N__16516\
        );

    \this_vga_signals.M_hcounter_q_4_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20073\,
            in1 => \N__18129\,
            in2 => \_gnd_net_\,
            in3 => \N__16189\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__40354\,
            ce => 'H',
            sr => \N__16516\
        );

    \this_vga_signals.M_hcounter_q_5_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20066\,
            in1 => \N__18197\,
            in2 => \_gnd_net_\,
            in3 => \N__16186\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__40354\,
            ce => 'H',
            sr => \N__16516\
        );

    \this_vga_signals.M_hcounter_q_6_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20074\,
            in1 => \N__19001\,
            in2 => \_gnd_net_\,
            in3 => \N__16429\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__40354\,
            ce => 'H',
            sr => \N__16516\
        );

    \this_vga_signals.M_hcounter_q_7_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20067\,
            in1 => \N__19069\,
            in2 => \_gnd_net_\,
            in3 => \N__16426\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__40354\,
            ce => 'H',
            sr => \N__16516\
        );

    \this_vga_signals.M_hcounter_q_8_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20075\,
            in1 => \N__18819\,
            in2 => \_gnd_net_\,
            in3 => \N__16423\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__40354\,
            ce => 'H',
            sr => \N__16516\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18924\,
            in2 => \_gnd_net_\,
            in3 => \N__16420\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40367\,
            ce => \N__16477\,
            sr => \N__16514\
        );

    \this_vga_signals.un4_haddress_if_m5_i_a4_0_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18534\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18400\,
            lcout => OPEN,
            ltout => \this_vga_signals.un4_hsynclto3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__18644\,
            in1 => \N__18209\,
            in2 => \N__16417\,
            in3 => \N__18140\,
            lcout => \this_vga_signals.un4_hsynclto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_d_0_sqmuxa_1_0_o2_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__16414\,
            in1 => \N__16687\,
            in2 => \_gnd_net_\,
            in3 => \N__16400\,
            lcout => \this_ppu.N_759_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16324\,
            lcout => \this_vga_signals_M_vcounter_q_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40387\,
            ce => \N__16300\,
            sr => \N__16257\
        );

    \this_vga_signals.M_hcounter_q_RNISKQ82_8_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__19092\,
            in1 => \N__16222\,
            in2 => \N__18853\,
            in3 => \N__19014\,
            lcout => \this_vga_signals.un4_hsynclt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_2_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110001100011"
        )
    port map (
            in0 => \N__16818\,
            in1 => \N__16681\,
            in2 => \N__17597\,
            in3 => \N__17343\,
            lcout => \this_vga_signals.g0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_1_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__16609\,
            in1 => \N__17344\,
            in2 => \_gnd_net_\,
            in3 => \N__16602\,
            lcout => \this_vga_signals.g0_0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__16495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20029\,
            lcout => \this_vga_signals.N_935_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16462\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18928\,
            in2 => \_gnd_net_\,
            in3 => \N__20478\,
            lcout => \this_vga_signals.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_0_9_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19718\,
            lcout => \M_vcounter_q_esr_RNIQJSA2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001011010"
        )
    port map (
            in0 => \N__17841\,
            in1 => \_gnd_net_\,
            in2 => \N__17901\,
            in3 => \N__17952\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010011"
        )
    port map (
            in0 => \N__17995\,
            in1 => \N__17960\,
            in2 => \N__17852\,
            in3 => \N__17897\,
            lcout => \this_vga_ramdac.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100010111"
        )
    port map (
            in0 => \N__17892\,
            in1 => \N__17853\,
            in2 => \N__17962\,
            in3 => \N__17997\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100100101011"
        )
    port map (
            in0 => \N__17998\,
            in1 => \N__17842\,
            in2 => \N__17961\,
            in3 => \N__17891\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18571\,
            in1 => \N__17671\,
            in2 => \N__17041\,
            in3 => \N__18444\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111101"
        )
    port map (
            in0 => \N__17996\,
            in1 => \N__17956\,
            in2 => \N__17857\,
            in3 => \N__17893\,
            lcout => \this_vga_ramdac.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIFBB7K_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111010"
        )
    port map (
            in0 => \N__18624\,
            in1 => \N__18383\,
            in2 => \N__18528\,
            in3 => \N__18427\,
            lcout => OPEN,
            ltout => \this_vga_signals.d_N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_am_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000011110000"
        )
    port map (
            in0 => \N__18384\,
            in1 => \N__18625\,
            in2 => \N__17032\,
            in3 => \N__17733\,
            lcout => \this_vga_signals.mult1_un89_sum_axbxc3_2_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__17029\,
            in1 => \N__17650\,
            in2 => \N__17019\,
            in3 => \N__23973\,
            lcout => \this_vga_ramdac.N_2687_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__17646\,
            in1 => \N__18049\,
            in2 => \N__16959\,
            in3 => \N__23956\,
            lcout => \this_vga_ramdac.N_28_i_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__17645\,
            in1 => \N__16924\,
            in2 => \N__16908\,
            in3 => \N__23955\,
            lcout => \this_vga_ramdac.N_2690_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100110011101"
        )
    port map (
            in0 => \N__16891\,
            in1 => \N__18116\,
            in2 => \N__18525\,
            in3 => \N__17706\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17707\,
            in1 => \N__18064\,
            in2 => \N__16873\,
            in3 => \N__18268\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__18607\,
            in1 => \N__17152\,
            in2 => \N__18524\,
            in3 => \N__18115\,
            lcout => \this_vga_signals.M_hcounter_d7lt7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18500\,
            in1 => \N__18117\,
            in2 => \_gnd_net_\,
            in3 => \N__17708\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__17644\,
            in1 => \N__17803\,
            in2 => \N__17139\,
            in3 => \N__23960\,
            lcout => \this_vga_ramdac.N_2691_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19159\,
            in2 => \_gnd_net_\,
            in3 => \N__18282\,
            lcout => \this_vga_signals.pixel_clk_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__17643\,
            in1 => \N__17122\,
            in2 => \N__17106\,
            in3 => \N__23959\,
            lcout => \this_vga_ramdac.N_2689_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17089\,
            in1 => \N__17080\,
            in2 => \_gnd_net_\,
            in3 => \N__17599\,
            lcout => \this_vga_signals.N_819_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__18196\,
            in1 => \N__19053\,
            in2 => \_gnd_net_\,
            in3 => \N__18997\,
            lcout => \this_vga_signals.M_lcounter_q_3_i_o2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNI4VLK7_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19179\,
            in1 => \N__19158\,
            in2 => \_gnd_net_\,
            in3 => \N__18281\,
            lcout => \M_pcounter_q_ret_1_RNI4VLK7\,
            ltout => \M_pcounter_q_ret_1_RNI4VLK7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__17052\,
            in1 => \N__17071\,
            in2 => \N__17062\,
            in3 => \N__23957\,
            lcout => \this_vga_ramdac.N_2686_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__23958\,
            in1 => \N__17659\,
            in2 => \N__17616\,
            in3 => \N__17642\,
            lcout => \this_vga_ramdac.N_2688_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40355\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17584\,
            in2 => \_gnd_net_\,
            in3 => \N__17391\,
            lcout => \this_vga_signals.g0_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__19134\,
            in1 => \N__20057\,
            in2 => \N__19183\,
            in3 => \N__19849\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40368\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__19098\,
            in1 => \N__18936\,
            in2 => \_gnd_net_\,
            in3 => \N__18848\,
            lcout => \M_hcounter_q_esr_RNIU8TO_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI63POP1_9_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18057\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI4UV2O8_9_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__17752\,
            in1 => \N__17179\,
            in2 => \N__18058\,
            in3 => \N__17782\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI4GRFM_9_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18051\,
            in2 => \_gnd_net_\,
            in3 => \N__18448\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI50QR8_9_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18056\,
            in2 => \_gnd_net_\,
            in3 => \N__17719\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI4T6U44_9_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__18052\,
            in1 => \N__17178\,
            in2 => \_gnd_net_\,
            in3 => \N__17772\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI7U1Q5_9_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18220\,
            in2 => \_gnd_net_\,
            in3 => \N__18050\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001001110101"
        )
    port map (
            in0 => \N__17994\,
            in1 => \N__17943\,
            in2 => \N__17902\,
            in3 => \N__17846\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001010110100"
        )
    port map (
            in0 => \N__18570\,
            in1 => \N__17670\,
            in2 => \N__17743\,
            in3 => \N__18443\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m5_i_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011001100100"
        )
    port map (
            in0 => \N__18646\,
            in1 => \N__18397\,
            in2 => \N__18547\,
            in3 => \N__18442\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_2_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.haddress_1_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__17677\,
            in1 => \N__17765\,
            in2 => \N__17791\,
            in3 => \N__17788\,
            lcout => \this_vga_signals.haddress_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000101111011"
        )
    port map (
            in0 => \N__17766\,
            in1 => \N__18398\,
            in2 => \N__18654\,
            in3 => \N__18292\,
            lcout => \this_vga_signals.mult1_un89_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_bm_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17739\,
            in1 => \N__18141\,
            in2 => \_gnd_net_\,
            in3 => \N__17715\,
            lcout => \this_vga_signals.mult1_un89_sum_axbxc3_2_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111011"
        )
    port map (
            in0 => \N__18542\,
            in1 => \N__18645\,
            in2 => \_gnd_net_\,
            in3 => \N__18428\,
            lcout => \this_vga_signals.mult1_un75_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_x4_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100110110"
        )
    port map (
            in0 => \N__18650\,
            in1 => \N__18563\,
            in2 => \N__18546\,
            in3 => \N__18429\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_8_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18399\,
            in2 => \N__18334\,
            in3 => \N__18330\,
            lcout => \this_vga_signals.if_N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18283\,
            lcout => \this_vga_signals.M_pcounter_q_i_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19135\,
            in1 => \N__19146\,
            in2 => \_gnd_net_\,
            in3 => \N__19839\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20006\,
            in1 => \_gnd_net_\,
            in2 => \N__18286\,
            in3 => \N__19108\,
            lcout => \this_vga_signals.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111010001100"
        )
    port map (
            in0 => \N__18267\,
            in1 => \N__18238\,
            in2 => \N__18211\,
            in3 => \N__19008\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110100110"
        )
    port map (
            in0 => \N__19009\,
            in1 => \N__18208\,
            in2 => \N__18145\,
            in3 => \N__18133\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIOSP33_9_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__18920\,
            in1 => \N__18840\,
            in2 => \N__19710\,
            in3 => \N__19097\,
            lcout => \N_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__18019\,
            in1 => \N__18919\,
            in2 => \N__19192\,
            in3 => \N__18839\,
            lcout => \this_vga_signals.N_83_1\,
            ltout => \this_vga_signals.N_83_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNIGO4F3_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__20030\,
            in1 => \N__19178\,
            in2 => \N__19162\,
            in3 => \N__19132\,
            lcout => \this_vga_signals.N_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19150\,
            in1 => \N__19133\,
            in2 => \_gnd_net_\,
            in3 => \N__19848\,
            lcout => \this_vga_signals.M_pcounter_q_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40356\,
            ce => \N__20063\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19096\,
            in2 => \_gnd_net_\,
            in3 => \N__19015\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_809_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIT8TC3_9_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__19711\,
            in1 => \N__18932\,
            in2 => \N__18856\,
            in3 => \N__18847\,
            lcout => \N_34_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI5I298_9_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__29229\,
            in1 => \N__37753\,
            in2 => \_gnd_net_\,
            in3 => \N__19719\,
            lcout => port_nmib_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_0_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22858\,
            in1 => \N__18729\,
            in2 => \N__22160\,
            in3 => \N__22136\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_1_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22864\,
            in1 => \N__18702\,
            in2 => \_gnd_net_\,
            in3 => \N__18688\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_2_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22859\,
            in1 => \N__18672\,
            in2 => \_gnd_net_\,
            in3 => \N__18658\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_3_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22865\,
            in1 => \N__19398\,
            in2 => \_gnd_net_\,
            in3 => \N__19384\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_4_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22860\,
            in1 => \N__19368\,
            in2 => \_gnd_net_\,
            in3 => \N__19354\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_5_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22862\,
            in1 => \N__19341\,
            in2 => \_gnd_net_\,
            in3 => \N__19327\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_6_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22861\,
            in1 => \N__19314\,
            in2 => \_gnd_net_\,
            in3 => \N__19300\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_7_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22863\,
            in1 => \N__19284\,
            in2 => \_gnd_net_\,
            in3 => \N__19270\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \N__40436\,
            ce => 'H',
            sr => \N__28898\
        );

    \M_this_map_address_q_8_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22866\,
            in1 => \N__19254\,
            in2 => \_gnd_net_\,
            in3 => \N__19240\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \N__40444\,
            ce => 'H',
            sr => \N__28896\
        );

    \M_this_map_address_q_9_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__19224\,
            in1 => \N__22867\,
            in2 => \_gnd_net_\,
            in3 => \N__19237\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40444\,
            ce => 'H',
            sr => \N__28896\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20024\,
            in1 => \N__19870\,
            in2 => \N__19449\,
            in3 => \N__20512\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_1_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__19445\,
            in1 => \N__19881\,
            in2 => \N__20608\,
            in3 => \N__20513\,
            lcout => \this_vga_signals.N_826_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__19666\,
            in1 => \N__19794\,
            in2 => \_gnd_net_\,
            in3 => \N__39882\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.G_406_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19665\,
            in1 => \N__19793\,
            in2 => \_gnd_net_\,
            in3 => \N__39881\,
            lcout => \this_vga_signals.GZ0Z_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_0_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35608\,
            in2 => \_gnd_net_\,
            in3 => \N__22162\,
            lcout => \M_this_map_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_3_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39517\,
            in2 => \_gnd_net_\,
            in3 => \N__22135\,
            lcout => \M_this_map_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_4_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41039\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22173\,
            lcout => \M_this_map_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI8K9F5_0_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29225\,
            lcout => dma_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__19450\,
            in1 => \N__19892\,
            in2 => \N__20552\,
            in3 => \N__20514\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_827_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010011001100"
        )
    port map (
            in0 => \N__19893\,
            in1 => \N__20607\,
            in2 => \N__19417\,
            in3 => \N__19987\,
            lcout => \this_vga_signals_M_lcounter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_1_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100011111000"
        )
    port map (
            in0 => \N__19414\,
            in1 => \N__19955\,
            in2 => \N__20554\,
            in3 => \N__19891\,
            lcout => \this_vga_signals_M_lcounter_q_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40345\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19795\,
            lcout => \this_pixel_clk_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40358\,
            ce => 'H',
            sr => \N__39784\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_1_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35504\,
            in2 => \_gnd_net_\,
            in3 => \N__22161\,
            lcout => \M_this_map_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_2_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38764\,
            lcout => \M_this_map_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_7_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22165\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36478\,
            lcout => \M_this_map_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_5_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__22164\,
            in1 => \N__40608\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_map_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIAJH46_5_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__21529\,
            in1 => \N__24174\,
            in2 => \N__31642\,
            in3 => \N__21646\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIITCPC_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__19720\,
            in1 => \N__23954\,
            in2 => \N__29224\,
            in3 => \N__29982\,
            lcout => \this_ppu.M_last_q_RNIITCPC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_0_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__24085\,
            in1 => \N__29148\,
            in2 => \N__31843\,
            in3 => \N__24031\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40312\,
            ce => 'H',
            sr => \N__29756\
        );

    \this_ppu.line_clk.M_last_q_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20606\,
            in1 => \N__20581\,
            in2 => \N__20553\,
            in3 => \N__20518\,
            lcout => \this_ppu.M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_srsts_0_i_o2_1_0_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20602\,
            in1 => \N__20580\,
            in2 => \N__20551\,
            in3 => \N__20511\,
            lcout => \this_ppu.N_5_4\,
            ltout => \this_ppu.N_5_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__24066\,
            in1 => \_gnd_net_\,
            in2 => \N__20404\,
            in3 => \N__29141\,
            lcout => \this_ppu.N_228_0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_0_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20401\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20383\,
            in1 => \N__34923\,
            in2 => \_gnd_net_\,
            in3 => \N__20377\,
            lcout => \M_this_ppu_spr_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_1_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__31862\,
            in1 => \N__31790\,
            in2 => \_gnd_net_\,
            in3 => \N__29968\,
            lcout => \this_ppu.M_vaddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40410\,
            ce => 'H',
            sr => \N__29769\
        );

    \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38914\,
            in1 => \N__20137\,
            in2 => \_gnd_net_\,
            in3 => \N__20122\,
            lcout => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIQER3C_9_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__29640\,
            in1 => \N__24769\,
            in2 => \_gnd_net_\,
            in3 => \N__29560\,
            lcout => \M_state_q_RNIQER3C_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNI1IH46_4_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__24172\,
            in1 => \N__21527\,
            in2 => \N__31687\,
            in3 => \N__21853\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIBKH46_6_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__21528\,
            in2 => \N__31594\,
            in3 => \N__21991\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNI0B6K1_3_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__28277\,
            in1 => \N__31734\,
            in2 => \_gnd_net_\,
            in3 => \N__24171\,
            lcout => \this_ppu.N_806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIF0FG4_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28278\,
            in1 => \N__24178\,
            in2 => \N__31738\,
            in3 => \N__21556\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38901\,
            in1 => \N__21499\,
            in2 => \_gnd_net_\,
            in3 => \N__21484\,
            lcout => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21715\,
            in1 => \N__21469\,
            in2 => \_gnd_net_\,
            in3 => \N__34975\,
            lcout => \M_this_ppu_spr_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27985\,
            in1 => \N__21256\,
            in2 => \_gnd_net_\,
            in3 => \N__34956\,
            lcout => \M_this_ppu_spr_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20614\,
            in1 => \N__21049\,
            in2 => \_gnd_net_\,
            in3 => \N__34957\,
            lcout => \M_this_ppu_spr_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29692\,
            in1 => \N__20857\,
            in2 => \_gnd_net_\,
            in3 => \N__34958\,
            lcout => \M_this_ppu_spr_addr_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_3_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20629\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_2_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21730\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_ram_write_data_0_a2_6_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36278\,
            in2 => \_gnd_net_\,
            in3 => \N__22166\,
            lcout => \M_this_map_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__22262\,
            in1 => \N__21598\,
            in2 => \N__22327\,
            in3 => \N__21697\,
            lcout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_1_RNISI5G_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21691\,
            in1 => \N__21670\,
            in2 => \_gnd_net_\,
            in3 => \N__38935\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_3_1_RNISI5GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__22264\,
            in1 => \N__38980\,
            in2 => \N__21655\,
            in3 => \N__21652\,
            lcout => \M_this_spr_ram_read_data_2\,
            ltout => \M_this_spr_ram_read_data_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vram_en_0_i_o2_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21990\,
            in1 => \N__21849\,
            in2 => \N__21637\,
            in3 => \N__21555\,
            lcout => \this_ppu.N_772_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38934\,
            in1 => \N__21634\,
            in2 => \_gnd_net_\,
            in3 => \N__21616\,
            lcout => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21592\,
            in1 => \N__21574\,
            in2 => \_gnd_net_\,
            in3 => \N__38943\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100100110001"
        )
    port map (
            in0 => \N__22263\,
            in1 => \N__21748\,
            in2 => \N__21559\,
            in3 => \N__38812\,
            lcout => \M_this_spr_ram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38944\,
            in1 => \N__21826\,
            in2 => \_gnd_net_\,
            in3 => \N__21808\,
            lcout => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38933\,
            in1 => \N__21793\,
            in2 => \_gnd_net_\,
            in3 => \N__21775\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__22323\,
            in1 => \N__22247\,
            in2 => \N__21757\,
            in3 => \N__21754\,
            lcout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_3_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__28275\,
            in1 => \N__28380\,
            in2 => \_gnd_net_\,
            in3 => \N__21909\,
            lcout => \M_this_ppu_vram_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40305\,
            ce => 'H',
            sr => \N__22414\
        );

    \this_delay_clk.M_pipe_q_2_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21742\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_1_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__24602\,
            in1 => \N__24698\,
            in2 => \N__25018\,
            in3 => \N__24655\,
            lcout => \M_this_oam_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40346\,
            ce => 'H',
            sr => \N__28895\
        );

    \this_ppu.M_state_q_8_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__24133\,
            in1 => \N__24757\,
            in2 => \N__28552\,
            in3 => \N__29580\,
            lcout => \this_ppu.M_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40359\,
            ce => 'H',
            sr => \N__39777\
        );

    \M_this_oam_address_q_RNI24IA1_1_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__24701\,
            in1 => \N__24657\,
            in2 => \N__24603\,
            in3 => \N__39883\,
            lcout => \N_1286_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_0_1_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__24702\,
            in1 => \N__24658\,
            in2 => \N__24604\,
            in3 => \N__39891\,
            lcout => \N_1294_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__21859\,
            in1 => \N__36127\,
            in2 => \N__22261\,
            in3 => \N__22030\,
            lcout => \M_this_spr_ram_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI1O64C_1_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27938\,
            in1 => \N__29330\,
            in2 => \N__28356\,
            in3 => \N__21928\,
            lcout => \this_ppu.un1_M_haddress_q_c3\,
            ltout => \this_ppu.un1_M_haddress_q_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIHAI4C_5_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28194\,
            in1 => \N__28117\,
            in2 => \N__21838\,
            in3 => \N__28285\,
            lcout => \this_ppu.un1_M_haddress_q_c6\,
            ltout => \this_ppu.un1_M_haddress_q_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_6_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21835\,
            in3 => \N__28067\,
            lcout => \M_this_ppu_vram_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40291\,
            ce => 'H',
            sr => \N__22409\
        );

    \this_ppu.M_state_q_RNIQER3C_0_9_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__29632\,
            in1 => \N__24765\,
            in2 => \_gnd_net_\,
            in3 => \N__29556\,
            lcout => \this_ppu.N_754_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_5_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__28195\,
            in1 => \N__28118\,
            in2 => \N__28295\,
            in3 => \N__21832\,
            lcout => \M_this_ppu_vram_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40291\,
            ce => 'H',
            sr => \N__22409\
        );

    \this_ppu.M_haddress_q_RNIJU24C_1_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__27942\,
            in1 => \N__29319\,
            in2 => \_gnd_net_\,
            in3 => \N__21929\,
            lcout => \this_ppu.un1_M_haddress_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__29139\,
            in1 => \N__24038\,
            in2 => \N__24099\,
            in3 => \N__39894\,
            lcout => \this_ppu.M_last_q_RNIGL6V4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_4_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__28276\,
            in1 => \N__28347\,
            in2 => \N__28196\,
            in3 => \N__21910\,
            lcout => \M_this_ppu_vram_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40300\,
            ce => 'H',
            sr => \N__22405\
        );

    \M_this_oam_address_q_0_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25006\,
            in1 => \N__24582\,
            in2 => \_gnd_net_\,
            in3 => \N__24643\,
            lcout => \M_this_oam_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40314\,
            ce => 'H',
            sr => \N__28897\
        );

    \this_ppu.M_state_q_9_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21898\,
            lcout => \this_ppu.M_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40347\,
            ce => 'H',
            sr => \N__39774\
        );

    \M_this_data_tmp_q_esr_13_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__40600\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40372\,
            ce => \N__29039\,
            sr => \N__39781\
        );

    \this_ppu.M_state_q_0_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__29115\,
            in1 => \N__23115\,
            in2 => \N__24103\,
            in3 => \N__24043\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40380\,
            ce => 'H',
            sr => \N__39785\
        );

    \this_ppu.M_count_q_7_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__23114\,
            in1 => \N__22504\,
            in2 => \_gnd_net_\,
            in3 => \N__30010\,
            lcout => \this_ppu.M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40380\,
            ce => 'H',
            sr => \N__39785\
        );

    \this_ppu.M_state_q_RNINUC91_4_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29448\,
            in2 => \_gnd_net_\,
            in3 => \N__29670\,
            lcout => \this_ppu.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_10_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40401\,
            ce => \N__29046\,
            sr => \N__39793\
        );

    \M_this_data_tmp_q_esr_12_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41054\,
            lcout => \M_this_data_tmp_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40411\,
            ce => \N__29057\,
            sr => \N__39794\
        );

    \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38932\,
            in1 => \N__21892\,
            in2 => \_gnd_net_\,
            in3 => \N__21877\,
            lcout => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38931\,
            in1 => \N__22066\,
            in2 => \_gnd_net_\,
            in3 => \N__22051\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__22318\,
            in1 => \N__22233\,
            in2 => \N__22033\,
            in3 => \N__21943\,
            lcout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_4_0_wclke_3_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__37549\,
            in1 => \N__37374\,
            in2 => \N__37477\,
            in3 => \N__37300\,
            lcout => \this_spr_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNITCNI1_12_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__22234\,
            in1 => \N__22000\,
            in2 => \N__22567\,
            in3 => \N__22319\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNINL8S2_11_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__22254\,
            in1 => \N__22525\,
            in2 => \N__21994\,
            in3 => \N__33550\,
            lcout => \M_this_spr_ram_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38930\,
            in1 => \N__21973\,
            in2 => \_gnd_net_\,
            in3 => \N__21958\,
            lcout => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_7_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__28032\,
            in1 => \N__28066\,
            in2 => \_gnd_net_\,
            in3 => \N__21937\,
            lcout => \this_ppu.M_haddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40290\,
            ce => 'H',
            sr => \N__22413\
        );

    \this_ppu.M_haddress_q_2_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001110011001100"
        )
    port map (
            in0 => \N__21931\,
            in1 => \N__28375\,
            in2 => \N__29338\,
            in3 => \N__27944\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40290\,
            ce => 'H',
            sr => \N__22413\
        );

    \this_ppu.M_haddress_q_1_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__27943\,
            in1 => \N__29323\,
            in2 => \_gnd_net_\,
            in3 => \N__21930\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40290\,
            ce => 'H',
            sr => \N__22413\
        );

    \this_ppu.M_haddress_q_0_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000011110"
        )
    port map (
            in0 => \N__29641\,
            in1 => \N__24764\,
            in2 => \N__29337\,
            in3 => \N__29579\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40290\,
            ce => 'H',
            sr => \N__22413\
        );

    \this_spr_ram.mem_mem_3_0_wclke_3_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__37358\,
            in1 => \N__37304\,
            in2 => \N__37462\,
            in3 => \N__37529\,
            lcout => \this_spr_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_12_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28969\,
            in1 => \N__22348\,
            in2 => \_gnd_net_\,
            in3 => \N__34976\,
            lcout => \this_spr_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40295\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22291\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_11_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22282\,
            in1 => \N__22975\,
            in2 => \_gnd_net_\,
            in3 => \N__34962\,
            lcout => \this_spr_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_1_i_0_0_a2_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__24454\,
            in1 => \N__36739\,
            in2 => \N__24487\,
            in3 => \N__24530\,
            lcout => \M_this_state_d_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__23026\,
            in1 => \N__24903\,
            in2 => \_gnd_net_\,
            in3 => \N__23046\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40326\,
            ce => \N__24815\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__24909\,
            in1 => \N__23809\,
            in2 => \N__39922\,
            in3 => \N__22827\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40335\,
            ce => \N__24823\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_6_11_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23047\,
            in2 => \_gnd_net_\,
            in3 => \N__23069\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100101"
        )
    port map (
            in0 => \N__23796\,
            in1 => \_gnd_net_\,
            in2 => \N__23782\,
            in3 => \N__24904\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40335\,
            ce => \N__24823\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_7_11_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23219\,
            in1 => \N__23795\,
            in2 => \N__24937\,
            in3 => \N__23820\,
            lcout => OPEN,
            ltout => \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_11_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23101\,
            in1 => \N__23128\,
            in2 => \N__22429\,
            in3 => \N__22426\,
            lcout => \this_ppu.N_934\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__23220\,
            in1 => \_gnd_net_\,
            in2 => \N__24910\,
            in3 => \N__23206\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40335\,
            ce => \N__24823\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__23056\,
            in1 => \N__24908\,
            in2 => \_gnd_net_\,
            in3 => \N__23070\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40335\,
            ce => \N__24823\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_6_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28545\,
            in2 => \_gnd_net_\,
            in3 => \N__24126\,
            lcout => \this_ppu.M_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40344\,
            ce => 'H',
            sr => \N__39775\
        );

    \M_this_data_tmp_q_esr_20_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41055\,
            lcout => \M_this_data_tmp_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40357\,
            ce => \N__32422\,
            sr => \N__39778\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25039\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23874\,
            in2 => \N__23768\,
            in3 => \N__22420\,
            lcout => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23759\,
            in2 => \N__22489\,
            in3 => \N__22417\,
            lcout => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22617\,
            in2 => \N__23769\,
            in3 => \N__22519\,
            lcout => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23763\,
            in2 => \N__22452\,
            in3 => \N__22516\,
            lcout => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23991\,
            in2 => \N__23770\,
            in3 => \N__22513\,
            lcout => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23767\,
            in2 => \N__22645\,
            in3 => \N__22510\,
            lcout => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_7_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110110"
        )
    port map (
            in0 => \N__29449\,
            in1 => \N__23857\,
            in2 => \N__30022\,
            in3 => \N__22507\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_2_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__22488\,
            in1 => \N__25093\,
            in2 => \N__22498\,
            in3 => \N__25063\,
            lcout => \this_ppu.M_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIDE0G_2_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23990\,
            in1 => \N__22445\,
            in2 => \N__22644\,
            in3 => \N__22484\,
            lcout => OPEN,
            ltout => \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIKM001_1_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22613\,
            in1 => \N__23873\,
            in2 => \N__22468\,
            in3 => \N__23842\,
            lcout => \this_ppu.M_hoffset_d_0_sqmuxa_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_4_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__22453\,
            in1 => \N__25094\,
            in2 => \N__22465\,
            in3 => \N__25065\,
            lcout => \this_ppu.M_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_6_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__25066\,
            in1 => \N__25096\,
            in2 => \N__22654\,
            in3 => \N__22640\,
            lcout => \this_ppu.M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_3_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000010"
        )
    port map (
            in0 => \N__25064\,
            in1 => \N__25095\,
            in2 => \N__22618\,
            in3 => \N__22624\,
            lcout => \this_ppu.M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_16_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35588\,
            lcout => \M_this_data_tmp_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40390\,
            ce => \N__32423\,
            sr => \N__39790\
        );

    \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39889\,
            lcout => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38936\,
            in1 => \N__22591\,
            in2 => \_gnd_net_\,
            in3 => \N__22579\,
            lcout => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_9_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__24234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22558\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_8_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__24187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24233\,
            lcout => \this_reset_cond.M_stage_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40287\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22552\,
            in1 => \N__22540\,
            in2 => \_gnd_net_\,
            in3 => \N__38937\,
            lcout => \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24255\,
            in2 => \_gnd_net_\,
            in3 => \N__22792\,
            lcout => \this_reset_cond.M_stage_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_6_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24258\,
            in2 => \_gnd_net_\,
            in3 => \N__22810\,
            lcout => \this_reset_cond.M_stage_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_5_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__24257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22798\,
            lcout => \this_reset_cond.M_stage_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_4_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24256\,
            in2 => \_gnd_net_\,
            in3 => \N__22804\,
            lcout => \this_reset_cond.M_stage_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__24260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22786\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22780\,
            in2 => \_gnd_net_\,
            in3 => \N__24259\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22774\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_wclke_3_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__37341\,
            in1 => \N__37273\,
            in2 => \N__37441\,
            in3 => \N__37500\,
            lcout => \this_spr_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__38791\,
            in1 => \N__37193\,
            in2 => \N__36294\,
            in3 => \N__36657\,
            lcout => \M_this_spr_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_5_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22993\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__24531\,
            in1 => \N__24449\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__35511\,
            in1 => \N__37183\,
            in2 => \N__40609\,
            in3 => \N__36678\,
            lcout => \M_this_spr_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_10_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24477\,
            in1 => \N__24511\,
            in2 => \_gnd_net_\,
            in3 => \N__24450\,
            lcout => \this_ppu.N_321_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_map_address_q_0_i_o2_0_a2_4_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40803\,
            lcout => \N_609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__23017\,
            in1 => \N__24900\,
            in2 => \_gnd_net_\,
            in3 => \N__23147\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40328\,
            ce => \N__24819\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__24901\,
            in1 => \N__23008\,
            in2 => \_gnd_net_\,
            in3 => \N__23193\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40328\,
            ce => \N__24819\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__23833\,
            in1 => \N__24902\,
            in2 => \_gnd_net_\,
            in3 => \N__23168\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40328\,
            ce => \N__24819\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__23091\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24899\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40328\,
            ce => \N__24819\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_9_11_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24387\,
            in1 => \N__24410\,
            in2 => \N__24357\,
            in3 => \N__23090\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_c_0_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23092\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_0_THRU_LUT4_0_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24411\,
            in2 => \N__23694\,
            in3 => \N__23077\,
            lcout => \M_this_data_count_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_1_THRU_LUT4_0_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23640\,
            in2 => \N__23074\,
            in3 => \N__23050\,
            lcout => \M_this_data_count_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_2_THRU_LUT4_0_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23045\,
            in2 => \N__23695\,
            in3 => \N__23020\,
            lcout => \M_this_data_count_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_3_THRU_LUT4_0_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23644\,
            in2 => \N__23152\,
            in3 => \N__23011\,
            lcout => \M_this_data_count_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_4_THRU_LUT4_0_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23192\,
            in2 => \N__23696\,
            in3 => \N__23002\,
            lcout => \M_this_data_count_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_5_THRU_LUT4_0_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23648\,
            in2 => \N__24388\,
            in3 => \N__22999\,
            lcout => \M_this_data_count_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_6_THRU_LUT4_0_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23697\,
            in2 => \N__24358\,
            in3 => \N__22996\,
            lcout => \M_this_data_count_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_8_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24835\,
            in2 => \N__23755\,
            in3 => \N__23836\,
            lcout => \M_this_data_count_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_8_THRU_LUT4_0_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23172\,
            in2 => \N__23749\,
            in3 => \N__23824\,
            lcout => \M_this_data_count_q_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_10_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23821\,
            in2 => \N__23754\,
            in3 => \N__23803\,
            lcout => \M_this_data_count_q_s_10\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_10_THRU_LUT4_0_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23735\,
            in2 => \N__23800\,
            in3 => \N__23773\,
            lcout => \M_this_data_count_q_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_11_THRU_LUT4_0_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23708\,
            in2 => \N__23224\,
            in3 => \N__23200\,
            lcout => \M_this_data_count_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_13_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__24933\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23197\,
            lcout => \M_this_data_count_q_s_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_8_11_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24834\,
            in1 => \N__23194\,
            in2 => \N__23173\,
            in3 => \N__23148\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_5_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__28511\,
            in1 => \N__23122\,
            in2 => \N__29455\,
            in3 => \N__29734\,
            lcout => \this_ppu.M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40360\,
            ce => 'H',
            sr => \N__39772\
        );

    \this_ppu.M_state_q_RNIEOOI_9_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29625\,
            in2 => \_gnd_net_\,
            in3 => \N__24729\,
            lcout => \this_ppu.N_760_0\,
            ltout => \this_ppu.N_760_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIKDTE1_5_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24124\,
            in1 => \N__29520\,
            in2 => \N__24181\,
            in3 => \N__41436\,
            lcout => \this_ppu.N_762_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNII6H51_5_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24730\,
            in1 => \N__24125\,
            in2 => \N__29447\,
            in3 => \N__28507\,
            lcout => \this_ppu.M_state_q_inv_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI7O615_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__24098\,
            in1 => \N__29443\,
            in2 => \N__29140\,
            in3 => \N__24039\,
            lcout => \this_ppu.N_268_i_0_0\,
            ltout => \this_ppu.N_268_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_5_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__23992\,
            in1 => \N__24001\,
            in2 => \N__23995\,
            in3 => \N__25062\,
            lcout => \this_ppu.M_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI7KJ86_0_4_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__29674\,
            in1 => \N__23953\,
            in2 => \N__29451\,
            in3 => \N__29983\,
            lcout => \this_ppu.N_1323_0\,
            ltout => \this_ppu.N_1323_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_1_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010010000"
        )
    port map (
            in0 => \N__23887\,
            in1 => \N__23875\,
            in2 => \N__23878\,
            in3 => \N__25092\,
            lcout => \this_ppu.M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40381\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIL508_7_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23856\,
            in2 => \_gnd_net_\,
            in3 => \N__25034\,
            lcout => \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_6_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24317\,
            in1 => \N__25011\,
            in2 => \_gnd_net_\,
            in3 => \N__25107\,
            lcout => \M_this_oam_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40392\,
            ce => 'H',
            sr => \N__28891\
        );

    \M_this_oam_address_q_7_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__24318\,
            in1 => \N__25013\,
            in2 => \N__24285\,
            in3 => \N__25108\,
            lcout => \M_this_oam_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40402\,
            ce => 'H',
            sr => \N__28890\
        );

    \M_this_oam_address_q_2_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25012\,
            in1 => \N__25295\,
            in2 => \_gnd_net_\,
            in3 => \N__25227\,
            lcout => \M_this_oam_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40402\,
            ce => 'H',
            sr => \N__28890\
        );

    \M_this_data_tmp_q_esr_9_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35491\,
            lcout => \M_this_data_tmp_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40412\,
            ce => \N__29053\,
            sr => \N__39791\
        );

    \M_this_data_tmp_q_esr_18_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38780\,
            lcout => \M_this_data_tmp_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40426\,
            ce => \N__32427\,
            sr => \N__39795\
        );

    \this_reset_cond.M_stage_q_7_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__24262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24193\,
            lcout => \this_reset_cond.M_stage_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_13_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32183\,
            in2 => \_gnd_net_\,
            in3 => \N__30634\,
            lcout => \this_ppu.N_324_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_9_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__40805\,
            in1 => \N__28950\,
            in2 => \_gnd_net_\,
            in3 => \N__39913\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_7_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30547\,
            in2 => \_gnd_net_\,
            in3 => \N__40804\,
            lcout => \N_332_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_en_1_sqmuxa_0_a2_i_o2_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__36799\,
            in1 => \N__24475\,
            in2 => \N__24541\,
            in3 => \N__24442\,
            lcout => \N_314_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.N_660_i_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__24476\,
            in1 => \N__30625\,
            in2 => \_gnd_net_\,
            in3 => \N__39897\,
            lcout => \N_660_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_address_q_0_i_o3_0_a2_0_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40819\,
            lcout => \N_611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_8_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__30329\,
            in1 => \N__32136\,
            in2 => \N__32275\,
            in3 => \N__28948\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__24540\,
            in1 => \N__24474\,
            in2 => \_gnd_net_\,
            in3 => \N__24441\,
            lcout => \N_309_0\,
            ltout => \N_309_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28947\,
            in2 => \N__24421\,
            in3 => \N__36656\,
            lcout => \N_260_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_data_count_qlde_0_i_i_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__40794\,
            in1 => \N__30664\,
            in2 => \N__40664\,
            in3 => \N__39890\,
            lcout => \N_257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_a2_1_0_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__28949\,
            in1 => \N__36677\,
            in2 => \_gnd_net_\,
            in3 => \N__40793\,
            lcout => \this_ppu.N_545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__24418\,
            in1 => \N__24873\,
            in2 => \_gnd_net_\,
            in3 => \N__24412\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40337\,
            ce => \N__24811\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__24394\,
            in1 => \N__24874\,
            in2 => \_gnd_net_\,
            in3 => \N__24386\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40337\,
            ce => \N__24811\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__24875\,
            in1 => \N__24364\,
            in2 => \_gnd_net_\,
            in3 => \N__24356\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40337\,
            ce => \N__24811\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__24876\,
            in1 => \N__30450\,
            in2 => \N__24949\,
            in3 => \N__39914\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40337\,
            ce => \N__24811\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a2_0_a2_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24645\,
            in1 => \N__24571\,
            in2 => \_gnd_net_\,
            in3 => \N__24700\,
            lcout => \M_this_oam_ram_write_data_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNIMU531_1_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24644\,
            in1 => \N__24699\,
            in2 => \N__36811\,
            in3 => \N__40836\,
            lcout => \un1_M_this_oam_address_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__24916\,
            in1 => \N__24898\,
            in2 => \N__25014\,
            in3 => \N__39915\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40361\,
            ce => \N__24804\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_7_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28515\,
            in2 => \_gnd_net_\,
            in3 => \N__29730\,
            lcout => \this_ppu.M_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40373\,
            ce => 'H',
            sr => \N__39767\
        );

    \this_ppu.M_oamcurr_q_3_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__30168\,
            in1 => \N__28437\,
            in2 => \_gnd_net_\,
            in3 => \N__28806\,
            lcout => \M_this_ppu_oam_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40382\,
            ce => 'H',
            sr => \N__28893\
        );

    \this_ppu.M_oamcurr_q_RNIRKBD7_4_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30164\,
            in1 => \N__25366\,
            in2 => \_gnd_net_\,
            in3 => \N__28804\,
            lcout => \this_ppu.un1_M_oamcurr_q_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIRE716_4_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29450\,
            in1 => \N__29683\,
            in2 => \_gnd_net_\,
            in3 => \N__30000\,
            lcout => \this_ppu.M_oamcurr_qc_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_1_1_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__24706\,
            in1 => \N__24656\,
            in2 => \N__24595\,
            in3 => \N__39896\,
            lcout => \N_1302_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_0_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__25038\,
            in1 => \N__25091\,
            in2 => \_gnd_net_\,
            in3 => \N__25061\,
            lcout => \this_ppu.M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_3_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__24993\,
            in1 => \N__25296\,
            in2 => \N__25254\,
            in3 => \N__25228\,
            lcout => \M_this_oam_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \this_ppu.M_oamcurr_q_1_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000001001000"
        )
    port map (
            in0 => \N__28736\,
            in1 => \N__28435\,
            in2 => \N__28674\,
            in3 => \N__28621\,
            lcout => \M_this_ppu_oam_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \M_this_oam_address_q_4_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__25203\,
            in1 => \_gnd_net_\,
            in2 => \N__25010\,
            in3 => \N__25130\,
            lcout => \M_this_oam_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \M_this_oam_address_q_5_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__25131\,
            in1 => \N__24994\,
            in2 => \N__25179\,
            in3 => \N__25204\,
            lcout => \M_this_oam_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \this_ppu.M_oamcurr_q_4_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__28436\,
            in1 => \N__25367\,
            in2 => \N__30183\,
            in3 => \N__28807\,
            lcout => \M_this_ppu_oam_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \this_ppu.M_oamcurr_q_0_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__28735\,
            in1 => \N__28432\,
            in2 => \_gnd_net_\,
            in3 => \N__28620\,
            lcout => \M_this_ppu_oam_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \this_ppu.M_oamcurr_q_5_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28434\,
            in1 => \N__28463\,
            in2 => \_gnd_net_\,
            in3 => \N__28407\,
            lcout => \M_this_ppu_oam_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \this_ppu.M_oamcurr_q_2_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28433\,
            in2 => \_gnd_net_\,
            in3 => \N__28840\,
            lcout => \M_this_ppu_oam_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40403\,
            ce => 'H',
            sr => \N__28892\
        );

    \this_ppu.M_oamcurr_q_RNI3AD1_4_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30066\,
            in1 => \N__28657\,
            in2 => \N__25377\,
            in3 => \N__28727\,
            lcout => \this_ppu.M_state_q_srsts_i_i_o2_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamidx_q_1_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__30286\,
            in1 => \N__39912\,
            in2 => \N__30259\,
            in3 => \N__30020\,
            lcout => \this_ppu.M_oamidx_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_13_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39269\,
            lcout => \M_this_oam_ram_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNILNG41_3_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25294\,
            in1 => \N__25247\,
            in2 => \_gnd_net_\,
            in3 => \N__25220\,
            lcout => \un1_M_this_oam_address_q_c4\,
            ltout => \un1_M_this_oam_address_q_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNIOKR51_5_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__25178\,
            in1 => \_gnd_net_\,
            in2 => \N__25153\,
            in3 => \N__25129\,
            lcout => \un1_M_this_oam_address_q_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_8_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35602\,
            lcout => \M_this_data_tmp_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40420\,
            ce => \N__29065\,
            sr => \N__39786\
        );

    \M_this_data_tmp_q_esr_15_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36472\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40420\,
            ce => \N__29065\,
            sr => \N__39786\
        );

    \M_this_data_tmp_q_esr_11_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39498\,
            lcout => \M_this_data_tmp_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40420\,
            ce => \N__29065\,
            sr => \N__39786\
        );

    \M_this_data_tmp_q_esr_21_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__40598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40427\,
            ce => \N__32438\,
            sr => \N__39792\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_18_LC_18_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27001\,
            in2 => \_gnd_net_\,
            in3 => \N__39270\,
            lcout => \M_this_oam_ram_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_21_LC_18_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26980\,
            in2 => \_gnd_net_\,
            in3 => \N__39271\,
            lcout => \M_this_oam_ram_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_spr_address_q_0_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30442\,
            in1 => \N__26772\,
            in2 => \N__28921\,
            in3 => \N__28920\,
            lcout => \M_this_spr_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_19_13_0_\,
            carryout => \un1_M_this_spr_address_q_cry_0\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_1_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30446\,
            in1 => \N__26576\,
            in2 => \_gnd_net_\,
            in3 => \N__26527\,
            lcout => \M_this_spr_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_0\,
            carryout => \un1_M_this_spr_address_q_cry_1\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_2_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30443\,
            in1 => \N__26340\,
            in2 => \_gnd_net_\,
            in3 => \N__26320\,
            lcout => \M_this_spr_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_1\,
            carryout => \un1_M_this_spr_address_q_cry_2\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_3_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30447\,
            in1 => \N__26090\,
            in2 => \_gnd_net_\,
            in3 => \N__26065\,
            lcout => \M_this_spr_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_2\,
            carryout => \un1_M_this_spr_address_q_cry_3\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_4_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30444\,
            in1 => \N__25889\,
            in2 => \_gnd_net_\,
            in3 => \N__25876\,
            lcout => \M_this_spr_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_3\,
            carryout => \un1_M_this_spr_address_q_cry_4\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_5_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30448\,
            in1 => \N__25687\,
            in2 => \_gnd_net_\,
            in3 => \N__25648\,
            lcout => \M_this_spr_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_4\,
            carryout => \un1_M_this_spr_address_q_cry_5\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_6_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30445\,
            in1 => \N__25407\,
            in2 => \_gnd_net_\,
            in3 => \N__25387\,
            lcout => \M_this_spr_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_5\,
            carryout => \un1_M_this_spr_address_q_cry_6\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_7_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30449\,
            in1 => \N__27695\,
            in2 => \_gnd_net_\,
            in3 => \N__27670\,
            lcout => \M_this_spr_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_6\,
            carryout => \un1_M_this_spr_address_q_cry_7\,
            clk => \N__40317\,
            ce => 'H',
            sr => \N__28900\
        );

    \M_this_spr_address_q_8_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30414\,
            in1 => \N__27484\,
            in2 => \_gnd_net_\,
            in3 => \N__27457\,
            lcout => \M_this_spr_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_19_14_0_\,
            carryout => \un1_M_this_spr_address_q_cry_8\,
            clk => \N__40322\,
            ce => 'H',
            sr => \N__28899\
        );

    \M_this_spr_address_q_9_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30417\,
            in1 => \N__27267\,
            in2 => \_gnd_net_\,
            in3 => \N__27250\,
            lcout => \M_this_spr_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_8\,
            carryout => \un1_M_this_spr_address_q_cry_9\,
            clk => \N__40322\,
            ce => 'H',
            sr => \N__28899\
        );

    \M_this_spr_address_q_10_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30412\,
            in1 => \N__27052\,
            in2 => \_gnd_net_\,
            in3 => \N__27013\,
            lcout => \M_this_spr_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_9\,
            carryout => \un1_M_this_spr_address_q_cry_10\,
            clk => \N__40322\,
            ce => 'H',
            sr => \N__28899\
        );

    \M_this_spr_address_q_11_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30416\,
            in1 => \N__37260\,
            in2 => \_gnd_net_\,
            in3 => \N__27010\,
            lcout => \M_this_spr_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_10\,
            carryout => \un1_M_this_spr_address_q_cry_11\,
            clk => \N__40322\,
            ce => 'H',
            sr => \N__28899\
        );

    \M_this_spr_address_q_12_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__30413\,
            in1 => \N__37340\,
            in2 => \_gnd_net_\,
            in3 => \N__27007\,
            lcout => \M_this_spr_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_11\,
            carryout => \un1_M_this_spr_address_q_cry_12\,
            clk => \N__40322\,
            ce => 'H',
            sr => \N__28899\
        );

    \M_this_spr_address_q_13_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__37421\,
            in1 => \N__30415\,
            in2 => \_gnd_net_\,
            in3 => \N__27004\,
            lcout => \M_this_spr_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40322\,
            ce => 'H',
            sr => \N__28899\
        );

    \M_this_state_q_RNILR691_2_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__32602\,
            in1 => \N__40827\,
            in2 => \_gnd_net_\,
            in3 => \N__39903\,
            lcout => \N_1310_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_scroll_q_esr_12_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41041\,
            lcout => \M_this_scroll_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40329\,
            ce => \N__27972\,
            sr => \N__39763\
        );

    \M_this_scroll_q_esr_15_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40338\,
            ce => \N__27973\,
            sr => \N__39760\
        );

    \M_this_scroll_q_esr_8_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35619\,
            lcout => \M_this_scroll_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40338\,
            ce => \N__27973\,
            sr => \N__39760\
        );

    \M_this_scroll_q_esr_9_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35512\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40338\,
            ce => \N__27973\,
            sr => \N__39760\
        );

    \M_this_scroll_q_esr_11_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39506\,
            lcout => \M_this_scroll_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40338\,
            ce => \N__27973\,
            sr => \N__39760\
        );

    \M_this_scroll_q_esr_14_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36269\,
            lcout => \M_this_scroll_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40338\,
            ce => \N__27973\,
            sr => \N__39760\
        );

    \M_this_scroll_q_esr_13_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40599\,
            lcout => \M_this_scroll_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40338\,
            ce => \N__27973\,
            sr => \N__39760\
        );

    \M_this_scroll_q_esr_10_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38784\,
            lcout => \M_this_scroll_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40338\,
            ce => \N__27973\,
            sr => \N__39760\
        );

    \this_ppu.un1_M_hoffset_d_cry_0_c_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29345\,
            in2 => \N__29271\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_17_0_\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_hoffset_q_esr_1_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27954\,
            in2 => \N__27910\,
            in3 => \N__27901\,
            lcout => \this_ppu.M_hoffset_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_d_cry_0\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_1\,
            clk => \N__40348\,
            ce => \N__32058\,
            sr => \N__39758\
        );

    \this_ppu.M_hoffset_q_esr_2_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28379\,
            in2 => \N__28315\,
            in3 => \N__28306\,
            lcout => \this_ppu.M_hoffset_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_d_cry_1\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_2\,
            clk => \N__40348\,
            ce => \N__32058\,
            sr => \N__39758\
        );

    \this_ppu.M_hoffset_q_esr_3_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28299\,
            in2 => \N__28225\,
            in3 => \N__28216\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_d_cry_2\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_3\,
            clk => \N__40348\,
            ce => \N__32058\,
            sr => \N__39758\
        );

    \this_ppu.M_hoffset_q_esr_4_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28206\,
            in2 => \N__28159\,
            in3 => \N__28147\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_d_cry_3\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_4\,
            clk => \N__40348\,
            ce => \N__32058\,
            sr => \N__39758\
        );

    \this_ppu.M_hoffset_q_esr_5_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28144\,
            in2 => \N__28131\,
            in3 => \N__28096\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_d_cry_4\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_5\,
            clk => \N__40348\,
            ce => \N__32058\,
            sr => \N__39758\
        );

    \this_ppu.M_hoffset_q_esr_6_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28093\,
            in2 => \N__28086\,
            in3 => \N__28039\,
            lcout => \M_this_ppu_map_addr_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_d_cry_5\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_6\,
            clk => \N__40348\,
            ce => \N__32058\,
            sr => \N__39758\
        );

    \this_ppu.M_hoffset_q_esr_7_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28036\,
            in2 => \N__28015\,
            in3 => \N__28006\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_d_cry_6\,
            carryout => \this_ppu.un1_M_hoffset_d_cry_7\,
            clk => \N__40348\,
            ce => \N__32058\,
            sr => \N__39758\
        );

    \this_ppu.M_hoffset_q_esr_8_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28003\,
            lcout => \this_ppu.M_hoffset_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40362\,
            ce => \N__32050\,
            sr => \N__39761\
        );

    \this_ppu.oam_cache.read_data_1_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28000\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamidx_q_RNIPAFC_1_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30300\,
            in2 => \_gnd_net_\,
            in3 => \N__28672\,
            lcout => OPEN,
            ltout => \this_ppu.N_61_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamidx_q_RNI8FTH1_0_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000100"
        )
    port map (
            in0 => \N__29892\,
            in1 => \N__30037\,
            in2 => \N__28555\,
            in3 => \N__28740\,
            lcout => \this_ppu.N_769_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_3_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__29847\,
            in1 => \N__33216\,
            in2 => \_gnd_net_\,
            in3 => \N__31548\,
            lcout => \this_ppu.M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40394\,
            ce => 'H',
            sr => \N__39768\
        );

    \this_ppu.M_state_q_2_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29521\,
            in2 => \_gnd_net_\,
            in3 => \N__29474\,
            lcout => \this_ppu.M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40394\,
            ce => 'H',
            sr => \N__39768\
        );

    \this_ppu.M_oamcurr_q_RNIMIF2_6_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__28528\,
            in1 => \N__28462\,
            in2 => \N__28395\,
            in3 => \N__30163\,
            lcout => \this_ppu.N_779_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIUUIB7_6_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__29729\,
            in1 => \N__41398\,
            in2 => \N__28519\,
            in3 => \N__29827\,
            lcout => \this_ppu.un1_M_state_q_2_0\,
            ltout => \this_ppu.un1_M_state_q_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamcurr_q_RNI6SKC7_2_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__28661\,
            in1 => \N__30070\,
            in2 => \N__28483\,
            in3 => \N__28728\,
            lcout => \this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamcurr_q_RNI6SKC7_0_2_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__28662\,
            in1 => \N__28729\,
            in2 => \N__30077\,
            in3 => \N__28617\,
            lcout => \this_ppu.un1_M_oamcurr_q_2_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamcurr_q_6_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__28464\,
            in1 => \N__28438\,
            in2 => \N__28396\,
            in3 => \N__28408\,
            lcout => \this_ppu.M_oamcurr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40404\,
            ce => 'H',
            sr => \N__28894\
        );

    \this_ppu.M_oamcurr_q_RNISRHKD_0_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__28764\,
            in1 => \N__28734\,
            in2 => \_gnd_net_\,
            in3 => \N__28618\,
            lcout => \this_ppu.N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI7KJ86_4_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001011"
        )
    port map (
            in0 => \N__29675\,
            in1 => \N__29415\,
            in2 => \N__39919\,
            in3 => \N__29998\,
            lcout => \this_ppu.N_329_0\,
            ltout => \this_ppu.N_329_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamcurr_q_RNIDG8LD_2_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28843\,
            in3 => \N__28839\,
            lcout => \this_ppu.N_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamcurr_q_RNI7SJLD_3_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__30178\,
            in1 => \N__28763\,
            in2 => \_gnd_net_\,
            in3 => \N__28805\,
            lcout => \this_ppu.N_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamcurr_q_RNIK5TKD_1_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000101000"
        )
    port map (
            in0 => \N__28765\,
            in1 => \N__28733\,
            in2 => \N__28673\,
            in3 => \N__28619\,
            lcout => \this_ppu.N_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIPG425_1_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__31799\,
            in1 => \N__31884\,
            in2 => \_gnd_net_\,
            in3 => \N__29999\,
            lcout => \this_ppu.un1_M_vaddress_q_c2\,
            ltout => \this_ppu.un1_M_vaddress_q_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31716\,
            in1 => \N__31669\,
            in2 => \N__28579\,
            in3 => \N__31758\,
            lcout => \this_ppu.un1_M_vaddress_q_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamidx_q_2_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__30219\,
            in1 => \N__39911\,
            in2 => \N__30244\,
            in3 => \N__30021\,
            lcout => \this_ppu.M_oamidx_qZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40421\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_8_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39328\,
            lcout => \M_this_oam_ram_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_9_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29083\,
            in2 => \_gnd_net_\,
            in3 => \N__39329\,
            lcout => \M_this_oam_ram_write_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_14_LC_19_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36293\,
            lcout => \M_this_data_tmp_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40437\,
            ce => \N__29064\,
            sr => \N__39787\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_14_LC_19_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29005\,
            in2 => \_gnd_net_\,
            in3 => \N__39368\,
            lcout => \M_this_oam_ram_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_6_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28981\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40318\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un20_i_a4_0_a3_0_a2_1_3_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30359\,
            in1 => \N__36721\,
            in2 => \N__36797\,
            in3 => \N__30502\,
            lcout => OPEN,
            ltout => \this_ppu.un20_i_a4_0_a3_0_a2_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un20_i_a4_0_a3_0_a2_3_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__36667\,
            in1 => \_gnd_net_\,
            in2 => \N__28960\,
            in3 => \N__28956\,
            lcout => dma_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_12_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__40845\,
            in1 => \N__29254\,
            in2 => \N__30367\,
            in3 => \N__28906\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40330\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_i_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__36668\,
            in1 => \N__28957\,
            in2 => \_gnd_net_\,
            in3 => \N__40844\,
            lcout => \N_260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_a2_12_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__30360\,
            in1 => \N__32314\,
            in2 => \N__36798\,
            in3 => \N__30632\,
            lcout => \this_ppu.N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_11_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__36727\,
            in1 => \N__32121\,
            in2 => \N__30334\,
            in3 => \N__30501\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_0_12_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__39893\,
            in1 => \N__32193\,
            in2 => \_gnd_net_\,
            in3 => \N__36796\,
            lcout => \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un20_i_a4_0_a3_0_a2_3_0_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30572\,
            in1 => \N__36726\,
            in2 => \N__36806\,
            in3 => \N__32262\,
            lcout => OPEN,
            ltout => \this_ppu_un20_i_a4_0_a3_0_a2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI8K9F5_1_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011001100"
        )
    port map (
            in0 => \N__30655\,
            in1 => \N__29248\,
            in2 => \N__29242\,
            in3 => \N__30508\,
            lcout => dma_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_o2_11_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40820\,
            in2 => \_gnd_net_\,
            in3 => \N__39892\,
            lcout => \this_ppu.N_328_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_1_10_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__40843\,
            in1 => \N__30499\,
            in2 => \N__32189\,
            in3 => \N__39904\,
            lcout => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_10_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30576\,
            in2 => \_gnd_net_\,
            in3 => \N__36731\,
            lcout => OPEN,
            ltout => \this_ppu.N_414_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_10_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001100"
        )
    port map (
            in0 => \N__30500\,
            in1 => \N__29158\,
            in2 => \N__29152\,
            in3 => \N__30633\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_1_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__41548\,
            in1 => \N__33223\,
            in2 => \N__29149\,
            in3 => \N__31549\,
            lcout => \this_ppu.N_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_1_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__29851\,
            in1 => \N__29362\,
            in2 => \N__41596\,
            in3 => \N__30019\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40363\,
            ce => 'H',
            sr => \N__39757\
        );

    \this_ppu.M_hoffset_q_0_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__29352\,
            in1 => \N__29820\,
            in2 => \N__29278\,
            in3 => \N__34135\,
            lcout => \this_ppu.hspr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40374\,
            ce => 'H',
            sr => \N__39759\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_0_c_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35785\,
            in2 => \N__34144\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_19_0_\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35885\,
            in2 => \N__32653\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_2_cry_0\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35325\,
            in2 => \N__34225\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_2_cry_1\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_3_c_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35020\,
            in2 => \N__33049\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_2_cry_2\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32978\,
            in2 => \N__32665\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_2_cry_3\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35178\,
            in2 => \N__32641\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_2_cry_4\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_6_c_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32860\,
            in2 => \N__32915\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_2_cry_5\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31102\,
            in2 => \N__34302\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_2_cry_6\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32677\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_20_0_\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNIH75J4_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101010001"
        )
    port map (
            in0 => \N__32689\,
            in1 => \N__31108\,
            in2 => \N__32797\,
            in3 => \N__29737\,
            lcout => \this_ppu.N_242_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIPRKS1_1_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__29813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39895\,
            lcout => \this_ppu.N_756_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_4_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29707\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_0_a2_2_6_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__36973\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37064\,
            lcout => \this_ppu.N_511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIDM8L1_1_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011110010"
        )
    port map (
            in0 => \N__29514\,
            in1 => \N__29476\,
            in2 => \N__29436\,
            in3 => \N__29682\,
            lcout => \this_ppu.N_756_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_4_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__29518\,
            in1 => \N__29633\,
            in2 => \_gnd_net_\,
            in3 => \N__29581\,
            lcout => OPEN,
            ltout => \this_ppu.N_799_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_4_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100000101"
        )
    port map (
            in0 => \N__29530\,
            in1 => \N__29519\,
            in2 => \N__29479\,
            in3 => \N__29475\,
            lcout => \this_ppu.M_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40405\,
            ce => 'H',
            sr => \N__39764\
        );

    \this_ppu.un1_oam_data_1_cry_8_c_RNI66L52_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__29843\,
            in1 => \N__33215\,
            in2 => \_gnd_net_\,
            in3 => \N__31538\,
            lcout => \this_ppu.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_voffset_q_0_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__31880\,
            in1 => \N__29821\,
            in2 => \N__33187\,
            in3 => \N__34839\,
            lcout => \this_ppu.vspr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40415\,
            ce => 'H',
            sr => \N__39769\
        );

    \this_ppu.M_vaddress_q_2_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__31807\,
            in1 => \N__31768\,
            in2 => \N__31885\,
            in3 => \N__30025\,
            lcout => \this_ppu.M_vaddress_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40422\,
            ce => 'H',
            sr => \N__29776\
        );

    \this_ppu.M_vaddress_q_3_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__31766\,
            in1 => \N__31718\,
            in2 => \_gnd_net_\,
            in3 => \N__29796\,
            lcout => \this_ppu.M_vaddress_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40422\,
            ce => 'H',
            sr => \N__29776\
        );

    \this_ppu.M_vaddress_q_4_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__29797\,
            in1 => \N__31673\,
            in2 => \N__31727\,
            in3 => \N__31767\,
            lcout => \this_ppu.M_vaddress_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40422\,
            ce => 'H',
            sr => \N__29776\
        );

    \this_ppu.M_vaddress_q_7_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__29788\,
            in1 => \N__32077\,
            in2 => \N__31632\,
            in3 => \N__31577\,
            lcout => \this_ppu.M_vaddress_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40422\,
            ce => 'H',
            sr => \N__29776\
        );

    \this_ppu.M_vaddress_q_5_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31621\,
            in2 => \_gnd_net_\,
            in3 => \N__29786\,
            lcout => \this_ppu.M_vaddress_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40422\,
            ce => 'H',
            sr => \N__29776\
        );

    \this_ppu.M_vaddress_q_6_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__29787\,
            in1 => \_gnd_net_\,
            in2 => \N__31631\,
            in3 => \N__31576\,
            lcout => \this_ppu.M_vaddress_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40422\,
            ce => 'H',
            sr => \N__29776\
        );

    \this_ppu.un1_M_oamidx_q_cry_0_c_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41437\,
            in2 => \N__29884\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_24_0_\,
            carryout => \this_ppu.un1_M_oamidx_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oamidx_q_cry_0_THRU_LUT4_0_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30299\,
            in3 => \N__30247\,
            lcout => \this_ppu.un1_M_oamidx_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oamidx_q_cry_0\,
            carryout => \this_ppu.un1_M_oamidx_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oamidx_q_cry_1_THRU_LUT4_0_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30218\,
            in2 => \_gnd_net_\,
            in3 => \N__30235\,
            lcout => \this_ppu.un1_M_oamidx_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oamidx_q_cry_1\,
            carryout => \this_ppu.un1_M_oamidx_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamidx_q_3_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__30024\,
            in1 => \N__39909\,
            in2 => \N__30120\,
            in3 => \N__30232\,
            lcout => \this_ppu.M_oamidx_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamidx_q_RNIORUO_3_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__30217\,
            in1 => \N__30182\,
            in2 => \N__30119\,
            in3 => \N__30081\,
            lcout => \this_ppu.M_state_q_srsts_0_a3_0_o2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oamidx_q_0_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__39910\,
            in1 => \N__41438\,
            in2 => \N__29885\,
            in3 => \N__30023\,
            lcout => \this_ppu.M_oamidx_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_2_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38779\,
            lcout => \M_this_data_tmp_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40438\,
            ce => \N__36015\,
            sr => \N__39779\
        );

    \M_this_data_tmp_q_esr_5_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40607\,
            lcout => \M_this_data_tmp_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40438\,
            ce => \N__36015\,
            sr => \N__39779\
        );

    \M_this_data_tmp_q_esr_19_LC_20_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39497\,
            lcout => \M_this_data_tmp_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40445\,
            ce => \N__32437\,
            sr => \N__39782\
        );

    \M_this_data_tmp_q_esr_23_LC_20_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36487\,
            lcout => \M_this_data_tmp_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40445\,
            ce => \N__32437\,
            sr => \N__39782\
        );

    \M_this_data_tmp_q_esr_17_LC_20_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40450\,
            ce => \N__32442\,
            sr => \N__39788\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_1_7_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__32266\,
            in1 => \N__30373\,
            in2 => \N__32194\,
            in3 => \N__39908\,
            lcout => OPEN,
            ltout => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__30451\,
            in1 => \N__36670\,
            in2 => \N__30376\,
            in3 => \N__32267\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_7_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__36669\,
            in1 => \N__30539\,
            in2 => \_gnd_net_\,
            in3 => \N__30626\,
            lcout => \this_ppu.N_405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un20_i_a4_0_a2_0_a2_0_2_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__36775\,
            in1 => \N__30364\,
            in2 => \_gnd_net_\,
            in3 => \N__32260\,
            lcout => this_ppu_un20_i_a4_0_a2_0_a2_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__33790\,
            in1 => \N__32111\,
            in2 => \N__32346\,
            in3 => \N__30543\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_data_count_qlde_0_i_o2_0_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__30366\,
            in1 => \N__32261\,
            in2 => \_gnd_net_\,
            in3 => \N__30498\,
            lcout => \this_ppu.N_341_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_i_0_1_13_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001010"
        )
    port map (
            in0 => \N__30365\,
            in1 => \N__40847\,
            in2 => \N__39921\,
            in3 => \N__36776\,
            lcout => OPEN,
            ltout => \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_13_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__36777\,
            in1 => \_gnd_net_\,
            in2 => \N__30337\,
            in3 => \N__30330\,
            lcout => \M_this_state_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_0_a2_5_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__30571\,
            in1 => \_gnd_net_\,
            in2 => \N__32122\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_ppu.N_424_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__36985\,
            in1 => \N__37078\,
            in2 => \N__30667\,
            in3 => \N__33789\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_data_count_qlde_0_i_a2_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__30645\,
            in1 => \N__32185\,
            in2 => \_gnd_net_\,
            in3 => \N__30627\,
            lcout => \this_ppu.N_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI1G0L_1_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__36508\,
            in1 => \N__36683\,
            in2 => \_gnd_net_\,
            in3 => \N__32626\,
            lcout => \M_this_state_q_RNI1G0LZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_i_1_0_0_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010001"
        )
    port map (
            in0 => \N__32107\,
            in1 => \N__32563\,
            in2 => \N__30649\,
            in3 => \N__30628\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_i_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un20_i_a4_0_a2_0_o2_2_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32301\,
            in1 => \N__30570\,
            in2 => \_gnd_net_\,
            in3 => \N__30538\,
            lcout => \N_311_0\,
            ltout => \N_311_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI244K2_10_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__32227\,
            in1 => \N__30517\,
            in2 => \N__30511\,
            in3 => \N__30466\,
            lcout => \M_this_state_q_RNI244K2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIR71E_10_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36722\,
            in2 => \_gnd_net_\,
            in3 => \N__30494\,
            lcout => \M_this_state_q_RNIR71EZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.hspr_cry_0_c_inv_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35784\,
            in1 => \N__34134\,
            in2 => \N__30460\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.hspr_cry_0_c_inv_RNI1203\,
            ltout => OPEN,
            carryin => \bfn_21_17_0_\,
            carryout => \this_ppu.hspr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.hspr_cry_0_c_RNISEIH1_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100110011100"
        )
    port map (
            in0 => \N__34966\,
            in1 => \N__35886\,
            in2 => \N__30676\,
            in3 => \N__30895\,
            lcout => \M_this_ppu_spr_addr_1\,
            ltout => OPEN,
            carryin => \this_ppu.hspr_cry_0\,
            carryout => \this_ppu.hspr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.hspr_cry_1_c_RNI6K8I1_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011001001"
        )
    port map (
            in0 => \N__34967\,
            in1 => \N__35324\,
            in2 => \N__36586\,
            in3 => \N__30892\,
            lcout => \M_this_ppu_spr_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNIUU07_9_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35848\,
            lcout => \this_ppu.M_oam_cache_read_data_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_0_c_inv_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35782\,
            in2 => \N__32538\,
            in3 => \N__34124\,
            lcout => \this_ppu.M_hoffset_q_i_0\,
            ltout => OPEN,
            carryin => \bfn_21_18_0_\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_1_c_inv_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35846\,
            in2 => \N__32520\,
            in3 => \N__35887\,
            lcout => \this_ppu.M_hoffset_q_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_2_cry_0\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_2_c_inv_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36582\,
            in2 => \N__32502\,
            in3 => \N__35332\,
            lcout => \this_ppu.M_hoffset_q_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_2_cry_1\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_3_c_inv_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35931\,
            in2 => \N__32481\,
            in3 => \N__33050\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_2_cry_2\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_4_c_inv_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35077\,
            in2 => \N__32463\,
            in3 => \N__32985\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_2_cry_3\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_5_c_inv_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35124\,
            in2 => \N__32739\,
            in3 => \N__35174\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_2_cry_4\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_6_c_inv_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34427\,
            in2 => \N__32721\,
            in3 => \N__32902\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_2_cry_5\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_7_c_inv_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32703\,
            in2 => \N__34368\,
            in3 => \N__34286\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_2_cry_6\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_2_cry_8_c_inv_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31117\,
            in2 => \_gnd_net_\,
            in3 => \N__32822\,
            lcout => \this_ppu.M_hoffset_q_i_8\,
            ltout => OPEN,
            carryin => \bfn_21_19_0_\,
            carryout => \this_ppu.un1_M_hoffset_q_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_2_cry_8_c_RNITUI32_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__34367\,
            in1 => \N__34393\,
            in2 => \_gnd_net_\,
            in3 => \N__31111\,
            lcout => \this_ppu.vspr12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNO_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__34366\,
            in1 => \N__34392\,
            in2 => \_gnd_net_\,
            in3 => \N__34296\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_0_c_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39061\,
            in2 => \N__34857\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_20_0_\,
            carryout => \this_ppu.un1_oam_data_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_1_c_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39010\,
            in2 => \N__33106\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_0\,
            carryout => \this_ppu.un1_oam_data_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_2_c_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38389\,
            in2 => \N__33538\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_1\,
            carryout => \this_ppu.un1_oam_data_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_3_c_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38182\,
            in2 => \N__33489\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_2\,
            carryout => \this_ppu.un1_oam_data_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_4_c_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38596\,
            in2 => \N__33438\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_3\,
            carryout => \this_ppu.un1_oam_data_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_5_c_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32746\,
            in2 => \N__33390\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_4\,
            carryout => \this_ppu.un1_oam_data_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_6_c_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32764\,
            in2 => \N__33345\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_5\,
            carryout => \this_ppu.un1_oam_data_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_7_c_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32752\,
            in2 => \N__33291\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_6\,
            carryout => \this_ppu.un1_oam_data_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_8_c_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32758\,
            in2 => \N__33250\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_21_0_\,
            carryout => \this_ppu.un1_oam_data_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_8_THRU_LUT4_0_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31552\,
            lcout => \this_ppu.un1_oam_data_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vspr_cry_0_c_inv_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34843\,
            in2 => \N__31522\,
            in3 => \N__35401\,
            lcout => \this_ppu.vspr_cry_0_c_inv_RNIFK43\,
            ltout => OPEN,
            carryin => \bfn_21_22_0_\,
            carryout => \this_ppu.vspr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vspr_cry_0_c_RNI75JG1_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100110011100"
        )
    port map (
            in0 => \N__34940\,
            in1 => \N__33102\,
            in2 => \N__31912\,
            in3 => \N__31315\,
            lcout => \M_this_ppu_spr_addr_4\,
            ltout => OPEN,
            carryin => \this_ppu.vspr_cry_0\,
            carryout => \this_ppu.vspr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vspr_cry_1_c_RNIA9KG1_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001011100001"
        )
    port map (
            in0 => \N__32770\,
            in1 => \N__34941\,
            in2 => \N__33537\,
            in3 => \N__31312\,
            lcout => \M_this_ppu_spr_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNID8M7_17_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31891\,
            lcout => \this_ppu.M_oam_cache_read_data_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_17_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31903\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40423\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_d_cry_0_c_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31876\,
            in2 => \N__33180\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_23_0_\,
            carryout => \this_ppu.un1_M_voffset_d_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_voffset_q_esr_1_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31806\,
            in2 => \N__33163\,
            in3 => \N__31771\,
            lcout => \this_ppu.M_voffset_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_d_cry_0\,
            carryout => \this_ppu.un1_M_voffset_d_cry_1\,
            clk => \N__40430\,
            ce => \N__32057\,
            sr => \N__39770\
        );

    \this_ppu.M_voffset_q_esr_2_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31757\,
            in2 => \N__33655\,
            in3 => \N__31741\,
            lcout => \this_ppu.M_voffset_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_d_cry_1\,
            carryout => \this_ppu.un1_M_voffset_d_cry_2\,
            clk => \N__40430\,
            ce => \N__32057\,
            sr => \N__39770\
        );

    \this_ppu.M_voffset_q_esr_3_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31717\,
            in2 => \N__33145\,
            in3 => \N__31690\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_d_cry_2\,
            carryout => \this_ppu.un1_M_voffset_d_cry_3\,
            clk => \N__40430\,
            ce => \N__32057\,
            sr => \N__39770\
        );

    \this_ppu.M_voffset_q_esr_4_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33136\,
            in2 => \N__31677\,
            in3 => \N__31645\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_d_cry_3\,
            carryout => \this_ppu.un1_M_voffset_d_cry_4\,
            clk => \N__40430\,
            ce => \N__32057\,
            sr => \N__39770\
        );

    \this_ppu.M_voffset_q_esr_5_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31617\,
            in2 => \N__33154\,
            in3 => \N__31597\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_d_cry_4\,
            carryout => \this_ppu.un1_M_voffset_d_cry_5\,
            clk => \N__40430\,
            ce => \N__32057\,
            sr => \N__39770\
        );

    \this_ppu.M_voffset_q_esr_6_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33130\,
            in2 => \N__31581\,
            in3 => \N__32080\,
            lcout => \M_this_ppu_map_addr_8\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_d_cry_5\,
            carryout => \this_ppu.un1_M_voffset_d_cry_6\,
            clk => \N__40430\,
            ce => \N__32057\,
            sr => \N__39770\
        );

    \this_ppu.M_voffset_q_esr_7_LC_21_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32076\,
            in2 => \N__33124\,
            in3 => \N__32065\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_d_cry_6\,
            carryout => \this_ppu.un1_M_voffset_d_cry_7\,
            clk => \N__40430\,
            ce => \N__32057\,
            sr => \N__39770\
        );

    \this_ppu.M_voffset_q_esr_8_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32062\,
            lcout => \this_ppu.M_voffset_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40439\,
            ce => \N__32059\,
            sr => \N__39773\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_2_LC_21_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32011\,
            lcout => \M_this_oam_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_16_LC_21_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39347\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31993\,
            lcout => \M_this_oam_ram_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_5_LC_21_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31966\,
            in2 => \_gnd_net_\,
            in3 => \N__39349\,
            lcout => \M_this_oam_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_15_LC_21_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31948\,
            in2 => \_gnd_net_\,
            in3 => \N__39346\,
            lcout => \M_this_oam_ram_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_19_LC_21_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39372\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31930\,
            lcout => \M_this_oam_ram_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_0_LC_21_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35563\,
            lcout => \M_this_data_tmp_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40454\,
            ce => \N__36028\,
            sr => \N__39783\
        );

    \M_this_data_tmp_q_esr_22_LC_21_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36307\,
            lcout => \M_this_data_tmp_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40460\,
            ce => \N__32446\,
            sr => \N__39789\
        );

    \this_spr_ram.mem_radreg_13_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34171\,
            in1 => \N__32365\,
            in2 => \_gnd_net_\,
            in3 => \N__34981\,
            lcout => \this_spr_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_0_i_1_6_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__39902\,
            in1 => \N__33751\,
            in2 => \N__32350\,
            in3 => \N__36885\,
            lcout => OPEN,
            ltout => \this_ppu.M_this_state_q_srsts_0_i_0_i_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__33715\,
            in1 => \N__32123\,
            in2 => \N__32317\,
            in3 => \N__32309\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_0_a2_1_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__36519\,
            in1 => \N__40846\,
            in2 => \N__36893\,
            in3 => \N__39901\,
            lcout => \this_ppu.N_416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32132\,
            in1 => \N__33778\,
            in2 => \N__32601\,
            in3 => \N__33802\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un20_i_a4_0_a3_0_a2_1_1_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32302\,
            in1 => \N__32586\,
            in2 => \N__32629\,
            in3 => \N__32268\,
            lcout => this_ppu_un20_i_a4_0_a3_0_a2_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_0_a2_3_6_LC_22_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__41269\,
            in1 => \N__32221\,
            in2 => \_gnd_net_\,
            in3 => \N__32184\,
            lcout => \this_ppu.N_916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32625\,
            in1 => \N__33796\,
            in2 => \N__32137\,
            in3 => \N__33779\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40375\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIKV6G1_2_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__39884\,
            in1 => \N__32628\,
            in2 => \N__32597\,
            in3 => \N__40848\,
            lcout => \N_1318_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_i_a2_1_0_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32627\,
            in1 => \N__32590\,
            in2 => \N__36518\,
            in3 => \N__39885\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0\,
            ltout => \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__36843\,
            in1 => \N__36886\,
            in2 => \N__32557\,
            in3 => \N__32554\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__36966\,
            in1 => \N__32548\,
            in2 => \N__37077\,
            in3 => \N__33774\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_0_c_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35783\,
            in2 => \N__32539\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_18_0_\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_1_c_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35847\,
            in2 => \N__32521\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_cry_0\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_2_c_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36581\,
            in2 => \N__32503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_cry_1\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_3_c_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35932\,
            in2 => \N__32485\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_cry_2\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_4_c_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35072\,
            in2 => \N__32464\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_cry_3\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_5_c_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35125\,
            in2 => \N__32740\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_cry_4\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_6_c_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34428\,
            in2 => \N__32722\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_cry_5\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_7_c_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32704\,
            in2 => \N__34369\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_hoffset_q_cry_6\,
            carryout => \this_ppu.un1_M_hoffset_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_hoffset_q_cry_7_c_RNIB1P42_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__34386\,
            in1 => \N__34354\,
            in2 => \_gnd_net_\,
            in3 => \N__32692\,
            lcout => \this_ppu.vspr16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_RNO_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34344\,
            in2 => \_gnd_net_\,
            in3 => \N__34385\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_ac0_13_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNO_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \N__32826\,
            in1 => \N__34343\,
            in2 => \_gnd_net_\,
            in3 => \N__34384\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNO_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__32989\,
            in1 => \N__35065\,
            in2 => \_gnd_net_\,
            in3 => \N__35229\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNO_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__35898\,
            in1 => \N__35826\,
            in2 => \_gnd_net_\,
            in3 => \N__35761\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNO_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001011111"
        )
    port map (
            in0 => \N__35230\,
            in1 => \N__35182\,
            in2 => \N__35073\,
            in3 => \N__35117\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_6_c_RNO_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001011111"
        )
    port map (
            in0 => \N__35693\,
            in1 => \_gnd_net_\,
            in2 => \N__34499\,
            in3 => \N__34558\,
            lcout => \this_ppu.un1_oam_data_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_8_c_RNO_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__34560\,
            in1 => \N__34495\,
            in2 => \N__35680\,
            in3 => \N__35695\,
            lcout => \this_ppu.un1_oam_data_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_7_c_RNO_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100110011"
        )
    port map (
            in0 => \N__35694\,
            in1 => \N__35675\,
            in2 => \N__34500\,
            in3 => \N__34559\,
            lcout => \this_ppu.un1_oam_data_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI3DGK1_14_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011100001111"
        )
    port map (
            in0 => \N__35228\,
            in1 => \N__35108\,
            in2 => \N__34429\,
            in3 => \N__35063\,
            lcout => \this_ppu.read_data_RNI3DGK1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_5_c_RNO_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34488\,
            in2 => \_gnd_net_\,
            in3 => \N__35692\,
            lcout => \this_ppu.un1_oam_data_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNO_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__35227\,
            in1 => \N__32990\,
            in2 => \_gnd_net_\,
            in3 => \N__35062\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_0_c_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35753\,
            in2 => \N__34154\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_21_0_\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35897\,
            in2 => \N__35704\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_3_cry_0\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35333\,
            in2 => \N__35275\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_3_cry_1\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_3_c_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35013\,
            in2 => \N__33063\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_3_cry_2\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33010\,
            in2 => \N__32994\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_3_cry_3\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35026\,
            in2 => \N__35199\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_3_cry_4\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_6_c_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32919\,
            in2 => \N__32856\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_3_cry_5\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34300\,
            in2 => \N__34237\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_read_data_3_cry_6\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32839\,
            in2 => \N__32830\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_22_0_\,
            carryout => \this_ppu.un1_M_oam_cache_read_data_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_LUT4_0_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32800\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_18_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32782\,
            lcout => \this_ppu.M_oam_cache_read_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_scroll_q_esr_0_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35569\,
            lcout => \M_this_scroll_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40440\,
            ce => \N__33633\,
            sr => \N__39765\
        );

    \M_this_scroll_q_esr_1_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35475\,
            lcout => \M_this_scroll_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40440\,
            ce => \N__33633\,
            sr => \N__39765\
        );

    \M_this_scroll_q_esr_5_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40574\,
            lcout => \M_this_scroll_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40440\,
            ce => \N__33633\,
            sr => \N__39765\
        );

    \M_this_scroll_q_esr_3_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39454\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40440\,
            ce => \N__33633\,
            sr => \N__39765\
        );

    \M_this_scroll_q_esr_4_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41016\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40440\,
            ce => \N__33633\,
            sr => \N__39765\
        );

    \M_this_scroll_q_esr_6_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36262\,
            lcout => \M_this_scroll_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40440\,
            ce => \N__33633\,
            sr => \N__39765\
        );

    \M_this_scroll_q_esr_7_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36462\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40440\,
            ce => \N__33633\,
            sr => \N__39765\
        );

    \this_ppu.un1_M_voffset_q_cry_0_c_inv_LC_22_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39057\,
            in2 => \N__33115\,
            in3 => \N__34850\,
            lcout => \this_ppu.M_voffset_q_i_0\,
            ltout => OPEN,
            carryin => \bfn_22_24_0_\,
            carryout => \this_ppu.un1_M_voffset_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_1_c_inv_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39103\,
            in2 => \N__33082\,
            in3 => \N__33098\,
            lcout => \this_ppu.M_voffset_q_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_q_cry_0\,
            carryout => \this_ppu.un1_M_voffset_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_2_c_inv_LC_22_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38441\,
            in2 => \N__33511\,
            in3 => \N__33527\,
            lcout => \this_ppu.M_voffset_q_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_q_cry_1\,
            carryout => \this_ppu.un1_M_voffset_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_3_c_inv_LC_22_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38565\,
            in2 => \N__33457\,
            in3 => \N__33476\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_q_cry_2\,
            carryout => \this_ppu.un1_M_voffset_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_4_c_inv_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38508\,
            in2 => \N__33406\,
            in3 => \N__33425\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_q_cry_3\,
            carryout => \this_ppu.un1_M_voffset_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_5_c_inv_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34484\,
            in2 => \N__33358\,
            in3 => \N__33377\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_7\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_q_cry_4\,
            carryout => \this_ppu.un1_M_voffset_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_6_c_inv_LC_22_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34554\,
            in2 => \N__33307\,
            in3 => \N__33326\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_8\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_q_cry_5\,
            carryout => \this_ppu.un1_M_voffset_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_7_c_inv_LC_22_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35671\,
            in2 => \N__33259\,
            in3 => \N__33278\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_9\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_voffset_q_cry_6\,
            carryout => \this_ppu.un1_M_voffset_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_8_c_inv_LC_22_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33232\,
            in2 => \_gnd_net_\,
            in3 => \N__33243\,
            lcout => \this_ppu.M_voffset_q_i_8\,
            ltout => OPEN,
            carryin => \bfn_22_25_0_\,
            carryout => \this_ppu.un1_M_voffset_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_voffset_q_cry_8_c_RNICN6N1_LC_22_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__38209\,
            in1 => \N__38044\,
            in2 => \_gnd_net_\,
            in3 => \N__33226\,
            lcout => \this_ppu.M_state_d14_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_24_LC_22_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35598\,
            in2 => \_gnd_net_\,
            in3 => \N__39333\,
            lcout => \N_433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_29_LC_22_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40575\,
            lcout => \N_438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_12_LC_22_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33673\,
            lcout => \M_this_oam_ram_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_scroll_q_esr_2_LC_22_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38765\,
            lcout => \M_this_scroll_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40455\,
            ce => \N__33640\,
            sr => \N__39776\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_0_LC_22_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33616\,
            in2 => \_gnd_net_\,
            in3 => \N__39370\,
            lcout => \M_this_oam_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_1_LC_22_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35470\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40461\,
            ce => \N__36029\,
            sr => \N__39780\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_1_LC_22_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33598\,
            lcout => \M_this_oam_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_25_LC_22_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39369\,
            lcout => \N_434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33571\,
            in1 => \N__33562\,
            in2 => \_gnd_net_\,
            in3 => \N__38900\,
            lcout => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__37373\,
            in1 => \N__37303\,
            in2 => \N__37474\,
            in3 => \N__37550\,
            lcout => \this_spr_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_7_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34186\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_hoffset_q_RNI91DA2_0_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__34977\,
            in1 => \N__34158\,
            in2 => \N__34159\,
            in3 => \N__35781\,
            lcout => \M_this_ppu_spr_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__37194\,
            in1 => \N__35623\,
            in2 => \N__41056\,
            in3 => \N__36688\,
            lcout => \M_this_spr_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_2_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__36986\,
            in1 => \N__37074\,
            in2 => \_gnd_net_\,
            in3 => \N__36830\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_3_LC_23_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36987\,
            in1 => \N__37075\,
            in2 => \_gnd_net_\,
            in3 => \N__36831\,
            lcout => \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__36829\,
            in1 => \N__41259\,
            in2 => \N__36919\,
            in3 => \N__33745\,
            lcout => \M_this_state_d_0_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_0_a2_1_1_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__36875\,
            in1 => \N__33714\,
            in2 => \N__39920\,
            in3 => \N__33746\,
            lcout => \this_ppu.N_510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_this_state_q_4_i_0_a2_0_a2_0_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__33747\,
            in1 => \N__36967\,
            in2 => \N__37076\,
            in3 => \N__33713\,
            lcout => \N_608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNIPMBQ1_16_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__34968\,
            in1 => \N__35400\,
            in2 => \_gnd_net_\,
            in3 => \N__34858\,
            lcout => \M_this_ppu_spr_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_15_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34588\,
            lcout => \this_ppu.un1_M_hoffset_q_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_14_LC_23_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34576\,
            lcout => \this_ppu.un1_M_hoffset_q_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41554\,
            in2 => \_gnd_net_\,
            in3 => \N__34564\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41553\,
            in2 => \_gnd_net_\,
            in3 => \N__34501\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI3DGK1_0_14_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35106\,
            in1 => \N__35061\,
            in2 => \N__34423\,
            in3 => \N__35226\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_c7\,
            ltout => \this_ppu.un1_M_oam_cache_read_data_c7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNO_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34342\,
            in2 => \N__34309\,
            in3 => \N__34301\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNO_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__36568\,
            in1 => \N__35832\,
            in2 => \N__35338\,
            in3 => \N__35762\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_12_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35350\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.un1_M_hoffset_q_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNO_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111111010"
        )
    port map (
            in0 => \N__35750\,
            in1 => \N__35334\,
            in2 => \N__35836\,
            in3 => \N__36562\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_9_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35266\,
            lcout => \this_ppu.un1_M_hoffset_q_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_8_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35254\,
            lcout => \this_ppu.un1_M_hoffset_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_13_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35242\,
            lcout => \this_ppu.un1_M_hoffset_q_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI80ET_0_11_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__36560\,
            in1 => \N__35820\,
            in2 => \N__35923\,
            in3 => \N__35749\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_c4\,
            ltout => \this_ppu.un1_M_oam_cache_read_data_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNO_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100110011"
        )
    port map (
            in0 => \N__35192\,
            in1 => \N__35107\,
            in2 => \N__35080\,
            in3 => \N__35064\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI80ET_11_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__36561\,
            in1 => \N__35824\,
            in2 => \N__35924\,
            in3 => \N__35751\,
            lcout => \this_ppu.read_data_RNI80ET_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35002\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_11_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35941\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.un1_M_hoffset_q_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40432\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNO_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__35899\,
            in1 => \N__35825\,
            in2 => \_gnd_net_\,
            in3 => \N__35752\,
            lcout => \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_4_c5_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010100000"
        )
    port map (
            in0 => \N__38566\,
            in1 => \N__38443\,
            in2 => \N__38512\,
            in3 => \N__38359\,
            lcout => \this_ppu.un1_oam_data_1_4_c5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41469\,
            in2 => \_gnd_net_\,
            in3 => \N__35679\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_14_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__40717\,
            in1 => \N__37984\,
            in2 => \N__36308\,
            in3 => \N__40887\,
            lcout => \M_this_ext_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40441\,
            ce => 'H',
            sr => \N__39762\
        );

    \M_this_ext_address_q_8_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__40885\,
            in1 => \N__40719\,
            in2 => \N__35618\,
            in3 => \N__37810\,
            lcout => \M_this_ext_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40441\,
            ce => 'H',
            sr => \N__39762\
        );

    \M_this_ext_address_q_9_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__40718\,
            in1 => \N__40886\,
            in2 => \N__37777\,
            in3 => \N__35498\,
            lcout => \M_this_ext_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40441\,
            ce => 'H',
            sr => \N__39762\
        );

    \this_ppu.oam_cache.read_data_16_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35413\,
            lcout => \this_ppu.M_oam_cache_read_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40446\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_20_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35380\,
            in2 => \_gnd_net_\,
            in3 => \N__39314\,
            lcout => \M_this_oam_ram_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_6_LC_23_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40451\,
            ce => \N__36030\,
            sr => \N__39766\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_7_LC_23_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36073\,
            in2 => \_gnd_net_\,
            in3 => \N__39315\,
            lcout => \M_this_oam_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_7_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36477\,
            lcout => \M_this_data_tmp_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40451\,
            ce => \N__36030\,
            sr => \N__39766\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_3_LC_23_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36055\,
            in2 => \_gnd_net_\,
            in3 => \N__39316\,
            lcout => \M_this_oam_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_3_LC_23_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39478\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40456\,
            ce => \N__36031\,
            sr => \N__39771\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_4_LC_23_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39317\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36037\,
            lcout => \M_this_oam_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_4_LC_23_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41029\,
            lcout => \M_this_data_tmp_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40456\,
            ce => \N__36031\,
            sr => \N__39771\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_23_LC_23_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35974\,
            in2 => \_gnd_net_\,
            in3 => \N__39318\,
            lcout => \M_this_oam_ram_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_23_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41584\,
            in2 => \_gnd_net_\,
            in3 => \N__39102\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_31_LC_23_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36486\,
            in2 => \_gnd_net_\,
            in3 => \N__39308\,
            lcout => \N_440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_28_LC_23_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40983\,
            in2 => \_gnd_net_\,
            in3 => \N__39307\,
            lcout => \N_437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_22_LC_23_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36331\,
            in2 => \_gnd_net_\,
            in3 => \N__39313\,
            lcout => \M_this_oam_ram_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_30_LC_23_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36313\,
            in2 => \_gnd_net_\,
            in3 => \N__39312\,
            lcout => \N_439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__37384\,
            in1 => \N__37476\,
            in2 => \N__37305\,
            in3 => \N__37555\,
            lcout => \this_spr_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__37379\,
            in1 => \N__37467\,
            in2 => \N__37306\,
            in3 => \N__37551\,
            lcout => \this_spr_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_24_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36145\,
            in1 => \N__36139\,
            in2 => \_gnd_net_\,
            in3 => \N__38899\,
            lcout => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37301\,
            in1 => \N__37375\,
            in2 => \N__37475\,
            in3 => \N__37547\,
            lcout => \this_spr_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__37548\,
            in1 => \N__37466\,
            in2 => \N__37383\,
            in3 => \N__37302\,
            lcout => \this_spr_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_24_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36429\,
            in1 => \N__37201\,
            in2 => \N__39516\,
            in3 => \N__36679\,
            lcout => \M_this_spr_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_i_0_a2_1_3_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__37063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36988\,
            lcout => \this_ppu.N_610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__36910\,
            in1 => \N__36832\,
            in2 => \N__36894\,
            in3 => \N__36844\,
            lcout => \M_this_substate_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40407\,
            ce => 'H',
            sr => \N__39754\
        );

    \this_ppu.un1_M_this_state_q_1_i_0_0_i_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__36810\,
            in1 => \N__36738\,
            in2 => \N__36687\,
            in3 => \N__40855\,
            lcout => \N_312_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_10_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36595\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.un1_M_hoffset_q_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41602\,
            in2 => \_gnd_net_\,
            in3 => \N__38442\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_15_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__40879\,
            in1 => \N__36476\,
            in2 => \N__40720\,
            in3 => \N__37945\,
            lcout => \M_this_ext_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40433\,
            ce => 'H',
            sr => \N__39755\
        );

    \M_this_ctrl_flags_q_7_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__37743\,
            in1 => \N__36523\,
            in2 => \N__36485\,
            in3 => \N__40882\,
            lcout => \M_this_ctrl_flags_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40433\,
            ce => 'H',
            sr => \N__39755\
        );

    \M_this_ext_address_q_0_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__40880\,
            in1 => \N__37700\,
            in2 => \N__40721\,
            in3 => \N__37731\,
            lcout => \M_this_ext_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40433\,
            ce => 'H',
            sr => \N__39755\
        );

    \M_this_ext_address_q_1_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__37668\,
            in1 => \N__40883\,
            in2 => \N__37651\,
            in3 => \N__40699\,
            lcout => \M_this_ext_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40433\,
            ce => 'H',
            sr => \N__39755\
        );

    \M_this_ext_address_q_2_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__40881\,
            in1 => \N__37626\,
            in2 => \N__40722\,
            in3 => \N__37609\,
            lcout => \M_this_ext_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40433\,
            ce => 'H',
            sr => \N__39755\
        );

    \M_this_ext_address_q_3_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__37584\,
            in1 => \N__40884\,
            in2 => \N__37567\,
            in3 => \N__40700\,
            lcout => \M_this_ext_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40433\,
            ce => 'H',
            sr => \N__39755\
        );

    \un1_M_this_ext_address_q_cry_0_c_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37732\,
            in2 => \N__37704\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_24_21_0_\,
            carryout => \un1_M_this_ext_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37667\,
            in2 => \_gnd_net_\,
            in3 => \N__37639\,
            lcout => \un1_M_this_ext_address_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_0\,
            carryout => \un1_M_this_ext_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37625\,
            in2 => \_gnd_net_\,
            in3 => \N__37603\,
            lcout => \un1_M_this_ext_address_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_1\,
            carryout => \un1_M_this_ext_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37583\,
            in2 => \_gnd_net_\,
            in3 => \N__37558\,
            lcout => \un1_M_this_ext_address_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_2\,
            carryout => \un1_M_this_ext_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38625\,
            in2 => \_gnd_net_\,
            in3 => \N__37849\,
            lcout => \un1_M_this_ext_address_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_3\,
            carryout => \un1_M_this_ext_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41229\,
            in2 => \_gnd_net_\,
            in3 => \N__37846\,
            lcout => \un1_M_this_ext_address_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_4\,
            carryout => \un1_M_this_ext_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41184\,
            in2 => \_gnd_net_\,
            in3 => \N__37843\,
            lcout => \un1_M_this_ext_address_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_5\,
            carryout => \un1_M_this_ext_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41136\,
            in3 => \N__37840\,
            lcout => \un1_M_this_ext_address_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_6\,
            carryout => \un1_M_this_ext_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37821\,
            in2 => \_gnd_net_\,
            in3 => \N__37804\,
            lcout => \un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0\,
            ltout => OPEN,
            carryin => \bfn_24_22_0_\,
            carryout => \un1_M_this_ext_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37788\,
            in2 => \_gnd_net_\,
            in3 => \N__37765\,
            lcout => \un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_8\,
            carryout => \un1_M_this_ext_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38652\,
            in2 => \_gnd_net_\,
            in3 => \N__37762\,
            lcout => \un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_9\,
            carryout => \un1_M_this_ext_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41082\,
            in2 => \_gnd_net_\,
            in3 => \N__37759\,
            lcout => \un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_10\,
            carryout => \un1_M_this_ext_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40929\,
            in2 => \_gnd_net_\,
            in3 => \N__37756\,
            lcout => \un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_11\,
            carryout => \un1_M_this_ext_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40488\,
            in3 => \N__38014\,
            lcout => \un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_12\,
            carryout => \un1_M_this_ext_address_q_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38001\,
            in3 => \N__37978\,
            lcout => \un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_13\,
            carryout => \un1_M_this_ext_address_q_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37965\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37948\,
            lcout => \un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37936\,
            in2 => \_gnd_net_\,
            in3 => \N__41564\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37918\,
            in2 => \_gnd_net_\,
            in3 => \N__41565\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38236\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41568\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37891\,
            in2 => \_gnd_net_\,
            in3 => \N__41566\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41569\,
            in2 => \_gnd_net_\,
            in3 => \N__39056\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37867\,
            in2 => \_gnd_net_\,
            in3 => \N__41567\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41574\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38149\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41575\,
            in2 => \_gnd_net_\,
            in3 => \N__38131\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_10_LC_24_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38113\,
            in2 => \_gnd_net_\,
            in3 => \N__39375\,
            lcout => \M_this_oam_ram_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_6_LC_24_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38095\,
            in2 => \_gnd_net_\,
            in3 => \N__39377\,
            lcout => \M_this_oam_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_11_LC_24_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38080\,
            in2 => \_gnd_net_\,
            in3 => \N__39376\,
            lcout => \M_this_oam_ram_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_24_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41573\,
            in2 => \_gnd_net_\,
            in3 => \N__38260\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un12lto7_4_LC_24_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38319\,
            in1 => \N__38340\,
            in2 => \N__38302\,
            in3 => \N__38034\,
            lcout => \this_ppu.un12lto7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_24_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__38035\,
            in1 => \_gnd_net_\,
            in2 => \N__41603\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_24_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41580\,
            in2 => \_gnd_net_\,
            in3 => \N__38341\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_24_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38320\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_24_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38301\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41582\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_24_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38218\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_24_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41576\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un12lto7_5_LC_24_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38256\,
            in1 => \N__38244\,
            in2 => \N__38235\,
            in3 => \N__38217\,
            lcout => \this_ppu.un12lto7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_24_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38200\,
            in2 => \_gnd_net_\,
            in3 => \N__41585\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_3_c_RNO_LC_24_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__38430\,
            in1 => \N__39092\,
            in2 => \N__38563\,
            in3 => \N__39046\,
            lcout => \this_ppu.un1_oam_data_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_24_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38167\,
            in2 => \_gnd_net_\,
            in3 => \N__41586\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_4_c_RNO_LC_24_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001111000011"
        )
    port map (
            in0 => \N__38431\,
            in1 => \N__38500\,
            in2 => \N__38564\,
            in3 => \N__38355\,
            lcout => \this_ppu.un1_oam_data_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_24_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38581\,
            in2 => \_gnd_net_\,
            in3 => \N__41587\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_24_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41589\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_24_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38501\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41588\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_24_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38461\,
            in2 => \_gnd_net_\,
            in3 => \N__41590\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_2_c_RNO_LC_24_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__38415\,
            in1 => \N__39083\,
            in2 => \_gnd_net_\,
            in3 => \N__39034\,
            lcout => \this_ppu.un1_oam_data_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_0_a2_17_LC_24_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38374\,
            in2 => \_gnd_net_\,
            in3 => \N__39374\,
            lcout => \M_this_oam_ram_write_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_4_ac0_1_LC_24_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39081\,
            in2 => \_gnd_net_\,
            in3 => \N__39032\,
            lcout => \this_ppu.un1_oam_data_1_4_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_24_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39154\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_24_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41591\,
            in2 => \_gnd_net_\,
            in3 => \N__39133\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_26_LC_24_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38754\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39373\,
            lcout => \N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_1_c_RNO_LC_24_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39082\,
            in2 => \_gnd_net_\,
            in3 => \N__39033\,
            lcout => \this_ppu.un1_oam_data_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_26_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38998\,
            in1 => \N__38992\,
            in2 => \_gnd_net_\,
            in3 => \N__38929\,
            lcout => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_26_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38965\,
            in1 => \N__38956\,
            in2 => \_gnd_net_\,
            in3 => \N__38928\,
            lcout => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_10_LC_26_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__40710\,
            in2 => \N__38760\,
            in3 => \N__40909\,
            lcout => \M_this_ext_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \M_this_ext_address_q_4_LC_26_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__40907\,
            in1 => \N__38615\,
            in2 => \N__40725\,
            in3 => \N__38638\,
            lcout => \M_this_ext_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \M_this_ext_address_q_5_LC_26_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000001100110"
        )
    port map (
            in0 => \N__41222\,
            in1 => \N__41245\,
            in2 => \N__40723\,
            in3 => \N__40911\,
            lcout => \M_this_ext_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \M_this_ext_address_q_6_LC_26_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__40908\,
            in1 => \N__41177\,
            in2 => \N__40726\,
            in3 => \N__41203\,
            lcout => \M_this_ext_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \M_this_ext_address_q_7_LC_26_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000001100110"
        )
    port map (
            in0 => \N__41120\,
            in1 => \N__41158\,
            in2 => \N__40724\,
            in3 => \N__40912\,
            lcout => \M_this_ext_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \M_this_ext_address_q_11_LC_26_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__40905\,
            in1 => \N__40702\,
            in2 => \N__39505\,
            in3 => \N__41101\,
            lcout => \M_this_ext_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \M_this_ext_address_q_12_LC_26_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__40701\,
            in1 => \N__41065\,
            in2 => \N__41040\,
            in3 => \N__40910\,
            lcout => \M_this_ext_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \M_this_ext_address_q_13_LC_26_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__40906\,
            in1 => \N__40703\,
            in2 => \N__40582\,
            in3 => \N__40501\,
            lcout => \M_this_ext_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40459\,
            ce => 'H',
            sr => \N__39756\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_26_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39538\,
            in2 => \_gnd_net_\,
            in3 => \N__41597\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_oam_ram_write_data_i_i_a2_27_LC_26_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__39440\,
            in1 => \N__39319\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_27_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41638\,
            in2 => \_gnd_net_\,
            in3 => \N__41605\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_28_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41617\,
            in2 => \_gnd_net_\,
            in3 => \N__41604\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1_0_LC_31_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__41344\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41326\,
            lcout => \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_0_LC_32_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__41317\,
            in1 => \N__41311\,
            in2 => \N__41299\,
            in3 => \N__41284\,
            lcout => \this_ppu.N_173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
