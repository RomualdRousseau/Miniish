-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 30 2022 08:36:05

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__35922\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35694\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_data_rw_0_i : std_logic;
signal rgb_c_0 : std_logic;
signal rgb_c_2 : std_logic;
signal rgb_c_4 : std_logic;
signal port_nmib_0_i : std_logic;
signal rgb_c_3 : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal rgb_c_5 : std_logic;
signal rgb_c_1 : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \bfn_7_24_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3\ : std_logic;
signal \this_vga_signals.N_219\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vga_signals.g1_1_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_1_0_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_i4_mux\ : std_logic;
signal \this_vga_signals.if_i4_mux_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_2\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \this_vga_signals.g1_4_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1\ : std_logic;
signal \this_vga_signals.g1_7_cascade_\ : std_logic;
signal \this_vga_signals.N_6_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.N_3_2_0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_3_cascade_\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_vga_signals.g0_0\ : std_logic;
signal \this_vga_signals.g0_5_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0_0_0_0\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal \this_vga_signals.g1_2_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_2\ : std_logic;
signal \this_vga_ramdac.N_24_mux\ : std_logic;
signal \this_vga_ramdac.N_2806_reto\ : std_logic;
signal \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_0_cascade_\ : std_logic;
signal \N_2_0_cascade_\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_vga_ramdac.N_2811_reto\ : std_logic;
signal \this_vga_ramdac.m16\ : std_logic;
signal \this_vga_ramdac.N_2809_reto\ : std_logic;
signal \this_vga_ramdac.i2_mux\ : std_logic;
signal \this_vga_ramdac.N_2808_reto\ : std_logic;
signal \this_vga_ramdac.m6\ : std_logic;
signal \G_463_cascade_\ : std_logic;
signal \this_vga_ramdac.N_2807_reto\ : std_logic;
signal \N_2_0\ : std_logic;
signal \M_this_vga_signals_pixel_clk_0_0\ : std_logic;
signal \G_463\ : std_logic;
signal \this_vga_ramdac.m19\ : std_logic;
signal \this_vga_ramdac.N_2810_reto\ : std_logic;
signal \M_this_map_ram_write_data_0\ : std_logic;
signal \M_this_map_ram_write_data_5\ : std_logic;
signal \M_this_map_ram_write_data_6\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.if_m2_0\ : std_logic;
signal \this_vga_signals.if_m2_1\ : std_logic;
signal \this_vga_signals.if_m2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\ : std_logic;
signal \M_this_vga_ramdac_en_0\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_4\ : std_logic;
signal this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0 : std_logic;
signal this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0 : std_logic;
signal \this_vga_signals.d_N_3_1_i\ : std_logic;
signal \this_vga_signals.M_hcounter_q_RNIO08E8Z0Z_3\ : std_logic;
signal this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3 : std_logic;
signal \this_vga_signals.g1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1_0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3_1_0_0_1\ : std_logic;
signal this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0 : std_logic;
signal \this_vga_signals.N_4_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1\ : std_logic;
signal \this_vga_signals.g1_7\ : std_logic;
signal \this_vga_signals.g0_i_x4_3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_3_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_3_1\ : std_logic;
signal \this_vga_signals.N_6_1_0\ : std_logic;
signal \this_vga_signals.N_234\ : std_logic;
signal \this_vga_signals.SUM_3_cascade_\ : std_logic;
signal \this_vga_signals.g0_6_1\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_1\ : std_logic;
signal \this_vga_signals.g1_2_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.SUM_3_0_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_0\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal this_vga_signals_hvisibility_i : std_logic;
signal \this_vga_signals.g3_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g3_0\ : std_logic;
signal \this_vga_signals.g3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_2\ : std_logic;
signal \this_vga_signals.g0_0_a2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_a2_1\ : std_logic;
signal \this_vga_signals.vaddress_1_5\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_ns\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_ns_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\ : std_logic;
signal \this_vga_signals.g0_i_x4_1\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_2_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_3\ : std_logic;
signal \this_vga_signals.g0_2_0_a2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_vga_signals.g0_1_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_x1\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.g0_i_x4_2_0_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_0\ : std_logic;
signal \this_vga_signals.N_3_cascade_\ : std_logic;
signal \this_vga_signals.N_4_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c2_0_0_0\ : std_logic;
signal \this_vga_signals.g0_2_1\ : std_logic;
signal \this_vga_signals.N_5_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_a0_0\ : std_logic;
signal \this_vga_signals.SUM_3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2\ : std_logic;
signal \this_vga_signals.if_N_6_0\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \this_vga_signals.un4_hsynclt9\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_1_cascade_\ : std_logic;
signal \N_3_0\ : std_logic;
signal \N_3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_3_1\ : std_logic;
signal \this_vga_signals.g1_2\ : std_logic;
signal \this_vga_signals.SUM_3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_0\ : std_logic;
signal \M_this_map_ram_write_data_4\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i_0\ : std_logic;
signal \this_vga_signals.N_18_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0_1\ : std_logic;
signal \this_vga_signals.vaddress_1_6\ : std_logic;
signal \this_vga_signals.N_6_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_661_cascade_\ : std_logic;
signal \this_vga_signals.g0_2_0_a2_1\ : std_logic;
signal \this_vga_signals.if_N_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.N_4_0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_0_a2_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1_661\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_a3_2\ : std_logic;
signal \this_vga_signals.vaddress_0_6\ : std_logic;
signal \this_vga_signals.g0_i_x4_0_a3_0\ : std_logic;
signal \this_vga_signals.vsync_1_3\ : std_logic;
signal \this_vga_signals.vsync_1_2_cascade_\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_vga_signals.un2_vsynclt8\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_0_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un2_hsynclto3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lto7_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt7_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.N_852_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.un2_hsynclt6_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.un2_hsynclt7\ : std_logic;
signal \this_vga_signals.un2_hsynclto3_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un4_hsynclto7_0\ : std_logic;
signal \M_this_map_ram_write_data_1\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_1_1_3\ : std_logic;
signal \this_vga_signals.N_1_3_1_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_2_3\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_2_3_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_1_3\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_i\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_N_2L1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_x1\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_d_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.g2_0_a2_5Z0Z_1_cascade_\ : std_logic;
signal \this_vga_signals.g2_0_a2_2\ : std_logic;
signal \this_vga_signals.g2_0_a2_5\ : std_logic;
signal \this_vga_signals.g2\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.g1_3\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.if_m2\ : std_logic;
signal \this_vga_signals.N_1098_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_0_N_2L1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.vaddress_c3_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.if_m8_0_a3_1_1_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylto8_0_cascade_\ : std_logic;
signal \this_vga_signals.un6_vvisibilitylt9_0_cascade_\ : std_logic;
signal \this_vga_signals_vvisibility_1_cascade_\ : std_logic;
signal \this_vga_signals.vvisibility\ : std_logic;
signal \this_vga_signals.vaddress_ac0_9_0_a0_0\ : std_logic;
signal \this_ppu.N_1195_0_1_cascade_\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_6_s1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal port_clk_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals.N_852_0\ : std_logic;
signal \this_vga_signals.N_1098_g\ : std_logic;
signal \this_ppu.N_1195_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_1195_0_1\ : std_logic;
signal \this_ppu.M_count_qZ0Z_0\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\ : std_logic;
signal \this_ppu.M_count_qZ0Z_5\ : std_logic;
signal \this_ppu.M_count_qZ0Z_4\ : std_logic;
signal \this_ppu.M_count_qZ0Z_6\ : std_logic;
signal \this_ppu.M_count_qZ0Z_2\ : std_logic;
signal \this_ppu.M_count_qZ0Z_1\ : std_logic;
signal \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4_cascade_\ : std_logic;
signal \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3\ : std_logic;
signal \this_ppu.un16_0\ : std_logic;
signal \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\ : std_logic;
signal \this_ppu.N_1195_0\ : std_logic;
signal \this_ppu.M_count_qZ0Z_3\ : std_logic;
signal \this_ppu.M_count_q_RNO_0Z0Z_7\ : std_logic;
signal \this_ppu.M_count_qZ0Z_7\ : std_logic;
signal \this_vga_signals.N_85_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_5\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0Z0Z_2_cascade_\ : std_logic;
signal \M_this_substate_qZ0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \M_this_map_ram_write_data_3\ : std_logic;
signal \M_this_map_ram_write_data_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lto8_1\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt8_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.line_clk_1_cascade_\ : std_logic;
signal \M_this_vga_signals_line_clk_0_cascade_\ : std_logic;
signal \this_vga_signals.un4_lvisibility_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.line_clk_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.CO0\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal \this_pixel_clk_M_counter_q_0\ : std_logic;
signal \this_vga_signals.N_152_0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_WE_6\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_i_1Z0Z_10\ : std_logic;
signal \this_sprites_ram.mem_WE_10\ : std_logic;
signal \this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_6\ : std_logic;
signal \this_vga_signals.N_85\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_4\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_1Z0Z_11\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0Z0Z_3\ : std_logic;
signal \M_this_state_d_0_sqmuxa_1\ : std_logic;
signal \M_this_map_ram_write_data_7\ : std_logic;
signal \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\ : std_logic;
signal \G_425\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_vcounter_d8\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d7_1_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_vga_signals.N_153_0_cascade_\ : std_logic;
signal \N_686_i_cascade_\ : std_logic;
signal \N_164\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_8\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_8_cascade_\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_8\ : std_logic;
signal \this_vga_signals.N_124_0\ : std_logic;
signal \this_vga_signals.N_154_cascade_\ : std_logic;
signal \this_vga_signals.N_97\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_2_0\ : std_logic;
signal \this_vga_signals.N_154\ : std_logic;
signal \this_vga_signals.N_62_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0\ : std_logic;
signal \M_this_map_ram_read_data_2\ : std_logic;
signal \M_this_ppu_sprites_addr_8\ : std_logic;
signal \M_this_map_ram_read_data_1\ : std_logic;
signal \M_this_ppu_sprites_addr_7\ : std_logic;
signal port_address_in_7 : std_logic;
signal led_c_1 : std_logic;
signal \N_84\ : std_logic;
signal port_address_in_1 : std_logic;
signal port_address_in_4 : std_logic;
signal port_address_in_0 : std_logic;
signal \N_36\ : std_logic;
signal port_dmab_c_i : std_logic;
signal \this_ppu.un1_M_oam_idx_q_1_c1_cascade_\ : std_logic;
signal \this_ppu.un1_M_oam_idx_q_1_c3_cascade_\ : std_logic;
signal \this_ppu.M_count_d_0_sqmuxa_1_7\ : std_logic;
signal \this_ppu.un1_M_oam_idx_q_1_c3\ : std_logic;
signal \this_ppu.un1_M_oam_idx_q_1_c1\ : std_logic;
signal \this_ppu.N_1156_0\ : std_logic;
signal \M_this_ppu_oam_addr_2\ : std_logic;
signal \M_this_ppu_oam_addr_1\ : std_logic;
signal \this_ppu.M_oam_idx_qZ0Z_4\ : std_logic;
signal \M_this_ppu_oam_addr_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c5\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_0\ : std_logic;
signal \this_ppu.un2_hscroll_axb_0_cascade_\ : std_logic;
signal \M_this_ppu_sprites_addr_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_3_c2\ : std_logic;
signal \this_ppu.M_state_q_RNIGL6V4Z0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_3\ : std_logic;
signal \this_sprites_ram.mem_WE_8\ : std_logic;
signal \N_686_i\ : std_logic;
signal \M_this_data_count_qlde_i_i\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_q_cry_1_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_data_count_q_s_6\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \M_this_data_count_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \M_this_data_count_q_cry_7_THRU_CO\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \M_this_data_count_q_cry_8_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \M_this_data_count_q_s_10\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_q_cry_10_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \M_this_data_count_q_cry_11_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal \M_this_data_count_q_s_13\ : std_logic;
signal \N_49\ : std_logic;
signal this_vga_signals_vvisibility_1 : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c5\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_1\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_2\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_3\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_5\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_6\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_cry_7\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_4\ : std_logic;
signal \this_ppu.N_148\ : std_logic;
signal \this_ppu.vscroll8\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_5\ : std_logic;
signal \this_ppu.M_state_qZ0Z_4\ : std_logic;
signal \M_this_ppu_oam_addr_3\ : std_logic;
signal \this_ppu.N_144_4\ : std_logic;
signal \this_ppu.M_state_qZ0Z_2\ : std_logic;
signal \this_ppu.N_144\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\ : std_logic;
signal \M_this_ppu_vram_data_0\ : std_logic;
signal \M_this_ppu_vram_data_0_cascade_\ : std_logic;
signal \this_ppu.N_156_cascade_\ : std_logic;
signal \M_this_ppu_vram_en_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_0\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_3\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_3\ : std_logic;
signal \this_ppu.N_156\ : std_logic;
signal \this_ppu.N_150\ : std_logic;
signal \this_ppu.M_state_qZ0Z_5\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_3\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_3\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \M_this_state_q_RNIH92SZ0Z_10_cascade_\ : std_logic;
signal \this_vga_signals.N_83\ : std_logic;
signal \this_vga_signals.N_94_0\ : std_logic;
signal \this_vga_signals.N_94_0_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_i_0Z0Z_12\ : std_logic;
signal \M_this_state_q_RNI373A1Z0Z_8\ : std_logic;
signal \this_vga_signals_un21_i_a3_1_1_cascade_\ : std_logic;
signal port_dmab_c : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_8\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_a3_0_7_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_0Z0Z_7_cascade_\ : std_logic;
signal \M_this_state_q_RNI6Q0SZ0Z_5\ : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \N_848\ : std_logic;
signal \this_vga_signals.N_93_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \M_this_vga_signals_line_clk_0\ : std_logic;
signal \this_ppu.M_last_q\ : std_logic;
signal \this_ppu.N_132_0\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_2_c2\ : std_logic;
signal \this_ppu.M_state_q_RNILG0GDZ0Z_0\ : std_logic;
signal \bfn_19_17_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_0\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_1\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_2\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_3\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_4\ : std_logic;
signal \M_this_ppu_map_addr_8\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_5\ : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_7\ : std_logic;
signal \bfn_19_18_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_3\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_0\ : std_logic;
signal \bfn_19_19_0_\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_0\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_1\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_0\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_2\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_1\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_3\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_2\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_4\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_3\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_4\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_haddress_q_cry_7\ : std_logic;
signal \bfn_19_20_0_\ : std_logic;
signal \this_ppu.vscroll8_1\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_4\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_1\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus7_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus3_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus4_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus0_2\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\ : std_logic;
signal \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\ : std_logic;
signal \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\ : std_logic;
signal \M_this_ppu_vram_data_2\ : std_logic;
signal \M_this_map_ram_read_data_0\ : std_logic;
signal \M_this_ppu_sprites_addr_6\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_2\ : std_logic;
signal \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\ : std_logic;
signal \N_792\ : std_logic;
signal \M_this_sprites_address_qc_0_0_0\ : std_logic;
signal \N_795\ : std_logic;
signal \N_773_0\ : std_logic;
signal \N_773_0_cascade_\ : std_logic;
signal \this_vga_signals.N_485\ : std_logic;
signal \N_17\ : std_logic;
signal \N_126\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \port_dmab_ac0_1_3_cascade_\ : std_logic;
signal port_dmab_ac0_1_4 : std_logic;
signal \N_15\ : std_logic;
signal \N_809_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \N_775_0\ : std_logic;
signal \N_775_0_cascade_\ : std_logic;
signal port_address_in_5 : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0Z0Z_0\ : std_logic;
signal \N_87_0_cascade_\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal port_enb_c : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_4\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \this_ppu.M_this_ppu_vram_addr_i_7\ : std_logic;
signal \bfn_20_19_0_\ : std_logic;
signal \this_ppu.M_vaddress_q_i_1\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_0\ : std_logic;
signal \this_ppu.M_vaddress_q_i_2\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_1\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_5\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_2\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_3\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_7\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_4\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_8\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_5\ : std_logic;
signal \this_ppu.M_this_ppu_map_addr_i_9\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_6\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_7\ : std_logic;
signal \bfn_20_20_0_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_11\ : std_logic;
signal \M_this_state_qZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_1\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_2\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_2\ : std_logic;
signal \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_0\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\ : std_logic;
signal \M_this_sprites_address_qc_0_0\ : std_logic;
signal \this_sprites_ram.mem_WE_14\ : std_logic;
signal \M_this_sprites_address_qZ0Z_0\ : std_logic;
signal \N_443_i\ : std_logic;
signal \M_this_sprites_address_q_RNO_0Z0Z_0\ : std_logic;
signal \bfn_21_13_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_1\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_2\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_3\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_5\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_6\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_7\ : std_logic;
signal \bfn_21_14_0_\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_8\ : std_logic;
signal \M_this_sprites_address_qZ0Z_10\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_9\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_11\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_10\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_11\ : std_logic;
signal \M_this_sprites_address_qc_2_1\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_12\ : std_logic;
signal \M_this_sprites_address_q_RNO_0Z0Z_12\ : std_logic;
signal \N_807_cascade_\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_7\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_8\ : std_logic;
signal \N_803_cascade_\ : std_logic;
signal \M_this_sprites_address_qc_10_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_8\ : std_logic;
signal \N_602\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_7\ : std_logic;
signal \M_this_sprites_address_qc_9_0\ : std_logic;
signal \M_this_oam_ram_read_data_i_19\ : std_logic;
signal \M_this_oam_ram_read_data_i_11\ : std_logic;
signal \M_this_oam_ram_read_data_15\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_7\ : std_logic;
signal \M_this_oam_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_oam_address_q_c4\ : std_logic;
signal \M_this_oam_address_qZ0Z_5\ : std_logic;
signal \M_this_oam_address_qZ0Z_3\ : std_logic;
signal \M_this_data_tmp_qZ0Z_2\ : std_logic;
signal \N_746_0\ : std_logic;
signal \M_this_oam_ram_write_data_28\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \un1_M_this_sprites_address_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_sprites_address_q_RNO_0Z0Z_2\ : std_logic;
signal \N_813\ : std_logic;
signal \N_799\ : std_logic;
signal \M_this_sprites_address_qc_11_0_cascade_\ : std_logic;
signal \M_this_sprites_address_q_RNO_1Z0Z_9\ : std_logic;
signal \M_this_sprites_address_qZ0Z_9\ : std_logic;
signal \M_this_sprites_address_q_RNO_0Z0Z_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_3\ : std_logic;
signal \N_50\ : std_logic;
signal \M_this_ppu_sprites_addr_3\ : std_logic;
signal \M_this_sprites_address_qZ0Z_2\ : std_logic;
signal \N_103\ : std_logic;
signal \M_this_sprites_ram_write_data_iv_i_i_1\ : std_logic;
signal port_address_in_3 : std_logic;
signal port_address_in_2 : std_logic;
signal port_rw_in : std_logic;
signal port_address_in_6 : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_4_0\ : std_logic;
signal \N_54_0\ : std_logic;
signal \this_ppu.un1_oam_data_1_c2\ : std_logic;
signal \N_163\ : std_logic;
signal \un1_M_this_oam_address_q_c2\ : std_logic;
signal \M_this_oam_address_qZ0Z_2\ : std_logic;
signal \N_1190_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_6\ : std_logic;
signal \N_742_0\ : std_logic;
signal \N_34_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_4\ : std_logic;
signal \N_744_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_7\ : std_logic;
signal \N_56_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_16\ : std_logic;
signal \N_738_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_22\ : std_logic;
signal \N_40_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus6_0\ : std_logic;
signal \this_sprites_ram.mem_out_bus2_0\ : std_logic;
signal \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\ : std_logic;
signal \N_102\ : std_logic;
signal \M_this_sprites_address_q_RNO_0Z0Z_4\ : std_logic;
signal \M_this_sprites_address_qZ0Z_4\ : std_logic;
signal \N_101_cascade_\ : std_logic;
signal \M_this_sprites_address_q_RNO_0Z0Z_6\ : std_logic;
signal \M_this_sprites_address_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_3_bmZ0Z_1\ : std_logic;
signal \M_this_sprites_address_qZ0Z_1\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \N_87_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_q_3_amZ0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_this_state_q_3_0_i_0_0\ : std_logic;
signal \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2\ : std_logic;
signal \M_this_sprites_ram_write_data_iv_i_i_3\ : std_logic;
signal \this_ppu.un2_vscroll_axb_0\ : std_logic;
signal \M_this_ppu_sprites_addr_1\ : std_logic;
signal \M_this_data_tmp_qZ0Z_8\ : std_logic;
signal \N_1182_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_3\ : std_logic;
signal \N_745_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_14\ : std_logic;
signal \N_739_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_5\ : std_logic;
signal \N_743_0\ : std_logic;
signal \N_32_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_11\ : std_logic;
signal \M_this_oam_ram_write_data_11\ : std_logic;
signal \M_this_data_tmp_qZ0Z_0\ : std_logic;
signal \N_748_0\ : std_logic;
signal \N_44_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_17\ : std_logic;
signal \N_1174_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_23\ : std_logic;
signal \M_this_oam_ram_write_data_23\ : std_logic;
signal \M_this_data_tmp_qZ0Z_20\ : std_logic;
signal \N_42_0\ : std_logic;
signal \M_this_oam_ram_write_data_30\ : std_logic;
signal \this_sprites_ram.mem_out_bus5_1\ : std_logic;
signal \this_sprites_ram.mem_out_bus1_1\ : std_logic;
signal \this_sprites_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\ : std_logic;
signal \M_this_ppu_sprites_addr_2\ : std_logic;
signal \this_sprites_ram.mem_WE_4\ : std_logic;
signal \this_sprites_ram.mem_WE_12\ : std_logic;
signal \M_this_ppu_sprites_addr_5\ : std_logic;
signal \N_809\ : std_logic;
signal \M_this_sprites_address_q_RNO_0Z0Z_5\ : std_logic;
signal \N_595\ : std_logic;
signal \N_383_0\ : std_logic;
signal \M_this_sprites_address_qZ0Z_5\ : std_logic;
signal \N_515_g\ : std_logic;
signal \this_sprites_ram.mem_WE_0\ : std_logic;
signal \M_this_ppu_sprites_addr_4\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \M_this_oam_ram_read_data_16\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_16\ : std_logic;
signal \bfn_24_16_0_\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_1\ : std_logic;
signal \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\ : std_logic;
signal \this_ppu.un2_vscroll_cry_0\ : std_logic;
signal \this_ppu.M_vaddress_qZ0Z_2\ : std_logic;
signal \M_this_oam_ram_read_data_18\ : std_logic;
signal \this_ppu.un2_vscroll_cry_1\ : std_logic;
signal \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \M_this_ppu_sprites_addr_10\ : std_logic;
signal \M_this_sprites_address_qZ0Z_11\ : std_logic;
signal \M_this_sprites_address_qZ0Z_12\ : std_logic;
signal \M_this_sprites_address_qZ0Z_13\ : std_logic;
signal \N_23_0\ : std_logic;
signal \this_sprites_ram.mem_WE_2\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_oam_ram_read_data_8\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\ : std_logic;
signal \bfn_24_19_0_\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\ : std_logic;
signal \this_ppu.un2_hscroll_cry_0\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \M_this_oam_ram_read_data_10\ : std_logic;
signal \this_ppu.un2_hscroll_cry_1\ : std_logic;
signal \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\ : std_logic;
signal \M_this_oam_ram_read_data_9\ : std_logic;
signal \M_this_oam_ram_read_data_i_9\ : std_logic;
signal \M_this_data_tmp_qZ0Z_1\ : std_logic;
signal \N_747_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_10\ : std_logic;
signal \M_this_oam_ram_write_data_10\ : std_logic;
signal \M_this_map_ram_read_data_3\ : std_logic;
signal \this_ppu.M_state_qZ0Z_6\ : std_logic;
signal \this_ppu.M_state_qZ0Z_7\ : std_logic;
signal \M_this_ppu_sprites_addr_9\ : std_logic;
signal \M_this_data_tmp_qZ0Z_12\ : std_logic;
signal \N_740_0\ : std_logic;
signal \M_this_oam_ram_read_data_13\ : std_logic;
signal \M_this_oam_ram_read_data_12\ : std_logic;
signal \M_this_oam_ram_read_data_14\ : std_logic;
signal \M_this_oam_ram_read_data_11\ : std_logic;
signal \this_ppu.un1_M_haddress_q_2_6\ : std_logic;
signal \M_this_data_tmp_qZ0Z_19\ : std_logic;
signal \M_this_oam_ram_write_data_19\ : std_logic;
signal \M_this_oam_ram_read_data_6\ : std_logic;
signal \M_this_oam_ram_read_data_5\ : std_logic;
signal \M_this_oam_ram_read_data_7\ : std_logic;
signal \M_this_oam_ram_read_data_4\ : std_logic;
signal \this_ppu.un9lto7Z0Z_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_9\ : std_logic;
signal \N_741_0\ : std_logic;
signal \M_this_oam_ram_read_data_23\ : std_logic;
signal \this_ppu.un1_oam_data_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_13\ : std_logic;
signal \M_this_oam_ram_write_data_13\ : std_logic;
signal \M_this_data_tmp_qZ0Z_15\ : std_logic;
signal \M_this_oam_ram_write_data_15\ : std_logic;
signal \N_123_0\ : std_logic;
signal \M_this_oam_ram_read_data_2\ : std_logic;
signal \M_this_oam_ram_read_data_1\ : std_logic;
signal \M_this_oam_ram_read_data_3\ : std_logic;
signal \M_this_oam_ram_read_data_0\ : std_logic;
signal \this_ppu.un9lto7Z0Z_5\ : std_logic;
signal \M_this_oam_ram_read_data_17\ : std_logic;
signal \M_this_oam_ram_read_data_i_17\ : std_logic;
signal \M_this_data_tmp_qZ0Z_18\ : std_logic;
signal \M_this_oam_ram_write_data_18\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_5\ : std_logic;
signal \N_38_0\ : std_logic;
signal \M_this_oam_ram_write_data_31\ : std_logic;
signal \N_736_0\ : std_logic;
signal \N_737_0\ : std_logic;
signal \M_this_oam_ram_read_data_21\ : std_logic;
signal \M_this_oam_ram_read_data_20\ : std_logic;
signal \M_this_oam_ram_read_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_19\ : std_logic;
signal \this_ppu.un1_M_vaddress_q_3_6\ : std_logic;
signal \M_this_oam_address_qZ0Z_0\ : std_logic;
signal \M_this_oam_address_qZ0Z_1\ : std_logic;
signal \M_this_data_tmp_qZ0Z_21\ : std_logic;
signal \N_122_0\ : std_logic;
signal \M_this_oam_ram_write_data_21\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_5\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_6\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_7\ : std_logic;
signal \un1_M_this_state_q_9_0_i\ : std_logic;
signal \M_this_external_address_qZ0Z_0\ : std_logic;
signal \bfn_28_21_0_\ : std_logic;
signal \M_this_external_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_external_address_q_cry_0\ : std_logic;
signal \M_this_external_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_external_address_q_cry_1\ : std_logic;
signal \M_this_external_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_external_address_q_cry_2\ : std_logic;
signal \M_this_external_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_external_address_q_cry_3\ : std_logic;
signal \M_this_external_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_external_address_q_cry_4\ : std_logic;
signal \M_this_external_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_5\ : std_logic;
signal \M_this_external_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_external_address_q_cry_6\ : std_logic;
signal \un1_M_this_external_address_q_cry_7\ : std_logic;
signal port_data_c_0 : std_logic;
signal \M_this_external_address_qZ0Z_8\ : std_logic;
signal \bfn_28_22_0_\ : std_logic;
signal port_data_c_1 : std_logic;
signal \M_this_external_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_external_address_q_cry_8\ : std_logic;
signal port_data_c_2 : std_logic;
signal \M_this_external_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_external_address_q_cry_9\ : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_external_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_external_address_q_cry_10\ : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_external_address_qZ0Z_12\ : std_logic;
signal \un1_M_this_external_address_q_cry_11\ : std_logic;
signal port_data_c_5 : std_logic;
signal \M_this_external_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_external_address_q_cry_12\ : std_logic;
signal port_data_c_6 : std_logic;
signal \M_this_external_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_external_address_q_cry_13\ : std_logic;
signal \N_749_0\ : std_logic;
signal port_data_c_7 : std_logic;
signal \un1_M_this_external_address_q_cry_14\ : std_logic;
signal \M_this_external_address_qZ0Z_15\ : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_8\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal clk_0_c_g : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_map_ram_read_data_3\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_2\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_1\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_0\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__22140\&\N__21819\&\N__21867\&\N__21906\&\N__21957\&\N__20424\&\N__20490\&\N__20568\&\N__20631\&\N__20271\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__11217\&\N__11250\&\N__11280\&\N__11310\&\N__11340\&\N__11370\&\N__11022\&\N__11052\&\N__11082\&\N__11109\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__16197\&'0'&'0'&'0'&\N__16185\&'0'&'0'&'0'&\N__13986\&'0'&'0'&'0'&\N__11958\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__22134\&\N__21813\&\N__21861\&\N__21900\&\N__21951\&\N__20418\&\N__20484\&\N__20562\&\N__20625\&\N__20265\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__11211\&\N__11244\&\N__11274\&\N__11304\&\N__11334\&\N__11364\&\N__11016\&\N__11046\&\N__11076\&\N__11103\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__17331\&'0'&'0'&'0'&\N__11940\&'0'&'0'&'0'&\N__11952\&'0'&'0'&'0'&\N__13215\&'0';
    \M_this_oam_ram_read_data_15\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_14\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_13\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_12\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_11\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_10\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_9\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_8\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_7\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_6\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_5\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_4\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_3\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_2\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_1\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_0\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20862\&\N__19056\&\N__19011\&\N__18954\;
    \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24822\&\N__24876\&\N__24789\&\N__26421\;
    \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ <= \N__32043\&\N__28149\&\N__32067\&\N__31074\&\N__28383\&\N__31713\&\N__32130\&\N__26517\&\N__26931\&\N__26343\&\N__28125\&\N__26952\&\N__28173\&\N__25278\&\N__31734\&\N__28362\;
    \M_this_oam_ram_read_data_23\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_22\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_21\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_20\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_19\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_18\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_17\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_16\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20856\&\N__19050\&\N__19005\&\N__18948\;
    \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__24816\&\N__24870\&\N__24783\&\N__26415\;
    \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ <= \N__33093\&\N__29685\&\N__33087\&\N__25263\&\N__28407\&\N__26331\&\N__33081\&\N__33102\&\N__28260\&\N__26889\&\N__32265\&\N__28239\&\N__30867\&\N__33132\&\N__28350\&\N__26910\;
    \this_sprites_ram.mem_out_bus0_1\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_0\ <= \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__30493\&\N__31334\&\N__18325\&\N__18096\&\N__22535\&\N__29315\&\N__28591\&\N__25785\&\N__29522\&\N__27180\&\N__18858\;
    \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__24366\&\N__26227\&\N__24711\&\N__25169\&\N__28101\&\N__28859\&\N__26821\&\N__26000\&\N__25544\&\N__27891\&\N__23988\;
    \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25370\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22818\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus0_3\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus0_2\ <= \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__30475\&\N__31314\&\N__18313\&\N__18092\&\N__22487\&\N__29297\&\N__28592\&\N__25784\&\N__29521\&\N__27179\&\N__18854\;
    \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__24365\&\N__26208\&\N__24707\&\N__25157\&\N__28100\&\N__28858\&\N__26820\&\N__26019\&\N__25590\&\N__27890\&\N__23987\;
    \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27273\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23100\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_1\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_0\ <= \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__30474\&\N__31325\&\N__18292\&\N__18085\&\N__22530\&\N__29299\&\N__28570\&\N__25776\&\N__29503\&\N__27172\&\N__18844\;
    \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__24357\&\N__26207\&\N__24698\&\N__25170\&\N__28091\&\N__28838\&\N__26801\&\N__26004\&\N__25584\&\N__27877\&\N__23977\;
    \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25362\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22813\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus1_3\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus1_2\ <= \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__30453\&\N__31291\&\N__18327\&\N__18075\&\N__22506\&\N__29268\&\N__28574\&\N__25761\&\N__29499\&\N__27161\&\N__18843\;
    \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__24343\&\N__26182\&\N__24679\&\N__25114\&\N__28090\&\N__28837\&\N__26800\&\N__25977\&\N__25569\&\N__27876\&\N__23976\;
    \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27276\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23095\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_1\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_0\ <= \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__30452\&\N__31307\&\N__18321\&\N__18063\&\N__22511\&\N__29277\&\N__28540\&\N__25739\&\N__29474\&\N__27144\&\N__18816\;
    \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__24319\&\N__26181\&\N__24650\&\N__25155\&\N__28065\&\N__28806\&\N__26749\&\N__26005\&\N__25547\&\N__27842\&\N__23950\;
    \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25349\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22800\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus2_3\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus2_2\ <= \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__30519\&\N__31335\&\N__18326\&\N__18021\&\N__22527\&\N__29325\&\N__28608\&\N__25783\&\N__29547\&\N__27097\&\N__18832\;
    \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__24356\&\N__26238\&\N__24706\&\N__25168\&\N__28099\&\N__28869\&\N__26822\&\N__26021\&\N__25589\&\N__27888\&\N__23985\;
    \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27275\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23099\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_1\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_0\ <= \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__30515\&\N__31261\&\N__18248\&\N__18020\&\N__22525\&\N__29324\&\N__28604\&\N__25772\&\N__29543\&\N__27160\&\N__18831\;
    \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__24339\&\N__26237\&\N__24705\&\N__25158\&\N__28086\&\N__28868\&\N__26811\&\N__26020\&\N__25588\&\N__27887\&\N__23984\;
    \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25371\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22817\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus3_3\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus3_2\ <= \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__30514\&\N__31330\&\N__18317\&\N__18019\&\N__22528\&\N__29316\&\N__28603\&\N__25771\&\N__29507\&\N__27159\&\N__18790\;
    \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__24270\&\N__26230\&\N__24691\&\N__25176\&\N__28085\&\N__28861\&\N__26810\&\N__26008\&\N__25577\&\N__27886\&\N__23964\;
    \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27274\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23091\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_1\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_0\ <= \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__30507\&\N__31329\&\N__18299\&\N__18018\&\N__22524\&\N__29284\&\N__28593\&\N__25751\&\N__29535\&\N__27137\&\N__18829\;
    \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__24337\&\N__26228\&\N__24690\&\N__25172\&\N__28083\&\N__28824\&\N__26808\&\N__26018\&\N__25531\&\N__27884\&\N__23963\;
    \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25366\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22807\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus4_3\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus4_2\ <= \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__30494\&\N__31315\&\N__18272\&\N__18017\&\N__22526\&\N__29323\&\N__28578\&\N__25701\&\N__29542\&\N__27171\&\N__18830\;
    \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__24338\&\N__26229\&\N__24689\&\N__25171\&\N__28084\&\N__28860\&\N__26809\&\N__26022\&\N__25576\&\N__27885\&\N__23925\;
    \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27262\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23077\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_1\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_0\ <= \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__30428\&\N__31262\&\N__18306\&\N__18051\&\N__22464\&\N__29229\&\N__28547\&\N__25713\&\N__29419\&\N__27122\&\N__18789\;
    \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__24215\&\N__26150\&\N__24616\&\N__25130\&\N__28064\&\N__28805\&\N__26750\&\N__25983\&\N__25519\&\N__27855\&\N__23949\;
    \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25348\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22811\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus5_3\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus5_2\ <= \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__30427\&\N__31281\&\N__18282\&\N__18038\&\N__22507\&\N__29191\&\N__28504\&\N__25682\&\N__29455\&\N__27098\&\N__18803\;
    \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__24283\&\N__26141\&\N__24642\&\N__25129\&\N__28020\&\N__28730\&\N__26748\&\N__25984\&\N__25471\&\N__27831\&\N__23948\;
    \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27251\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23072\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_1\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_0\ <= \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__30394\&\N__31227\&\N__18249\&\N__18022\&\N__22480\&\N__29236\&\N__28469\&\N__25651\&\N__29491\&\N__27073\&\N__18833\;
    \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__24297\&\N__26142\&\N__24603\&\N__25127\&\N__28039\&\N__28765\&\N__26790\&\N__25982\&\N__25511\&\N__27832\&\N__23938\;
    \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25330\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22793\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus6_3\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus6_2\ <= \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__30367\&\N__31248\&\N__18180\&\N__17999\&\N__22529\&\N__29272\&\N__28514\&\N__25694\&\N__29492\&\N__27046\&\N__18851\;
    \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__24332\&\N__26143\&\N__24643\&\N__25128\&\N__28078\&\N__28819\&\N__26815\&\N__25981\&\N__25512\&\N__27871\&\N__23971\;
    \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27252\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23073\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_1\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_0\ <= \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__30425\&\N__31190\&\N__18261\&\N__18034\&\N__22531\&\N__29273\&\N__28554\&\N__25725\&\N__29519\&\N__27020\&\N__18852\;
    \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__24333\&\N__26179\&\N__24677\&\N__25113\&\N__28079\&\N__28820\&\N__26816\&\N__26006\&\N__25545\&\N__27872\&\N__23972\;
    \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__25342\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__22812\&'0'&'0'&'0';
    \this_sprites_ram.mem_out_bus7_3\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_sprites_ram.mem_out_bus7_2\ <= \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__30426\&\N__31133\&\N__18262\&\N__18050\&\N__22536\&\N__29298\&\N__28555\&\N__25726\&\N__29520\&\N__27061\&\N__18853\;
    \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__24364\&\N__26180\&\N__24678\&\N__25156\&\N__28098\&\N__28845\&\N__26823\&\N__26007\&\N__25546\&\N__27889\&\N__23986\;
    \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__27269\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23090\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__12195\&\N__11457\&\N__11190\&\N__11181\&\N__11499\&\N__12084\&\N__11469\&\N__11529\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__30855\&\N__20480\&\N__20561\&\N__20618\&\N__20264\&\N__29757\&\N__29836\&\N__29969\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21138\&\N__22581\&\N__22713\&\N__20763\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34633\,
            RE => \N__19658\,
            WCLKE => \N__17434\,
            WCLK => \N__34634\,
            WE => \N__19667\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34640\,
            RE => \N__19581\,
            WCLKE => \N__17435\,
            WCLK => \N__34641\,
            WE => \N__19617\
        );

    \this_oam_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34629\,
            RE => \N__19822\,
            WCLKE => \N__32033\,
            WCLK => \N__34630\,
            WE => \N__19746\
        );

    \this_oam_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34635\,
            RE => \N__19744\,
            WCLKE => \N__32037\,
            WCLK => \N__34636\,
            WE => \N__19745\
        );

    \this_sprites_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34518\,
            RE => \N__20100\,
            WCLKE => \N__24018\,
            WCLK => \N__34519\,
            WE => \N__20012\
        );

    \this_sprites_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34528\,
            RE => \N__19887\,
            WCLKE => \N__24017\,
            WCLK => \N__34529\,
            WE => \N__20092\
        );

    \this_sprites_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34542\,
            RE => \N__20097\,
            WCLKE => \N__29343\,
            WCLK => \N__34543\,
            WE => \N__20091\
        );

    \this_sprites_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34558\,
            RE => \N__20096\,
            WCLKE => \N__29342\,
            WCLK => \N__34559\,
            WE => \N__20057\
        );

    \this_sprites_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34573\,
            RE => \N__20068\,
            WCLKE => \N__16955\,
            WCLK => \N__34572\,
            WE => \N__20056\
        );

    \this_sprites_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34550\,
            RE => \N__20080\,
            WCLKE => \N__16962\,
            WCLK => \N__34551\,
            WE => \N__20076\
        );

    \this_sprites_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34565\,
            RE => \N__19809\,
            WCLKE => \N__19080\,
            WCLK => \N__34564\,
            WE => \N__20075\
        );

    \this_sprites_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34578\,
            RE => \N__20023\,
            WCLKE => \N__19076\,
            WCLK => \N__34579\,
            WE => \N__19878\
        );

    \this_sprites_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34592\,
            RE => \N__20013\,
            WCLKE => \N__16995\,
            WCLK => \N__34593\,
            WE => \N__19877\
        );

    \this_sprites_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34603\,
            RE => \N__19865\,
            WCLKE => \N__16991\,
            WCLK => \N__34604\,
            WE => \N__19802\
        );

    \this_sprites_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34586\,
            RE => \N__20067\,
            WCLKE => \N__29354\,
            WCLK => \N__34587\,
            WE => \N__20085\
        );

    \this_sprites_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34599\,
            RE => \N__20099\,
            WCLKE => \N__29361\,
            WCLK => \N__34600\,
            WE => \N__19987\
        );

    \this_sprites_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34607\,
            RE => \N__19913\,
            WCLKE => \N__29985\,
            WCLK => \N__34608\,
            WE => \N__20087\
        );

    \this_sprites_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34613\,
            RE => \N__20042\,
            WCLKE => \N__29984\,
            WCLK => \N__34614\,
            WE => \N__20086\
        );

    \this_sprites_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34620\,
            RE => \N__20046\,
            WCLKE => \N__28625\,
            WCLK => \N__34621\,
            WE => \N__19986\
        );

    \this_sprites_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_sprites_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_sprites_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_sprites_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_sprites_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_sprites_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34626\,
            RE => \N__19968\,
            WCLKE => \N__28626\,
            WCLK => \N__34627\,
            WE => \N__19975\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__34534\,
            RE => \N__20098\,
            WCLKE => \N__20736\,
            WCLK => \N__34535\,
            WE => \N__19964\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__35920\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35922\,
            DIN => \N__35921\,
            DOUT => \N__35920\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35922\,
            PADOUT => \N__35921\,
            PADIN => \N__35920\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35911\,
            DIN => \N__35910\,
            DOUT => \N__35909\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35911\,
            PADOUT => \N__35910\,
            PADIN => \N__35909\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35902\,
            DIN => \N__35901\,
            DOUT => \N__35900\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35902\,
            PADOUT => \N__35901\,
            PADIN => \N__35900\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35893\,
            DIN => \N__35892\,
            DOUT => \N__35891\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35893\,
            PADOUT => \N__35892\,
            PADIN => \N__35891\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12537\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35884\,
            DIN => \N__35883\,
            DOUT => \N__35882\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35884\,
            PADOUT => \N__35883\,
            PADIN => \N__35882\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12558\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35875\,
            DIN => \N__35874\,
            DOUT => \N__35873\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35875\,
            PADOUT => \N__35874\,
            PADIN => \N__35873\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__20041\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35866\,
            DIN => \N__35865\,
            DOUT => \N__35864\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35866\,
            PADOUT => \N__35865\,
            PADIN => \N__35864\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__17889\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35857\,
            DIN => \N__35856\,
            DOUT => \N__35855\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35857\,
            PADOUT => \N__35856\,
            PADIN => \N__35855\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35848\,
            DIN => \N__35847\,
            DOUT => \N__35846\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35848\,
            PADOUT => \N__35847\,
            PADIN => \N__35846\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35839\,
            DIN => \N__35838\,
            DOUT => \N__35837\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35839\,
            PADOUT => \N__35838\,
            PADIN => \N__35837\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35830\,
            DIN => \N__35829\,
            DOUT => \N__35828\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35830\,
            PADOUT => \N__35829\,
            PADIN => \N__35828\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35821\,
            DIN => \N__35820\,
            DOUT => \N__35819\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35821\,
            PADOUT => \N__35820\,
            PADIN => \N__35819\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35812\,
            DIN => \N__35811\,
            DOUT => \N__35810\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35812\,
            PADOUT => \N__35811\,
            PADIN => \N__35810\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35803\,
            DIN => \N__35802\,
            DOUT => \N__35801\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35803\,
            PADOUT => \N__35802\,
            PADIN => \N__35801\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__33282\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18556\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35794\,
            DIN => \N__35793\,
            DOUT => \N__35792\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35794\,
            PADOUT => \N__35793\,
            PADIN => \N__35792\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__33258\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18643\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35785\,
            DIN => \N__35784\,
            DOUT => \N__35783\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35785\,
            PADOUT => \N__35784\,
            PADIN => \N__35783\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__33231\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18626\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35776\,
            DIN => \N__35775\,
            DOUT => \N__35774\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35776\,
            PADOUT => \N__35775\,
            PADIN => \N__35774\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__33210\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18647\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35767\,
            DIN => \N__35766\,
            DOUT => \N__35765\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35767\,
            PADOUT => \N__35766\,
            PADIN => \N__35765\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__33186\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18613\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35758\,
            DIN => \N__35757\,
            DOUT => \N__35756\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35758\,
            PADOUT => \N__35757\,
            PADIN => \N__35756\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__33165\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18611\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35749\,
            DIN => \N__35748\,
            DOUT => \N__35747\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35749\,
            PADOUT => \N__35748\,
            PADIN => \N__35747\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__34251\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18609\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35740\,
            DIN => \N__35739\,
            DOUT => \N__35738\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35740\,
            PADOUT => \N__35739\,
            PADIN => \N__35738\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__34227\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18641\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35731\,
            DIN => \N__35730\,
            DOUT => \N__35729\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35731\,
            PADOUT => \N__35730\,
            PADIN => \N__35729\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33786\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18597\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35722\,
            DIN => \N__35721\,
            DOUT => \N__35720\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35722\,
            PADOUT => \N__35721\,
            PADIN => \N__35720\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33639\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18648\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35713\,
            DIN => \N__35712\,
            DOUT => \N__35711\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35713\,
            PADOUT => \N__35712\,
            PADIN => \N__35711\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33492\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18636\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35704\,
            DIN => \N__35703\,
            DOUT => \N__35702\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35704\,
            PADOUT => \N__35703\,
            PADIN => \N__35702\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33348\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18612\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35695\,
            DIN => \N__35694\,
            DOUT => \N__35693\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35695\,
            PADOUT => \N__35694\,
            PADIN => \N__35693\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__35337\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18610\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35686\,
            DIN => \N__35685\,
            DOUT => \N__35684\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35686\,
            PADOUT => \N__35685\,
            PADIN => \N__35684\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__35124\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18640\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35677\,
            DIN => \N__35676\,
            DOUT => \N__35675\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35677\,
            PADOUT => \N__35676\,
            PADIN => \N__35675\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__34083\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18596\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35668\,
            DIN => \N__35667\,
            DOUT => \N__35666\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35668\,
            PADOUT => \N__35667\,
            PADIN => \N__35666\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__33939\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18642\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35659\,
            DIN => \N__35658\,
            DOUT => \N__35657\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35659\,
            PADOUT => \N__35658\,
            PADIN => \N__35657\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35650\,
            DIN => \N__35649\,
            DOUT => \N__35648\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35650\,
            PADOUT => \N__35649\,
            PADIN => \N__35648\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35641\,
            DIN => \N__35640\,
            DOUT => \N__35639\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35641\,
            PADOUT => \N__35640\,
            PADIN => \N__35639\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35632\,
            DIN => \N__35631\,
            DOUT => \N__35630\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35632\,
            PADOUT => \N__35631\,
            PADIN => \N__35630\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35623\,
            DIN => \N__35622\,
            DOUT => \N__35621\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35623\,
            PADOUT => \N__35622\,
            PADIN => \N__35621\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35614\,
            DIN => \N__35613\,
            DOUT => \N__35612\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35614\,
            PADOUT => \N__35613\,
            PADIN => \N__35612\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35605\,
            DIN => \N__35604\,
            DOUT => \N__35603\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35605\,
            PADOUT => \N__35604\,
            PADIN => \N__35603\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35596\,
            DIN => \N__35595\,
            DOUT => \N__35594\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35596\,
            PADOUT => \N__35595\,
            PADIN => \N__35594\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35587\,
            DIN => \N__35586\,
            DOUT => \N__35585\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35587\,
            PADOUT => \N__35586\,
            PADIN => \N__35585\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35578\,
            DIN => \N__35577\,
            DOUT => \N__35576\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35578\,
            PADOUT => \N__35577\,
            PADIN => \N__35576\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10992\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35569\,
            DIN => \N__35568\,
            DOUT => \N__35567\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35569\,
            PADOUT => \N__35568\,
            PADIN => \N__35567\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__21400\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35560\,
            DIN => \N__35559\,
            DOUT => \N__35558\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35560\,
            PADOUT => \N__35559\,
            PADIN => \N__35558\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35551\,
            DIN => \N__35550\,
            DOUT => \N__35549\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35551\,
            PADOUT => \N__35550\,
            PADIN => \N__35549\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10932\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35542\,
            DIN => \N__35541\,
            DOUT => \N__35540\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__35542\,
            PADOUT => \N__35541\,
            PADIN => \N__35540\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__19729\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__18590\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35533\,
            DIN => \N__35532\,
            DOUT => \N__35531\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35533\,
            PADOUT => \N__35532\,
            PADIN => \N__35531\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10977\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35524\,
            DIN => \N__35523\,
            DOUT => \N__35522\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35524\,
            PADOUT => \N__35523\,
            PADIN => \N__35522\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11124\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35515\,
            DIN => \N__35514\,
            DOUT => \N__35513\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35515\,
            PADOUT => \N__35514\,
            PADIN => \N__35513\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10962\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35506\,
            DIN => \N__35505\,
            DOUT => \N__35504\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35506\,
            PADOUT => \N__35505\,
            PADIN => \N__35504\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11172\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35497\,
            DIN => \N__35496\,
            DOUT => \N__35495\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35497\,
            PADOUT => \N__35496\,
            PADIN => \N__35495\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10950\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35488\,
            DIN => \N__35487\,
            DOUT => \N__35486\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35488\,
            PADOUT => \N__35487\,
            PADIN => \N__35486\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11145\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35479\,
            DIN => \N__35478\,
            DOUT => \N__35477\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35479\,
            PADOUT => \N__35478\,
            PADIN => \N__35477\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35470\,
            DIN => \N__35469\,
            DOUT => \N__35468\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35470\,
            PADOUT => \N__35469\,
            PADIN => \N__35468\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11154\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35461\,
            DIN => \N__35460\,
            DOUT => \N__35459\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35461\,
            PADOUT => \N__35460\,
            PADIN => \N__35459\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__13956\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__8978\ : InMux
    port map (
            O => \N__35442\,
            I => \un1_M_this_external_address_q_cry_12\
        );

    \I__8977\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35434\
        );

    \I__8976\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35431\
        );

    \I__8975\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35428\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__35434\,
            I => \N__35422\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__35431\,
            I => \N__35417\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__35428\,
            I => \N__35417\
        );

    \I__8971\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35414\
        );

    \I__8970\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35411\
        );

    \I__8969\ : CascadeMux
    port map (
            O => \N__35425\,
            I => \N__35407\
        );

    \I__8968\ : Span4Mux_v
    port map (
            O => \N__35422\,
            I => \N__35403\
        );

    \I__8967\ : Span4Mux_v
    port map (
            O => \N__35417\,
            I => \N__35396\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__35414\,
            I => \N__35396\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__35411\,
            I => \N__35396\
        );

    \I__8964\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35393\
        );

    \I__8963\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35390\
        );

    \I__8962\ : CascadeMux
    port map (
            O => \N__35406\,
            I => \N__35387\
        );

    \I__8961\ : Sp12to4
    port map (
            O => \N__35403\,
            I => \N__35384\
        );

    \I__8960\ : Span4Mux_v
    port map (
            O => \N__35396\,
            I => \N__35380\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__35393\,
            I => \N__35375\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__35390\,
            I => \N__35375\
        );

    \I__8957\ : InMux
    port map (
            O => \N__35387\,
            I => \N__35372\
        );

    \I__8956\ : Span12Mux_h
    port map (
            O => \N__35384\,
            I => \N__35369\
        );

    \I__8955\ : InMux
    port map (
            O => \N__35383\,
            I => \N__35366\
        );

    \I__8954\ : Span4Mux_v
    port map (
            O => \N__35380\,
            I => \N__35359\
        );

    \I__8953\ : Span4Mux_h
    port map (
            O => \N__35375\,
            I => \N__35359\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__35372\,
            I => \N__35359\
        );

    \I__8951\ : Span12Mux_v
    port map (
            O => \N__35369\,
            I => \N__35356\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35353\
        );

    \I__8949\ : Span4Mux_v
    port map (
            O => \N__35359\,
            I => \N__35350\
        );

    \I__8948\ : Span12Mux_h
    port map (
            O => \N__35356\,
            I => \N__35345\
        );

    \I__8947\ : Span12Mux_v
    port map (
            O => \N__35353\,
            I => \N__35345\
        );

    \I__8946\ : Sp12to4
    port map (
            O => \N__35350\,
            I => \N__35342\
        );

    \I__8945\ : Odrv12
    port map (
            O => \N__35345\,
            I => port_data_c_6
        );

    \I__8944\ : Odrv12
    port map (
            O => \N__35342\,
            I => port_data_c_6
        );

    \I__8943\ : IoInMux
    port map (
            O => \N__35337\,
            I => \N__35334\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__35334\,
            I => \N__35330\
        );

    \I__8941\ : CascadeMux
    port map (
            O => \N__35333\,
            I => \N__35327\
        );

    \I__8940\ : Span12Mux_s4_h
    port map (
            O => \N__35330\,
            I => \N__35324\
        );

    \I__8939\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35321\
        );

    \I__8938\ : Odrv12
    port map (
            O => \N__35324\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__35321\,
            I => \M_this_external_address_qZ0Z_14\
        );

    \I__8936\ : InMux
    port map (
            O => \N__35316\,
            I => \un1_M_this_external_address_q_cry_13\
        );

    \I__8935\ : InMux
    port map (
            O => \N__35313\,
            I => \N__35289\
        );

    \I__8934\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35289\
        );

    \I__8933\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35289\
        );

    \I__8932\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35289\
        );

    \I__8931\ : InMux
    port map (
            O => \N__35309\,
            I => \N__35280\
        );

    \I__8930\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35280\
        );

    \I__8929\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35280\
        );

    \I__8928\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35280\
        );

    \I__8927\ : InMux
    port map (
            O => \N__35305\,
            I => \N__35271\
        );

    \I__8926\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35271\
        );

    \I__8925\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35271\
        );

    \I__8924\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35271\
        );

    \I__8923\ : InMux
    port map (
            O => \N__35301\,
            I => \N__35262\
        );

    \I__8922\ : InMux
    port map (
            O => \N__35300\,
            I => \N__35262\
        );

    \I__8921\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35262\
        );

    \I__8920\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35262\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__35289\,
            I => \N__35256\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35256\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35251\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__35262\,
            I => \N__35251\
        );

    \I__8915\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35248\
        );

    \I__8914\ : Span4Mux_v
    port map (
            O => \N__35256\,
            I => \N__35243\
        );

    \I__8913\ : Span4Mux_v
    port map (
            O => \N__35251\,
            I => \N__35243\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__35248\,
            I => \N__35240\
        );

    \I__8911\ : Span4Mux_h
    port map (
            O => \N__35243\,
            I => \N__35237\
        );

    \I__8910\ : Span4Mux_v
    port map (
            O => \N__35240\,
            I => \N__35234\
        );

    \I__8909\ : Span4Mux_h
    port map (
            O => \N__35237\,
            I => \N__35231\
        );

    \I__8908\ : Odrv4
    port map (
            O => \N__35234\,
            I => \N_749_0\
        );

    \I__8907\ : Odrv4
    port map (
            O => \N__35231\,
            I => \N_749_0\
        );

    \I__8906\ : InMux
    port map (
            O => \N__35226\,
            I => \N__35223\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__35223\,
            I => \N__35218\
        );

    \I__8904\ : InMux
    port map (
            O => \N__35222\,
            I => \N__35215\
        );

    \I__8903\ : CascadeMux
    port map (
            O => \N__35221\,
            I => \N__35212\
        );

    \I__8902\ : Span4Mux_v
    port map (
            O => \N__35218\,
            I => \N__35208\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__35215\,
            I => \N__35205\
        );

    \I__8900\ : InMux
    port map (
            O => \N__35212\,
            I => \N__35202\
        );

    \I__8899\ : CascadeMux
    port map (
            O => \N__35211\,
            I => \N__35197\
        );

    \I__8898\ : Span4Mux_h
    port map (
            O => \N__35208\,
            I => \N__35192\
        );

    \I__8897\ : Span4Mux_v
    port map (
            O => \N__35205\,
            I => \N__35192\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__35202\,
            I => \N__35189\
        );

    \I__8895\ : CascadeMux
    port map (
            O => \N__35201\,
            I => \N__35186\
        );

    \I__8894\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35183\
        );

    \I__8893\ : InMux
    port map (
            O => \N__35197\,
            I => \N__35180\
        );

    \I__8892\ : Span4Mux_h
    port map (
            O => \N__35192\,
            I => \N__35175\
        );

    \I__8891\ : Span4Mux_v
    port map (
            O => \N__35189\,
            I => \N__35175\
        );

    \I__8890\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35172\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__35183\,
            I => \N__35169\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__35165\
        );

    \I__8887\ : Sp12to4
    port map (
            O => \N__35175\,
            I => \N__35160\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__35172\,
            I => \N__35160\
        );

    \I__8885\ : Span4Mux_v
    port map (
            O => \N__35169\,
            I => \N__35157\
        );

    \I__8884\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35154\
        );

    \I__8883\ : Span4Mux_v
    port map (
            O => \N__35165\,
            I => \N__35151\
        );

    \I__8882\ : Span12Mux_s6_h
    port map (
            O => \N__35160\,
            I => \N__35148\
        );

    \I__8881\ : Sp12to4
    port map (
            O => \N__35157\,
            I => \N__35143\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__35154\,
            I => \N__35143\
        );

    \I__8879\ : Span4Mux_v
    port map (
            O => \N__35151\,
            I => \N__35140\
        );

    \I__8878\ : Span12Mux_v
    port map (
            O => \N__35148\,
            I => \N__35137\
        );

    \I__8877\ : Span12Mux_v
    port map (
            O => \N__35143\,
            I => \N__35132\
        );

    \I__8876\ : Sp12to4
    port map (
            O => \N__35140\,
            I => \N__35132\
        );

    \I__8875\ : Odrv12
    port map (
            O => \N__35137\,
            I => port_data_c_7
        );

    \I__8874\ : Odrv12
    port map (
            O => \N__35132\,
            I => port_data_c_7
        );

    \I__8873\ : InMux
    port map (
            O => \N__35127\,
            I => \un1_M_this_external_address_q_cry_14\
        );

    \I__8872\ : IoInMux
    port map (
            O => \N__35124\,
            I => \N__35121\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__35118\
        );

    \I__8870\ : Span4Mux_s0_h
    port map (
            O => \N__35118\,
            I => \N__35115\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__35115\,
            I => \N__35112\
        );

    \I__8868\ : Sp12to4
    port map (
            O => \N__35112\,
            I => \N__35109\
        );

    \I__8867\ : Span12Mux_v
    port map (
            O => \N__35109\,
            I => \N__35105\
        );

    \I__8866\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35102\
        );

    \I__8865\ : Odrv12
    port map (
            O => \N__35105\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__35102\,
            I => \M_this_external_address_qZ0Z_15\
        );

    \I__8863\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35065\
        );

    \I__8862\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35065\
        );

    \I__8861\ : InMux
    port map (
            O => \N__35095\,
            I => \N__35058\
        );

    \I__8860\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35058\
        );

    \I__8859\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35058\
        );

    \I__8858\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35055\
        );

    \I__8857\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35050\
        );

    \I__8856\ : InMux
    port map (
            O => \N__35090\,
            I => \N__35050\
        );

    \I__8855\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35047\
        );

    \I__8854\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35044\
        );

    \I__8853\ : InMux
    port map (
            O => \N__35087\,
            I => \N__35041\
        );

    \I__8852\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35038\
        );

    \I__8851\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35033\
        );

    \I__8850\ : InMux
    port map (
            O => \N__35084\,
            I => \N__35033\
        );

    \I__8849\ : InMux
    port map (
            O => \N__35083\,
            I => \N__35030\
        );

    \I__8848\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35027\
        );

    \I__8847\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35024\
        );

    \I__8846\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35019\
        );

    \I__8845\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35019\
        );

    \I__8844\ : InMux
    port map (
            O => \N__35078\,
            I => \N__35014\
        );

    \I__8843\ : InMux
    port map (
            O => \N__35077\,
            I => \N__35014\
        );

    \I__8842\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35011\
        );

    \I__8841\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35008\
        );

    \I__8840\ : InMux
    port map (
            O => \N__35074\,
            I => \N__35001\
        );

    \I__8839\ : InMux
    port map (
            O => \N__35073\,
            I => \N__35001\
        );

    \I__8838\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35001\
        );

    \I__8837\ : InMux
    port map (
            O => \N__35071\,
            I => \N__34996\
        );

    \I__8836\ : InMux
    port map (
            O => \N__35070\,
            I => \N__34996\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__35065\,
            I => \N__34978\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__35058\,
            I => \N__34975\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__35055\,
            I => \N__34972\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__34969\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__35047\,
            I => \N__34966\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__35044\,
            I => \N__34963\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__35041\,
            I => \N__34960\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__35038\,
            I => \N__34957\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__35033\,
            I => \N__34954\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__35030\,
            I => \N__34951\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__35027\,
            I => \N__34948\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__35024\,
            I => \N__34945\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__35019\,
            I => \N__34942\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__35014\,
            I => \N__34939\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__35011\,
            I => \N__34936\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__35008\,
            I => \N__34933\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__35001\,
            I => \N__34930\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__34996\,
            I => \N__34927\
        );

    \I__8817\ : SRMux
    port map (
            O => \N__34995\,
            I => \N__34860\
        );

    \I__8816\ : SRMux
    port map (
            O => \N__34994\,
            I => \N__34860\
        );

    \I__8815\ : SRMux
    port map (
            O => \N__34993\,
            I => \N__34860\
        );

    \I__8814\ : SRMux
    port map (
            O => \N__34992\,
            I => \N__34860\
        );

    \I__8813\ : SRMux
    port map (
            O => \N__34991\,
            I => \N__34860\
        );

    \I__8812\ : SRMux
    port map (
            O => \N__34990\,
            I => \N__34860\
        );

    \I__8811\ : SRMux
    port map (
            O => \N__34989\,
            I => \N__34860\
        );

    \I__8810\ : SRMux
    port map (
            O => \N__34988\,
            I => \N__34860\
        );

    \I__8809\ : SRMux
    port map (
            O => \N__34987\,
            I => \N__34860\
        );

    \I__8808\ : SRMux
    port map (
            O => \N__34986\,
            I => \N__34860\
        );

    \I__8807\ : SRMux
    port map (
            O => \N__34985\,
            I => \N__34860\
        );

    \I__8806\ : SRMux
    port map (
            O => \N__34984\,
            I => \N__34860\
        );

    \I__8805\ : SRMux
    port map (
            O => \N__34983\,
            I => \N__34860\
        );

    \I__8804\ : SRMux
    port map (
            O => \N__34982\,
            I => \N__34860\
        );

    \I__8803\ : SRMux
    port map (
            O => \N__34981\,
            I => \N__34860\
        );

    \I__8802\ : Glb2LocalMux
    port map (
            O => \N__34978\,
            I => \N__34860\
        );

    \I__8801\ : Glb2LocalMux
    port map (
            O => \N__34975\,
            I => \N__34860\
        );

    \I__8800\ : Glb2LocalMux
    port map (
            O => \N__34972\,
            I => \N__34860\
        );

    \I__8799\ : Glb2LocalMux
    port map (
            O => \N__34969\,
            I => \N__34860\
        );

    \I__8798\ : Glb2LocalMux
    port map (
            O => \N__34966\,
            I => \N__34860\
        );

    \I__8797\ : Glb2LocalMux
    port map (
            O => \N__34963\,
            I => \N__34860\
        );

    \I__8796\ : Glb2LocalMux
    port map (
            O => \N__34960\,
            I => \N__34860\
        );

    \I__8795\ : Glb2LocalMux
    port map (
            O => \N__34957\,
            I => \N__34860\
        );

    \I__8794\ : Glb2LocalMux
    port map (
            O => \N__34954\,
            I => \N__34860\
        );

    \I__8793\ : Glb2LocalMux
    port map (
            O => \N__34951\,
            I => \N__34860\
        );

    \I__8792\ : Glb2LocalMux
    port map (
            O => \N__34948\,
            I => \N__34860\
        );

    \I__8791\ : Glb2LocalMux
    port map (
            O => \N__34945\,
            I => \N__34860\
        );

    \I__8790\ : Glb2LocalMux
    port map (
            O => \N__34942\,
            I => \N__34860\
        );

    \I__8789\ : Glb2LocalMux
    port map (
            O => \N__34939\,
            I => \N__34860\
        );

    \I__8788\ : Glb2LocalMux
    port map (
            O => \N__34936\,
            I => \N__34860\
        );

    \I__8787\ : Glb2LocalMux
    port map (
            O => \N__34933\,
            I => \N__34860\
        );

    \I__8786\ : Glb2LocalMux
    port map (
            O => \N__34930\,
            I => \N__34860\
        );

    \I__8785\ : Glb2LocalMux
    port map (
            O => \N__34927\,
            I => \N__34860\
        );

    \I__8784\ : GlobalMux
    port map (
            O => \N__34860\,
            I => \N__34857\
        );

    \I__8783\ : gio2CtrlBuf
    port map (
            O => \N__34857\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__8782\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34851\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__34851\,
            I => \N__34845\
        );

    \I__8780\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34838\
        );

    \I__8779\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34838\
        );

    \I__8778\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34838\
        );

    \I__8777\ : Span4Mux_s3_h
    port map (
            O => \N__34845\,
            I => \N__34832\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__34838\,
            I => \N__34832\
        );

    \I__8775\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34826\
        );

    \I__8774\ : Span4Mux_h
    port map (
            O => \N__34832\,
            I => \N__34823\
        );

    \I__8773\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34820\
        );

    \I__8772\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34817\
        );

    \I__8771\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34813\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34810\
        );

    \I__8769\ : Span4Mux_h
    port map (
            O => \N__34823\,
            I => \N__34803\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34803\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__34817\,
            I => \N__34803\
        );

    \I__8766\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34800\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__34813\,
            I => \N__34797\
        );

    \I__8764\ : Span4Mux_h
    port map (
            O => \N__34810\,
            I => \N__34792\
        );

    \I__8763\ : Span4Mux_h
    port map (
            O => \N__34803\,
            I => \N__34792\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__34800\,
            I => \N__34789\
        );

    \I__8761\ : Span4Mux_h
    port map (
            O => \N__34797\,
            I => \N__34786\
        );

    \I__8760\ : Span4Mux_v
    port map (
            O => \N__34792\,
            I => \N__34781\
        );

    \I__8759\ : Span4Mux_h
    port map (
            O => \N__34789\,
            I => \N__34781\
        );

    \I__8758\ : Span4Mux_v
    port map (
            O => \N__34786\,
            I => \N__34777\
        );

    \I__8757\ : Span4Mux_v
    port map (
            O => \N__34781\,
            I => \N__34774\
        );

    \I__8756\ : InMux
    port map (
            O => \N__34780\,
            I => \N__34771\
        );

    \I__8755\ : Span4Mux_v
    port map (
            O => \N__34777\,
            I => \N__34768\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__34774\,
            I => \N__34765\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34762\
        );

    \I__8752\ : Span4Mux_v
    port map (
            O => \N__34768\,
            I => \N__34759\
        );

    \I__8751\ : Span4Mux_v
    port map (
            O => \N__34765\,
            I => \N__34756\
        );

    \I__8750\ : Span12Mux_v
    port map (
            O => \N__34762\,
            I => \N__34753\
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__34759\,
            I => rst_n_c
        );

    \I__8748\ : Odrv4
    port map (
            O => \N__34756\,
            I => rst_n_c
        );

    \I__8747\ : Odrv12
    port map (
            O => \N__34753\,
            I => rst_n_c
        );

    \I__8746\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34743\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__34743\,
            I => \N__34740\
        );

    \I__8744\ : Span4Mux_s2_h
    port map (
            O => \N__34740\,
            I => \N__34737\
        );

    \I__8743\ : Odrv4
    port map (
            O => \N__34737\,
            I => \this_reset_cond.M_stage_qZ0Z_8\
        );

    \I__8742\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34730\
        );

    \I__8741\ : InMux
    port map (
            O => \N__34733\,
            I => \N__34727\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__34730\,
            I => \N__34716\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__34727\,
            I => \N__34716\
        );

    \I__8738\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34705\
        );

    \I__8737\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34705\
        );

    \I__8736\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34705\
        );

    \I__8735\ : InMux
    port map (
            O => \N__34723\,
            I => \N__34705\
        );

    \I__8734\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34705\
        );

    \I__8733\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34702\
        );

    \I__8732\ : Span4Mux_h
    port map (
            O => \N__34716\,
            I => \N__34696\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__34705\,
            I => \N__34696\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__34702\,
            I => \N__34692\
        );

    \I__8729\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34689\
        );

    \I__8728\ : Span4Mux_v
    port map (
            O => \N__34696\,
            I => \N__34686\
        );

    \I__8727\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34683\
        );

    \I__8726\ : Span4Mux_h
    port map (
            O => \N__34692\,
            I => \N__34678\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__34689\,
            I => \N__34678\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__34686\,
            I => \N__34675\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__34683\,
            I => \N__34672\
        );

    \I__8722\ : Sp12to4
    port map (
            O => \N__34678\,
            I => \N__34669\
        );

    \I__8721\ : Span4Mux_h
    port map (
            O => \N__34675\,
            I => \N__34664\
        );

    \I__8720\ : Span4Mux_v
    port map (
            O => \N__34672\,
            I => \N__34664\
        );

    \I__8719\ : Span12Mux_v
    port map (
            O => \N__34669\,
            I => \N__34661\
        );

    \I__8718\ : Sp12to4
    port map (
            O => \N__34664\,
            I => \N__34658\
        );

    \I__8717\ : Span12Mux_h
    port map (
            O => \N__34661\,
            I => \N__34654\
        );

    \I__8716\ : Span12Mux_h
    port map (
            O => \N__34658\,
            I => \N__34651\
        );

    \I__8715\ : IoInMux
    port map (
            O => \N__34657\,
            I => \N__34648\
        );

    \I__8714\ : Odrv12
    port map (
            O => \N__34654\,
            I => \M_this_reset_cond_out_0\
        );

    \I__8713\ : Odrv12
    port map (
            O => \N__34651\,
            I => \M_this_reset_cond_out_0\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__34648\,
            I => \M_this_reset_cond_out_0\
        );

    \I__8711\ : ClkMux
    port map (
            O => \N__34641\,
            I => \N__34257\
        );

    \I__8710\ : ClkMux
    port map (
            O => \N__34640\,
            I => \N__34257\
        );

    \I__8709\ : ClkMux
    port map (
            O => \N__34639\,
            I => \N__34257\
        );

    \I__8708\ : ClkMux
    port map (
            O => \N__34638\,
            I => \N__34257\
        );

    \I__8707\ : ClkMux
    port map (
            O => \N__34637\,
            I => \N__34257\
        );

    \I__8706\ : ClkMux
    port map (
            O => \N__34636\,
            I => \N__34257\
        );

    \I__8705\ : ClkMux
    port map (
            O => \N__34635\,
            I => \N__34257\
        );

    \I__8704\ : ClkMux
    port map (
            O => \N__34634\,
            I => \N__34257\
        );

    \I__8703\ : ClkMux
    port map (
            O => \N__34633\,
            I => \N__34257\
        );

    \I__8702\ : ClkMux
    port map (
            O => \N__34632\,
            I => \N__34257\
        );

    \I__8701\ : ClkMux
    port map (
            O => \N__34631\,
            I => \N__34257\
        );

    \I__8700\ : ClkMux
    port map (
            O => \N__34630\,
            I => \N__34257\
        );

    \I__8699\ : ClkMux
    port map (
            O => \N__34629\,
            I => \N__34257\
        );

    \I__8698\ : ClkMux
    port map (
            O => \N__34628\,
            I => \N__34257\
        );

    \I__8697\ : ClkMux
    port map (
            O => \N__34627\,
            I => \N__34257\
        );

    \I__8696\ : ClkMux
    port map (
            O => \N__34626\,
            I => \N__34257\
        );

    \I__8695\ : ClkMux
    port map (
            O => \N__34625\,
            I => \N__34257\
        );

    \I__8694\ : ClkMux
    port map (
            O => \N__34624\,
            I => \N__34257\
        );

    \I__8693\ : ClkMux
    port map (
            O => \N__34623\,
            I => \N__34257\
        );

    \I__8692\ : ClkMux
    port map (
            O => \N__34622\,
            I => \N__34257\
        );

    \I__8691\ : ClkMux
    port map (
            O => \N__34621\,
            I => \N__34257\
        );

    \I__8690\ : ClkMux
    port map (
            O => \N__34620\,
            I => \N__34257\
        );

    \I__8689\ : ClkMux
    port map (
            O => \N__34619\,
            I => \N__34257\
        );

    \I__8688\ : ClkMux
    port map (
            O => \N__34618\,
            I => \N__34257\
        );

    \I__8687\ : ClkMux
    port map (
            O => \N__34617\,
            I => \N__34257\
        );

    \I__8686\ : ClkMux
    port map (
            O => \N__34616\,
            I => \N__34257\
        );

    \I__8685\ : ClkMux
    port map (
            O => \N__34615\,
            I => \N__34257\
        );

    \I__8684\ : ClkMux
    port map (
            O => \N__34614\,
            I => \N__34257\
        );

    \I__8683\ : ClkMux
    port map (
            O => \N__34613\,
            I => \N__34257\
        );

    \I__8682\ : ClkMux
    port map (
            O => \N__34612\,
            I => \N__34257\
        );

    \I__8681\ : ClkMux
    port map (
            O => \N__34611\,
            I => \N__34257\
        );

    \I__8680\ : ClkMux
    port map (
            O => \N__34610\,
            I => \N__34257\
        );

    \I__8679\ : ClkMux
    port map (
            O => \N__34609\,
            I => \N__34257\
        );

    \I__8678\ : ClkMux
    port map (
            O => \N__34608\,
            I => \N__34257\
        );

    \I__8677\ : ClkMux
    port map (
            O => \N__34607\,
            I => \N__34257\
        );

    \I__8676\ : ClkMux
    port map (
            O => \N__34606\,
            I => \N__34257\
        );

    \I__8675\ : ClkMux
    port map (
            O => \N__34605\,
            I => \N__34257\
        );

    \I__8674\ : ClkMux
    port map (
            O => \N__34604\,
            I => \N__34257\
        );

    \I__8673\ : ClkMux
    port map (
            O => \N__34603\,
            I => \N__34257\
        );

    \I__8672\ : ClkMux
    port map (
            O => \N__34602\,
            I => \N__34257\
        );

    \I__8671\ : ClkMux
    port map (
            O => \N__34601\,
            I => \N__34257\
        );

    \I__8670\ : ClkMux
    port map (
            O => \N__34600\,
            I => \N__34257\
        );

    \I__8669\ : ClkMux
    port map (
            O => \N__34599\,
            I => \N__34257\
        );

    \I__8668\ : ClkMux
    port map (
            O => \N__34598\,
            I => \N__34257\
        );

    \I__8667\ : ClkMux
    port map (
            O => \N__34597\,
            I => \N__34257\
        );

    \I__8666\ : ClkMux
    port map (
            O => \N__34596\,
            I => \N__34257\
        );

    \I__8665\ : ClkMux
    port map (
            O => \N__34595\,
            I => \N__34257\
        );

    \I__8664\ : ClkMux
    port map (
            O => \N__34594\,
            I => \N__34257\
        );

    \I__8663\ : ClkMux
    port map (
            O => \N__34593\,
            I => \N__34257\
        );

    \I__8662\ : ClkMux
    port map (
            O => \N__34592\,
            I => \N__34257\
        );

    \I__8661\ : ClkMux
    port map (
            O => \N__34591\,
            I => \N__34257\
        );

    \I__8660\ : ClkMux
    port map (
            O => \N__34590\,
            I => \N__34257\
        );

    \I__8659\ : ClkMux
    port map (
            O => \N__34589\,
            I => \N__34257\
        );

    \I__8658\ : ClkMux
    port map (
            O => \N__34588\,
            I => \N__34257\
        );

    \I__8657\ : ClkMux
    port map (
            O => \N__34587\,
            I => \N__34257\
        );

    \I__8656\ : ClkMux
    port map (
            O => \N__34586\,
            I => \N__34257\
        );

    \I__8655\ : ClkMux
    port map (
            O => \N__34585\,
            I => \N__34257\
        );

    \I__8654\ : ClkMux
    port map (
            O => \N__34584\,
            I => \N__34257\
        );

    \I__8653\ : ClkMux
    port map (
            O => \N__34583\,
            I => \N__34257\
        );

    \I__8652\ : ClkMux
    port map (
            O => \N__34582\,
            I => \N__34257\
        );

    \I__8651\ : ClkMux
    port map (
            O => \N__34581\,
            I => \N__34257\
        );

    \I__8650\ : ClkMux
    port map (
            O => \N__34580\,
            I => \N__34257\
        );

    \I__8649\ : ClkMux
    port map (
            O => \N__34579\,
            I => \N__34257\
        );

    \I__8648\ : ClkMux
    port map (
            O => \N__34578\,
            I => \N__34257\
        );

    \I__8647\ : ClkMux
    port map (
            O => \N__34577\,
            I => \N__34257\
        );

    \I__8646\ : ClkMux
    port map (
            O => \N__34576\,
            I => \N__34257\
        );

    \I__8645\ : ClkMux
    port map (
            O => \N__34575\,
            I => \N__34257\
        );

    \I__8644\ : ClkMux
    port map (
            O => \N__34574\,
            I => \N__34257\
        );

    \I__8643\ : ClkMux
    port map (
            O => \N__34573\,
            I => \N__34257\
        );

    \I__8642\ : ClkMux
    port map (
            O => \N__34572\,
            I => \N__34257\
        );

    \I__8641\ : ClkMux
    port map (
            O => \N__34571\,
            I => \N__34257\
        );

    \I__8640\ : ClkMux
    port map (
            O => \N__34570\,
            I => \N__34257\
        );

    \I__8639\ : ClkMux
    port map (
            O => \N__34569\,
            I => \N__34257\
        );

    \I__8638\ : ClkMux
    port map (
            O => \N__34568\,
            I => \N__34257\
        );

    \I__8637\ : ClkMux
    port map (
            O => \N__34567\,
            I => \N__34257\
        );

    \I__8636\ : ClkMux
    port map (
            O => \N__34566\,
            I => \N__34257\
        );

    \I__8635\ : ClkMux
    port map (
            O => \N__34565\,
            I => \N__34257\
        );

    \I__8634\ : ClkMux
    port map (
            O => \N__34564\,
            I => \N__34257\
        );

    \I__8633\ : ClkMux
    port map (
            O => \N__34563\,
            I => \N__34257\
        );

    \I__8632\ : ClkMux
    port map (
            O => \N__34562\,
            I => \N__34257\
        );

    \I__8631\ : ClkMux
    port map (
            O => \N__34561\,
            I => \N__34257\
        );

    \I__8630\ : ClkMux
    port map (
            O => \N__34560\,
            I => \N__34257\
        );

    \I__8629\ : ClkMux
    port map (
            O => \N__34559\,
            I => \N__34257\
        );

    \I__8628\ : ClkMux
    port map (
            O => \N__34558\,
            I => \N__34257\
        );

    \I__8627\ : ClkMux
    port map (
            O => \N__34557\,
            I => \N__34257\
        );

    \I__8626\ : ClkMux
    port map (
            O => \N__34556\,
            I => \N__34257\
        );

    \I__8625\ : ClkMux
    port map (
            O => \N__34555\,
            I => \N__34257\
        );

    \I__8624\ : ClkMux
    port map (
            O => \N__34554\,
            I => \N__34257\
        );

    \I__8623\ : ClkMux
    port map (
            O => \N__34553\,
            I => \N__34257\
        );

    \I__8622\ : ClkMux
    port map (
            O => \N__34552\,
            I => \N__34257\
        );

    \I__8621\ : ClkMux
    port map (
            O => \N__34551\,
            I => \N__34257\
        );

    \I__8620\ : ClkMux
    port map (
            O => \N__34550\,
            I => \N__34257\
        );

    \I__8619\ : ClkMux
    port map (
            O => \N__34549\,
            I => \N__34257\
        );

    \I__8618\ : ClkMux
    port map (
            O => \N__34548\,
            I => \N__34257\
        );

    \I__8617\ : ClkMux
    port map (
            O => \N__34547\,
            I => \N__34257\
        );

    \I__8616\ : ClkMux
    port map (
            O => \N__34546\,
            I => \N__34257\
        );

    \I__8615\ : ClkMux
    port map (
            O => \N__34545\,
            I => \N__34257\
        );

    \I__8614\ : ClkMux
    port map (
            O => \N__34544\,
            I => \N__34257\
        );

    \I__8613\ : ClkMux
    port map (
            O => \N__34543\,
            I => \N__34257\
        );

    \I__8612\ : ClkMux
    port map (
            O => \N__34542\,
            I => \N__34257\
        );

    \I__8611\ : ClkMux
    port map (
            O => \N__34541\,
            I => \N__34257\
        );

    \I__8610\ : ClkMux
    port map (
            O => \N__34540\,
            I => \N__34257\
        );

    \I__8609\ : ClkMux
    port map (
            O => \N__34539\,
            I => \N__34257\
        );

    \I__8608\ : ClkMux
    port map (
            O => \N__34538\,
            I => \N__34257\
        );

    \I__8607\ : ClkMux
    port map (
            O => \N__34537\,
            I => \N__34257\
        );

    \I__8606\ : ClkMux
    port map (
            O => \N__34536\,
            I => \N__34257\
        );

    \I__8605\ : ClkMux
    port map (
            O => \N__34535\,
            I => \N__34257\
        );

    \I__8604\ : ClkMux
    port map (
            O => \N__34534\,
            I => \N__34257\
        );

    \I__8603\ : ClkMux
    port map (
            O => \N__34533\,
            I => \N__34257\
        );

    \I__8602\ : ClkMux
    port map (
            O => \N__34532\,
            I => \N__34257\
        );

    \I__8601\ : ClkMux
    port map (
            O => \N__34531\,
            I => \N__34257\
        );

    \I__8600\ : ClkMux
    port map (
            O => \N__34530\,
            I => \N__34257\
        );

    \I__8599\ : ClkMux
    port map (
            O => \N__34529\,
            I => \N__34257\
        );

    \I__8598\ : ClkMux
    port map (
            O => \N__34528\,
            I => \N__34257\
        );

    \I__8597\ : ClkMux
    port map (
            O => \N__34527\,
            I => \N__34257\
        );

    \I__8596\ : ClkMux
    port map (
            O => \N__34526\,
            I => \N__34257\
        );

    \I__8595\ : ClkMux
    port map (
            O => \N__34525\,
            I => \N__34257\
        );

    \I__8594\ : ClkMux
    port map (
            O => \N__34524\,
            I => \N__34257\
        );

    \I__8593\ : ClkMux
    port map (
            O => \N__34523\,
            I => \N__34257\
        );

    \I__8592\ : ClkMux
    port map (
            O => \N__34522\,
            I => \N__34257\
        );

    \I__8591\ : ClkMux
    port map (
            O => \N__34521\,
            I => \N__34257\
        );

    \I__8590\ : ClkMux
    port map (
            O => \N__34520\,
            I => \N__34257\
        );

    \I__8589\ : ClkMux
    port map (
            O => \N__34519\,
            I => \N__34257\
        );

    \I__8588\ : ClkMux
    port map (
            O => \N__34518\,
            I => \N__34257\
        );

    \I__8587\ : ClkMux
    port map (
            O => \N__34517\,
            I => \N__34257\
        );

    \I__8586\ : ClkMux
    port map (
            O => \N__34516\,
            I => \N__34257\
        );

    \I__8585\ : ClkMux
    port map (
            O => \N__34515\,
            I => \N__34257\
        );

    \I__8584\ : ClkMux
    port map (
            O => \N__34514\,
            I => \N__34257\
        );

    \I__8583\ : GlobalMux
    port map (
            O => \N__34257\,
            I => \N__34254\
        );

    \I__8582\ : gio2CtrlBuf
    port map (
            O => \N__34254\,
            I => clk_0_c_g
        );

    \I__8581\ : IoInMux
    port map (
            O => \N__34251\,
            I => \N__34248\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__34248\,
            I => \N__34245\
        );

    \I__8579\ : Span4Mux_s1_h
    port map (
            O => \N__34245\,
            I => \N__34242\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__34242\,
            I => \N__34238\
        );

    \I__8577\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34235\
        );

    \I__8576\ : Odrv4
    port map (
            O => \N__34238\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__34235\,
            I => \M_this_external_address_qZ0Z_6\
        );

    \I__8574\ : InMux
    port map (
            O => \N__34230\,
            I => \un1_M_this_external_address_q_cry_5\
        );

    \I__8573\ : IoInMux
    port map (
            O => \N__34227\,
            I => \N__34224\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__8571\ : Span4Mux_s0_h
    port map (
            O => \N__34221\,
            I => \N__34218\
        );

    \I__8570\ : Span4Mux_h
    port map (
            O => \N__34218\,
            I => \N__34215\
        );

    \I__8569\ : Sp12to4
    port map (
            O => \N__34215\,
            I => \N__34212\
        );

    \I__8568\ : Span12Mux_v
    port map (
            O => \N__34212\,
            I => \N__34208\
        );

    \I__8567\ : InMux
    port map (
            O => \N__34211\,
            I => \N__34205\
        );

    \I__8566\ : Odrv12
    port map (
            O => \N__34208\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__34205\,
            I => \M_this_external_address_qZ0Z_7\
        );

    \I__8564\ : InMux
    port map (
            O => \N__34200\,
            I => \un1_M_this_external_address_q_cry_6\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__8562\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34188\
        );

    \I__8561\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34185\
        );

    \I__8560\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34182\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__34191\,
            I => \N__34179\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__34188\,
            I => \N__34174\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__34185\,
            I => \N__34174\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__34182\,
            I => \N__34170\
        );

    \I__8555\ : InMux
    port map (
            O => \N__34179\,
            I => \N__34167\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__34174\,
            I => \N__34163\
        );

    \I__8553\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34160\
        );

    \I__8552\ : Span4Mux_v
    port map (
            O => \N__34170\,
            I => \N__34155\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34152\
        );

    \I__8550\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34149\
        );

    \I__8549\ : Span4Mux_h
    port map (
            O => \N__34163\,
            I => \N__34144\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__34160\,
            I => \N__34144\
        );

    \I__8547\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34141\
        );

    \I__8546\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34138\
        );

    \I__8545\ : Span4Mux_h
    port map (
            O => \N__34155\,
            I => \N__34133\
        );

    \I__8544\ : Span4Mux_v
    port map (
            O => \N__34152\,
            I => \N__34133\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__34149\,
            I => \N__34130\
        );

    \I__8542\ : Span4Mux_v
    port map (
            O => \N__34144\,
            I => \N__34127\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__34141\,
            I => \N__34124\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34120\
        );

    \I__8539\ : Span4Mux_h
    port map (
            O => \N__34133\,
            I => \N__34117\
        );

    \I__8538\ : Span4Mux_v
    port map (
            O => \N__34130\,
            I => \N__34110\
        );

    \I__8537\ : Span4Mux_v
    port map (
            O => \N__34127\,
            I => \N__34110\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__34124\,
            I => \N__34110\
        );

    \I__8535\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34107\
        );

    \I__8534\ : Span4Mux_v
    port map (
            O => \N__34120\,
            I => \N__34104\
        );

    \I__8533\ : Sp12to4
    port map (
            O => \N__34117\,
            I => \N__34097\
        );

    \I__8532\ : Sp12to4
    port map (
            O => \N__34110\,
            I => \N__34097\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__34107\,
            I => \N__34097\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__34104\,
            I => \N__34094\
        );

    \I__8529\ : Span12Mux_h
    port map (
            O => \N__34097\,
            I => \N__34091\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__34094\,
            I => \N__34088\
        );

    \I__8527\ : Odrv12
    port map (
            O => \N__34091\,
            I => port_data_c_0
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__34088\,
            I => port_data_c_0
        );

    \I__8525\ : IoInMux
    port map (
            O => \N__34083\,
            I => \N__34080\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__34080\,
            I => \N__34077\
        );

    \I__8523\ : Span4Mux_s2_v
    port map (
            O => \N__34077\,
            I => \N__34074\
        );

    \I__8522\ : Sp12to4
    port map (
            O => \N__34074\,
            I => \N__34071\
        );

    \I__8521\ : Span12Mux_v
    port map (
            O => \N__34071\,
            I => \N__34067\
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__34070\,
            I => \N__34064\
        );

    \I__8519\ : Span12Mux_h
    port map (
            O => \N__34067\,
            I => \N__34061\
        );

    \I__8518\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34058\
        );

    \I__8517\ : Odrv12
    port map (
            O => \N__34061\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__34058\,
            I => \M_this_external_address_qZ0Z_8\
        );

    \I__8515\ : InMux
    port map (
            O => \N__34053\,
            I => \bfn_28_22_0_\
        );

    \I__8514\ : CascadeMux
    port map (
            O => \N__34050\,
            I => \N__34047\
        );

    \I__8513\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34043\
        );

    \I__8512\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34038\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__34043\,
            I => \N__34033\
        );

    \I__8510\ : InMux
    port map (
            O => \N__34042\,
            I => \N__34030\
        );

    \I__8509\ : CascadeMux
    port map (
            O => \N__34041\,
            I => \N__34027\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__34038\,
            I => \N__34024\
        );

    \I__8507\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34021\
        );

    \I__8506\ : CascadeMux
    port map (
            O => \N__34036\,
            I => \N__34017\
        );

    \I__8505\ : Span4Mux_v
    port map (
            O => \N__34033\,
            I => \N__34011\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__34030\,
            I => \N__34011\
        );

    \I__8503\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34008\
        );

    \I__8502\ : Span4Mux_v
    port map (
            O => \N__34024\,
            I => \N__34005\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__34021\,
            I => \N__34002\
        );

    \I__8500\ : InMux
    port map (
            O => \N__34020\,
            I => \N__33999\
        );

    \I__8499\ : InMux
    port map (
            O => \N__34017\,
            I => \N__33996\
        );

    \I__8498\ : InMux
    port map (
            O => \N__34016\,
            I => \N__33993\
        );

    \I__8497\ : Span4Mux_v
    port map (
            O => \N__34011\,
            I => \N__33990\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__33987\
        );

    \I__8495\ : Span4Mux_h
    port map (
            O => \N__34005\,
            I => \N__33980\
        );

    \I__8494\ : Span4Mux_v
    port map (
            O => \N__34002\,
            I => \N__33980\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__33999\,
            I => \N__33980\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__33996\,
            I => \N__33974\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__33993\,
            I => \N__33974\
        );

    \I__8490\ : Span4Mux_v
    port map (
            O => \N__33990\,
            I => \N__33971\
        );

    \I__8489\ : Span4Mux_v
    port map (
            O => \N__33987\,
            I => \N__33966\
        );

    \I__8488\ : Span4Mux_v
    port map (
            O => \N__33980\,
            I => \N__33966\
        );

    \I__8487\ : InMux
    port map (
            O => \N__33979\,
            I => \N__33963\
        );

    \I__8486\ : Span12Mux_h
    port map (
            O => \N__33974\,
            I => \N__33960\
        );

    \I__8485\ : Sp12to4
    port map (
            O => \N__33971\,
            I => \N__33955\
        );

    \I__8484\ : Sp12to4
    port map (
            O => \N__33966\,
            I => \N__33955\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__33963\,
            I => \N__33952\
        );

    \I__8482\ : Span12Mux_v
    port map (
            O => \N__33960\,
            I => \N__33947\
        );

    \I__8481\ : Span12Mux_h
    port map (
            O => \N__33955\,
            I => \N__33947\
        );

    \I__8480\ : Sp12to4
    port map (
            O => \N__33952\,
            I => \N__33944\
        );

    \I__8479\ : Odrv12
    port map (
            O => \N__33947\,
            I => port_data_c_1
        );

    \I__8478\ : Odrv12
    port map (
            O => \N__33944\,
            I => port_data_c_1
        );

    \I__8477\ : IoInMux
    port map (
            O => \N__33939\,
            I => \N__33936\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__33936\,
            I => \N__33933\
        );

    \I__8475\ : IoSpan4Mux
    port map (
            O => \N__33933\,
            I => \N__33930\
        );

    \I__8474\ : Span4Mux_s2_v
    port map (
            O => \N__33930\,
            I => \N__33926\
        );

    \I__8473\ : CascadeMux
    port map (
            O => \N__33929\,
            I => \N__33923\
        );

    \I__8472\ : Sp12to4
    port map (
            O => \N__33926\,
            I => \N__33920\
        );

    \I__8471\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33917\
        );

    \I__8470\ : Odrv12
    port map (
            O => \N__33920\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__33917\,
            I => \M_this_external_address_qZ0Z_9\
        );

    \I__8468\ : InMux
    port map (
            O => \N__33912\,
            I => \un1_M_this_external_address_q_cry_8\
        );

    \I__8467\ : CascadeMux
    port map (
            O => \N__33909\,
            I => \N__33905\
        );

    \I__8466\ : CascadeMux
    port map (
            O => \N__33908\,
            I => \N__33901\
        );

    \I__8465\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33898\
        );

    \I__8464\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33893\
        );

    \I__8463\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33889\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33886\
        );

    \I__8461\ : InMux
    port map (
            O => \N__33897\,
            I => \N__33883\
        );

    \I__8460\ : CascadeMux
    port map (
            O => \N__33896\,
            I => \N__33880\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__33893\,
            I => \N__33876\
        );

    \I__8458\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33873\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__33889\,
            I => \N__33870\
        );

    \I__8456\ : Span4Mux_v
    port map (
            O => \N__33886\,
            I => \N__33865\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__33883\,
            I => \N__33865\
        );

    \I__8454\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33862\
        );

    \I__8453\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33859\
        );

    \I__8452\ : Span4Mux_v
    port map (
            O => \N__33876\,
            I => \N__33854\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__33873\,
            I => \N__33854\
        );

    \I__8450\ : Span4Mux_h
    port map (
            O => \N__33870\,
            I => \N__33851\
        );

    \I__8449\ : Span4Mux_v
    port map (
            O => \N__33865\,
            I => \N__33846\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__33862\,
            I => \N__33846\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__33859\,
            I => \N__33841\
        );

    \I__8446\ : Span4Mux_v
    port map (
            O => \N__33854\,
            I => \N__33838\
        );

    \I__8445\ : Span4Mux_h
    port map (
            O => \N__33851\,
            I => \N__33835\
        );

    \I__8444\ : Span4Mux_v
    port map (
            O => \N__33846\,
            I => \N__33832\
        );

    \I__8443\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33829\
        );

    \I__8442\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33826\
        );

    \I__8441\ : Span4Mux_v
    port map (
            O => \N__33841\,
            I => \N__33823\
        );

    \I__8440\ : Sp12to4
    port map (
            O => \N__33838\,
            I => \N__33820\
        );

    \I__8439\ : Sp12to4
    port map (
            O => \N__33835\,
            I => \N__33817\
        );

    \I__8438\ : Span4Mux_h
    port map (
            O => \N__33832\,
            I => \N__33814\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__33829\,
            I => \N__33809\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__33826\,
            I => \N__33809\
        );

    \I__8435\ : Span4Mux_v
    port map (
            O => \N__33823\,
            I => \N__33806\
        );

    \I__8434\ : Span12Mux_h
    port map (
            O => \N__33820\,
            I => \N__33803\
        );

    \I__8433\ : Span12Mux_v
    port map (
            O => \N__33817\,
            I => \N__33796\
        );

    \I__8432\ : Sp12to4
    port map (
            O => \N__33814\,
            I => \N__33796\
        );

    \I__8431\ : Span12Mux_h
    port map (
            O => \N__33809\,
            I => \N__33796\
        );

    \I__8430\ : IoSpan4Mux
    port map (
            O => \N__33806\,
            I => \N__33793\
        );

    \I__8429\ : Odrv12
    port map (
            O => \N__33803\,
            I => port_data_c_2
        );

    \I__8428\ : Odrv12
    port map (
            O => \N__33796\,
            I => port_data_c_2
        );

    \I__8427\ : Odrv4
    port map (
            O => \N__33793\,
            I => port_data_c_2
        );

    \I__8426\ : IoInMux
    port map (
            O => \N__33786\,
            I => \N__33783\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__33783\,
            I => \N__33780\
        );

    \I__8424\ : Span4Mux_s3_v
    port map (
            O => \N__33780\,
            I => \N__33777\
        );

    \I__8423\ : Span4Mux_h
    port map (
            O => \N__33777\,
            I => \N__33774\
        );

    \I__8422\ : Span4Mux_h
    port map (
            O => \N__33774\,
            I => \N__33770\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__33773\,
            I => \N__33767\
        );

    \I__8420\ : Span4Mux_v
    port map (
            O => \N__33770\,
            I => \N__33764\
        );

    \I__8419\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33761\
        );

    \I__8418\ : Odrv4
    port map (
            O => \N__33764\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__33761\,
            I => \M_this_external_address_qZ0Z_10\
        );

    \I__8416\ : InMux
    port map (
            O => \N__33756\,
            I => \un1_M_this_external_address_q_cry_9\
        );

    \I__8415\ : CascadeMux
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__8414\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33746\
        );

    \I__8413\ : CascadeMux
    port map (
            O => \N__33749\,
            I => \N__33743\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33739\
        );

    \I__8411\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33736\
        );

    \I__8410\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33733\
        );

    \I__8409\ : Span4Mux_v
    port map (
            O => \N__33739\,
            I => \N__33725\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__33736\,
            I => \N__33725\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__33733\,
            I => \N__33722\
        );

    \I__8406\ : InMux
    port map (
            O => \N__33732\,
            I => \N__33719\
        );

    \I__8405\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33715\
        );

    \I__8404\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33712\
        );

    \I__8403\ : Span4Mux_h
    port map (
            O => \N__33725\,
            I => \N__33705\
        );

    \I__8402\ : Span4Mux_v
    port map (
            O => \N__33722\,
            I => \N__33705\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33705\
        );

    \I__8400\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33702\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__33715\,
            I => \N__33698\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__33712\,
            I => \N__33694\
        );

    \I__8397\ : Span4Mux_v
    port map (
            O => \N__33705\,
            I => \N__33691\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__33702\,
            I => \N__33688\
        );

    \I__8395\ : CascadeMux
    port map (
            O => \N__33701\,
            I => \N__33685\
        );

    \I__8394\ : Span4Mux_h
    port map (
            O => \N__33698\,
            I => \N__33682\
        );

    \I__8393\ : InMux
    port map (
            O => \N__33697\,
            I => \N__33679\
        );

    \I__8392\ : Span4Mux_v
    port map (
            O => \N__33694\,
            I => \N__33676\
        );

    \I__8391\ : Span4Mux_v
    port map (
            O => \N__33691\,
            I => \N__33673\
        );

    \I__8390\ : Span4Mux_v
    port map (
            O => \N__33688\,
            I => \N__33670\
        );

    \I__8389\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33667\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__33682\,
            I => \N__33662\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__33679\,
            I => \N__33662\
        );

    \I__8386\ : Sp12to4
    port map (
            O => \N__33676\,
            I => \N__33653\
        );

    \I__8385\ : Sp12to4
    port map (
            O => \N__33673\,
            I => \N__33653\
        );

    \I__8384\ : Sp12to4
    port map (
            O => \N__33670\,
            I => \N__33653\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__33667\,
            I => \N__33653\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__33662\,
            I => \N__33650\
        );

    \I__8381\ : Span12Mux_h
    port map (
            O => \N__33653\,
            I => \N__33647\
        );

    \I__8380\ : Span4Mux_v
    port map (
            O => \N__33650\,
            I => \N__33644\
        );

    \I__8379\ : Odrv12
    port map (
            O => \N__33647\,
            I => port_data_c_3
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__33644\,
            I => port_data_c_3
        );

    \I__8377\ : IoInMux
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__33636\,
            I => \N__33633\
        );

    \I__8375\ : IoSpan4Mux
    port map (
            O => \N__33633\,
            I => \N__33630\
        );

    \I__8374\ : Span4Mux_s3_v
    port map (
            O => \N__33630\,
            I => \N__33626\
        );

    \I__8373\ : CascadeMux
    port map (
            O => \N__33629\,
            I => \N__33623\
        );

    \I__8372\ : Span4Mux_v
    port map (
            O => \N__33626\,
            I => \N__33620\
        );

    \I__8371\ : InMux
    port map (
            O => \N__33623\,
            I => \N__33617\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__33620\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__33617\,
            I => \M_this_external_address_qZ0Z_11\
        );

    \I__8368\ : InMux
    port map (
            O => \N__33612\,
            I => \un1_M_this_external_address_q_cry_10\
        );

    \I__8367\ : CascadeMux
    port map (
            O => \N__33609\,
            I => \N__33601\
        );

    \I__8366\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33598\
        );

    \I__8365\ : CascadeMux
    port map (
            O => \N__33607\,
            I => \N__33595\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__33606\,
            I => \N__33592\
        );

    \I__8363\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33589\
        );

    \I__8362\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33586\
        );

    \I__8361\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33581\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__33598\,
            I => \N__33578\
        );

    \I__8359\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33575\
        );

    \I__8358\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33571\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33568\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33565\
        );

    \I__8355\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33562\
        );

    \I__8354\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33559\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__33581\,
            I => \N__33556\
        );

    \I__8352\ : Span4Mux_h
    port map (
            O => \N__33578\,
            I => \N__33553\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__33575\,
            I => \N__33550\
        );

    \I__8350\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33547\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__33571\,
            I => \N__33544\
        );

    \I__8348\ : Span4Mux_v
    port map (
            O => \N__33568\,
            I => \N__33537\
        );

    \I__8347\ : Span4Mux_h
    port map (
            O => \N__33565\,
            I => \N__33537\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__33562\,
            I => \N__33537\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__33559\,
            I => \N__33534\
        );

    \I__8344\ : Span12Mux_h
    port map (
            O => \N__33556\,
            I => \N__33531\
        );

    \I__8343\ : Sp12to4
    port map (
            O => \N__33553\,
            I => \N__33526\
        );

    \I__8342\ : Span12Mux_v
    port map (
            O => \N__33550\,
            I => \N__33526\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__33547\,
            I => \N__33523\
        );

    \I__8340\ : Span4Mux_v
    port map (
            O => \N__33544\,
            I => \N__33520\
        );

    \I__8339\ : Span4Mux_v
    port map (
            O => \N__33537\,
            I => \N__33517\
        );

    \I__8338\ : Span4Mux_v
    port map (
            O => \N__33534\,
            I => \N__33514\
        );

    \I__8337\ : Span12Mux_v
    port map (
            O => \N__33531\,
            I => \N__33511\
        );

    \I__8336\ : Span12Mux_v
    port map (
            O => \N__33526\,
            I => \N__33502\
        );

    \I__8335\ : Span12Mux_h
    port map (
            O => \N__33523\,
            I => \N__33502\
        );

    \I__8334\ : Sp12to4
    port map (
            O => \N__33520\,
            I => \N__33502\
        );

    \I__8333\ : Sp12to4
    port map (
            O => \N__33517\,
            I => \N__33502\
        );

    \I__8332\ : Span4Mux_v
    port map (
            O => \N__33514\,
            I => \N__33499\
        );

    \I__8331\ : Odrv12
    port map (
            O => \N__33511\,
            I => port_data_c_4
        );

    \I__8330\ : Odrv12
    port map (
            O => \N__33502\,
            I => port_data_c_4
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__33499\,
            I => port_data_c_4
        );

    \I__8328\ : IoInMux
    port map (
            O => \N__33492\,
            I => \N__33489\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__33489\,
            I => \N__33485\
        );

    \I__8326\ : CascadeMux
    port map (
            O => \N__33488\,
            I => \N__33482\
        );

    \I__8325\ : Span4Mux_s3_h
    port map (
            O => \N__33485\,
            I => \N__33479\
        );

    \I__8324\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33476\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__33479\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__33476\,
            I => \M_this_external_address_qZ0Z_12\
        );

    \I__8321\ : InMux
    port map (
            O => \N__33471\,
            I => \un1_M_this_external_address_q_cry_11\
        );

    \I__8320\ : CascadeMux
    port map (
            O => \N__33468\,
            I => \N__33464\
        );

    \I__8319\ : CascadeMux
    port map (
            O => \N__33467\,
            I => \N__33460\
        );

    \I__8318\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33454\
        );

    \I__8317\ : InMux
    port map (
            O => \N__33463\,
            I => \N__33451\
        );

    \I__8316\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33448\
        );

    \I__8315\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33444\
        );

    \I__8314\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33441\
        );

    \I__8313\ : CascadeMux
    port map (
            O => \N__33457\,
            I => \N__33438\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__33454\,
            I => \N__33435\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__33451\,
            I => \N__33432\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__33448\,
            I => \N__33429\
        );

    \I__8309\ : InMux
    port map (
            O => \N__33447\,
            I => \N__33426\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__33444\,
            I => \N__33423\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__33441\,
            I => \N__33420\
        );

    \I__8306\ : InMux
    port map (
            O => \N__33438\,
            I => \N__33417\
        );

    \I__8305\ : Span4Mux_v
    port map (
            O => \N__33435\,
            I => \N__33413\
        );

    \I__8304\ : Span4Mux_h
    port map (
            O => \N__33432\,
            I => \N__33406\
        );

    \I__8303\ : Span4Mux_v
    port map (
            O => \N__33429\,
            I => \N__33406\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33406\
        );

    \I__8301\ : Sp12to4
    port map (
            O => \N__33423\,
            I => \N__33402\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__33420\,
            I => \N__33399\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__33417\,
            I => \N__33396\
        );

    \I__8298\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33393\
        );

    \I__8297\ : Span4Mux_v
    port map (
            O => \N__33413\,
            I => \N__33388\
        );

    \I__8296\ : Span4Mux_v
    port map (
            O => \N__33406\,
            I => \N__33388\
        );

    \I__8295\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33385\
        );

    \I__8294\ : Span12Mux_v
    port map (
            O => \N__33402\,
            I => \N__33382\
        );

    \I__8293\ : Span4Mux_v
    port map (
            O => \N__33399\,
            I => \N__33377\
        );

    \I__8292\ : Span4Mux_v
    port map (
            O => \N__33396\,
            I => \N__33377\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__33393\,
            I => \N__33374\
        );

    \I__8290\ : Span4Mux_h
    port map (
            O => \N__33388\,
            I => \N__33371\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__33385\,
            I => \N__33368\
        );

    \I__8288\ : Span12Mux_h
    port map (
            O => \N__33382\,
            I => \N__33361\
        );

    \I__8287\ : Sp12to4
    port map (
            O => \N__33377\,
            I => \N__33361\
        );

    \I__8286\ : Span12Mux_v
    port map (
            O => \N__33374\,
            I => \N__33361\
        );

    \I__8285\ : Span4Mux_h
    port map (
            O => \N__33371\,
            I => \N__33358\
        );

    \I__8284\ : Span4Mux_v
    port map (
            O => \N__33368\,
            I => \N__33355\
        );

    \I__8283\ : Odrv12
    port map (
            O => \N__33361\,
            I => port_data_c_5
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__33358\,
            I => port_data_c_5
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__33355\,
            I => port_data_c_5
        );

    \I__8280\ : IoInMux
    port map (
            O => \N__33348\,
            I => \N__33345\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__33345\,
            I => \N__33341\
        );

    \I__8278\ : CascadeMux
    port map (
            O => \N__33344\,
            I => \N__33338\
        );

    \I__8277\ : Span4Mux_s3_h
    port map (
            O => \N__33341\,
            I => \N__33335\
        );

    \I__8276\ : InMux
    port map (
            O => \N__33338\,
            I => \N__33332\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__33335\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__33332\,
            I => \M_this_external_address_qZ0Z_13\
        );

    \I__8273\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33324\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__33324\,
            I => \N__33321\
        );

    \I__8271\ : Odrv12
    port map (
            O => \N__33321\,
            I => \this_reset_cond.M_stage_qZ0Z_5\
        );

    \I__8270\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33315\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__33315\,
            I => \this_reset_cond.M_stage_qZ0Z_6\
        );

    \I__8268\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33309\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__33309\,
            I => \this_reset_cond.M_stage_qZ0Z_7\
        );

    \I__8266\ : CascadeMux
    port map (
            O => \N__33306\,
            I => \N__33302\
        );

    \I__8265\ : InMux
    port map (
            O => \N__33305\,
            I => \N__33299\
        );

    \I__8264\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33296\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__33299\,
            I => \N__33291\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__33296\,
            I => \N__33291\
        );

    \I__8261\ : Span4Mux_h
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__8260\ : Span4Mux_h
    port map (
            O => \N__33288\,
            I => \N__33285\
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__33285\,
            I => \un1_M_this_state_q_9_0_i\
        );

    \I__8258\ : IoInMux
    port map (
            O => \N__33282\,
            I => \N__33279\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__33279\,
            I => \N__33276\
        );

    \I__8256\ : Span4Mux_s3_v
    port map (
            O => \N__33276\,
            I => \N__33273\
        );

    \I__8255\ : Sp12to4
    port map (
            O => \N__33273\,
            I => \N__33270\
        );

    \I__8254\ : Span12Mux_h
    port map (
            O => \N__33270\,
            I => \N__33266\
        );

    \I__8253\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33263\
        );

    \I__8252\ : Odrv12
    port map (
            O => \N__33266\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__33263\,
            I => \M_this_external_address_qZ0Z_0\
        );

    \I__8250\ : IoInMux
    port map (
            O => \N__33258\,
            I => \N__33255\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33252\
        );

    \I__8248\ : Span4Mux_s3_v
    port map (
            O => \N__33252\,
            I => \N__33249\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__33249\,
            I => \N__33246\
        );

    \I__8246\ : Span4Mux_v
    port map (
            O => \N__33246\,
            I => \N__33242\
        );

    \I__8245\ : InMux
    port map (
            O => \N__33245\,
            I => \N__33239\
        );

    \I__8244\ : Odrv4
    port map (
            O => \N__33242\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__33239\,
            I => \M_this_external_address_qZ0Z_1\
        );

    \I__8242\ : InMux
    port map (
            O => \N__33234\,
            I => \un1_M_this_external_address_q_cry_0\
        );

    \I__8241\ : IoInMux
    port map (
            O => \N__33231\,
            I => \N__33228\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__33228\,
            I => \N__33225\
        );

    \I__8239\ : Span12Mux_s11_v
    port map (
            O => \N__33225\,
            I => \N__33221\
        );

    \I__8238\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33218\
        );

    \I__8237\ : Odrv12
    port map (
            O => \N__33221\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__33218\,
            I => \M_this_external_address_qZ0Z_2\
        );

    \I__8235\ : InMux
    port map (
            O => \N__33213\,
            I => \un1_M_this_external_address_q_cry_1\
        );

    \I__8234\ : IoInMux
    port map (
            O => \N__33210\,
            I => \N__33207\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__33207\,
            I => \N__33204\
        );

    \I__8232\ : Span4Mux_s3_h
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__8231\ : Span4Mux_v
    port map (
            O => \N__33201\,
            I => \N__33197\
        );

    \I__8230\ : InMux
    port map (
            O => \N__33200\,
            I => \N__33194\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__33197\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__33194\,
            I => \M_this_external_address_qZ0Z_3\
        );

    \I__8227\ : InMux
    port map (
            O => \N__33189\,
            I => \un1_M_this_external_address_q_cry_2\
        );

    \I__8226\ : IoInMux
    port map (
            O => \N__33186\,
            I => \N__33183\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33180\
        );

    \I__8224\ : Span4Mux_s3_h
    port map (
            O => \N__33180\,
            I => \N__33176\
        );

    \I__8223\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33173\
        );

    \I__8222\ : Odrv4
    port map (
            O => \N__33176\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__33173\,
            I => \M_this_external_address_qZ0Z_4\
        );

    \I__8220\ : InMux
    port map (
            O => \N__33168\,
            I => \un1_M_this_external_address_q_cry_3\
        );

    \I__8219\ : IoInMux
    port map (
            O => \N__33165\,
            I => \N__33162\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__33162\,
            I => \N__33158\
        );

    \I__8217\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33155\
        );

    \I__8216\ : Odrv12
    port map (
            O => \N__33158\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__33155\,
            I => \M_this_external_address_qZ0Z_5\
        );

    \I__8214\ : InMux
    port map (
            O => \N__33150\,
            I => \un1_M_this_external_address_q_cry_4\
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__33147\,
            I => \N__33144\
        );

    \I__8212\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33141\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__33141\,
            I => \N__33138\
        );

    \I__8210\ : Span4Mux_h
    port map (
            O => \N__33138\,
            I => \N__33135\
        );

    \I__8209\ : Odrv4
    port map (
            O => \N__33135\,
            I => \M_this_data_tmp_qZ0Z_18\
        );

    \I__8208\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33129\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__33129\,
            I => \N__33126\
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__33126\,
            I => \M_this_oam_ram_write_data_18\
        );

    \I__8205\ : CascadeMux
    port map (
            O => \N__33123\,
            I => \N__33120\
        );

    \I__8204\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33117\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33114\
        );

    \I__8202\ : Span4Mux_v
    port map (
            O => \N__33114\,
            I => \N__33111\
        );

    \I__8201\ : Span4Mux_v
    port map (
            O => \N__33111\,
            I => \N__33108\
        );

    \I__8200\ : Span4Mux_h
    port map (
            O => \N__33108\,
            I => \N__33105\
        );

    \I__8199\ : Odrv4
    port map (
            O => \N__33105\,
            I => \this_ppu.un1_M_vaddress_q_3_5\
        );

    \I__8198\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33099\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33096\
        );

    \I__8196\ : Odrv4
    port map (
            O => \N__33096\,
            I => \N_38_0\
        );

    \I__8195\ : InMux
    port map (
            O => \N__33093\,
            I => \N__33090\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__33090\,
            I => \M_this_oam_ram_write_data_31\
        );

    \I__8193\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N_736_0\
        );

    \I__8191\ : InMux
    port map (
            O => \N__33081\,
            I => \N__33078\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__33078\,
            I => \N_737_0\
        );

    \I__8189\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33072\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__33072\,
            I => \N__33068\
        );

    \I__8187\ : InMux
    port map (
            O => \N__33071\,
            I => \N__33063\
        );

    \I__8186\ : Span4Mux_v
    port map (
            O => \N__33068\,
            I => \N__33060\
        );

    \I__8185\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33057\
        );

    \I__8184\ : InMux
    port map (
            O => \N__33066\,
            I => \N__33054\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__33063\,
            I => \N__33047\
        );

    \I__8182\ : Span4Mux_h
    port map (
            O => \N__33060\,
            I => \N__33047\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__33057\,
            I => \N__33047\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__33054\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__8179\ : Odrv4
    port map (
            O => \N__33047\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__8178\ : InMux
    port map (
            O => \N__33042\,
            I => \N__33038\
        );

    \I__8177\ : InMux
    port map (
            O => \N__33041\,
            I => \N__33035\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__33031\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__33035\,
            I => \N__33026\
        );

    \I__8174\ : InMux
    port map (
            O => \N__33034\,
            I => \N__33023\
        );

    \I__8173\ : Span4Mux_v
    port map (
            O => \N__33031\,
            I => \N__33020\
        );

    \I__8172\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33017\
        );

    \I__8171\ : InMux
    port map (
            O => \N__33029\,
            I => \N__33014\
        );

    \I__8170\ : Span12Mux_h
    port map (
            O => \N__33026\,
            I => \N__33011\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__33023\,
            I => \N__33004\
        );

    \I__8168\ : Span4Mux_h
    port map (
            O => \N__33020\,
            I => \N__33004\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__33017\,
            I => \N__33004\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__33014\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__8165\ : Odrv12
    port map (
            O => \N__33011\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__8164\ : Odrv4
    port map (
            O => \N__33004\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__8163\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32992\
        );

    \I__8162\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32989\
        );

    \I__8161\ : CascadeMux
    port map (
            O => \N__32995\,
            I => \N__32986\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__32992\,
            I => \N__32983\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__32989\,
            I => \N__32980\
        );

    \I__8158\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32977\
        );

    \I__8157\ : Span12Mux_v
    port map (
            O => \N__32983\,
            I => \N__32974\
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__32980\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__32977\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__8154\ : Odrv12
    port map (
            O => \N__32974\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__8153\ : InMux
    port map (
            O => \N__32967\,
            I => \N__32962\
        );

    \I__8152\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32959\
        );

    \I__8151\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32956\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__32962\,
            I => \N__32953\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__32959\,
            I => \N__32950\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32944\
        );

    \I__8147\ : Span4Mux_v
    port map (
            O => \N__32953\,
            I => \N__32944\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__32950\,
            I => \N__32939\
        );

    \I__8145\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32936\
        );

    \I__8144\ : Span4Mux_v
    port map (
            O => \N__32944\,
            I => \N__32933\
        );

    \I__8143\ : InMux
    port map (
            O => \N__32943\,
            I => \N__32930\
        );

    \I__8142\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32927\
        );

    \I__8141\ : Span4Mux_h
    port map (
            O => \N__32939\,
            I => \N__32924\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__32936\,
            I => \N__32917\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__32933\,
            I => \N__32917\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__32930\,
            I => \N__32917\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__32927\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__32924\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__8135\ : Odrv4
    port map (
            O => \N__32917\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__8134\ : CascadeMux
    port map (
            O => \N__32910\,
            I => \N__32907\
        );

    \I__8133\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32904\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__8131\ : Span12Mux_h
    port map (
            O => \N__32901\,
            I => \N__32898\
        );

    \I__8130\ : Odrv12
    port map (
            O => \N__32898\,
            I => \this_ppu.un1_M_vaddress_q_3_6\
        );

    \I__8129\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32887\
        );

    \I__8128\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32887\
        );

    \I__8127\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32882\
        );

    \I__8126\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32882\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__32887\,
            I => \N__32871\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__32882\,
            I => \N__32871\
        );

    \I__8123\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32866\
        );

    \I__8122\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32866\
        );

    \I__8121\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32837\
        );

    \I__8120\ : InMux
    port map (
            O => \N__32878\,
            I => \N__32837\
        );

    \I__8119\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32832\
        );

    \I__8118\ : InMux
    port map (
            O => \N__32876\,
            I => \N__32832\
        );

    \I__8117\ : Span4Mux_v
    port map (
            O => \N__32871\,
            I => \N__32827\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__32866\,
            I => \N__32827\
        );

    \I__8115\ : InMux
    port map (
            O => \N__32865\,
            I => \N__32820\
        );

    \I__8114\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32820\
        );

    \I__8113\ : InMux
    port map (
            O => \N__32863\,
            I => \N__32820\
        );

    \I__8112\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32817\
        );

    \I__8111\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32808\
        );

    \I__8110\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32808\
        );

    \I__8109\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32808\
        );

    \I__8108\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32808\
        );

    \I__8107\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32803\
        );

    \I__8106\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32803\
        );

    \I__8105\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32798\
        );

    \I__8104\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32798\
        );

    \I__8103\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32789\
        );

    \I__8102\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32789\
        );

    \I__8101\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32789\
        );

    \I__8100\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32789\
        );

    \I__8099\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32780\
        );

    \I__8098\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32780\
        );

    \I__8097\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32780\
        );

    \I__8096\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32780\
        );

    \I__8095\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32775\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__32844\,
            I => \N__32770\
        );

    \I__8093\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32766\
        );

    \I__8092\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32763\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__32837\,
            I => \N__32754\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__32832\,
            I => \N__32754\
        );

    \I__8089\ : Span4Mux_h
    port map (
            O => \N__32827\,
            I => \N__32754\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__32820\,
            I => \N__32754\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__32817\,
            I => \N__32747\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__32808\,
            I => \N__32747\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__32803\,
            I => \N__32747\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__32798\,
            I => \N__32744\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__32789\,
            I => \N__32739\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__32780\,
            I => \N__32739\
        );

    \I__8081\ : InMux
    port map (
            O => \N__32779\,
            I => \N__32736\
        );

    \I__8080\ : InMux
    port map (
            O => \N__32778\,
            I => \N__32733\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__32775\,
            I => \N__32730\
        );

    \I__8078\ : InMux
    port map (
            O => \N__32774\,
            I => \N__32721\
        );

    \I__8077\ : InMux
    port map (
            O => \N__32773\,
            I => \N__32721\
        );

    \I__8076\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32721\
        );

    \I__8075\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32721\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__32766\,
            I => \N__32710\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__32763\,
            I => \N__32710\
        );

    \I__8072\ : Span4Mux_v
    port map (
            O => \N__32754\,
            I => \N__32710\
        );

    \I__8071\ : Span4Mux_v
    port map (
            O => \N__32747\,
            I => \N__32710\
        );

    \I__8070\ : Span4Mux_v
    port map (
            O => \N__32744\,
            I => \N__32710\
        );

    \I__8069\ : Span4Mux_h
    port map (
            O => \N__32739\,
            I => \N__32707\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__32736\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__32733\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8066\ : Odrv12
    port map (
            O => \N__32730\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__32721\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__32710\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8063\ : Odrv4
    port map (
            O => \N__32707\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__32694\,
            I => \N__32673\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__32693\,
            I => \N__32670\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__32692\,
            I => \N__32661\
        );

    \I__8059\ : CascadeMux
    port map (
            O => \N__32691\,
            I => \N__32658\
        );

    \I__8058\ : CascadeMux
    port map (
            O => \N__32690\,
            I => \N__32649\
        );

    \I__8057\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32646\
        );

    \I__8056\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32641\
        );

    \I__8055\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32641\
        );

    \I__8054\ : InMux
    port map (
            O => \N__32686\,
            I => \N__32638\
        );

    \I__8053\ : InMux
    port map (
            O => \N__32685\,
            I => \N__32633\
        );

    \I__8052\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32633\
        );

    \I__8051\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32628\
        );

    \I__8050\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32628\
        );

    \I__8049\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32623\
        );

    \I__8048\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32623\
        );

    \I__8047\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32618\
        );

    \I__8046\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32618\
        );

    \I__8045\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32613\
        );

    \I__8044\ : InMux
    port map (
            O => \N__32676\,
            I => \N__32613\
        );

    \I__8043\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32606\
        );

    \I__8042\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32606\
        );

    \I__8041\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32606\
        );

    \I__8040\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32601\
        );

    \I__8039\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32601\
        );

    \I__8038\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32598\
        );

    \I__8037\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32591\
        );

    \I__8036\ : InMux
    port map (
            O => \N__32664\,
            I => \N__32591\
        );

    \I__8035\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32591\
        );

    \I__8034\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32588\
        );

    \I__8033\ : CascadeMux
    port map (
            O => \N__32657\,
            I => \N__32583\
        );

    \I__8032\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32575\
        );

    \I__8031\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32575\
        );

    \I__8030\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32575\
        );

    \I__8029\ : InMux
    port map (
            O => \N__32653\,
            I => \N__32566\
        );

    \I__8028\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32566\
        );

    \I__8027\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32563\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__32646\,
            I => \N__32560\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32557\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32538\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__32633\,
            I => \N__32538\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__32628\,
            I => \N__32538\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__32623\,
            I => \N__32538\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__32618\,
            I => \N__32538\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32538\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__32606\,
            I => \N__32538\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__32601\,
            I => \N__32538\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__32598\,
            I => \N__32538\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__32591\,
            I => \N__32533\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__32588\,
            I => \N__32533\
        );

    \I__8013\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32524\
        );

    \I__8012\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32524\
        );

    \I__8011\ : InMux
    port map (
            O => \N__32583\,
            I => \N__32524\
        );

    \I__8010\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32524\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__32575\,
            I => \N__32521\
        );

    \I__8008\ : InMux
    port map (
            O => \N__32574\,
            I => \N__32516\
        );

    \I__8007\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32516\
        );

    \I__8006\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32513\
        );

    \I__8005\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32510\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32507\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__32563\,
            I => \N__32502\
        );

    \I__8002\ : Span4Mux_v
    port map (
            O => \N__32560\,
            I => \N__32502\
        );

    \I__8001\ : Span4Mux_v
    port map (
            O => \N__32557\,
            I => \N__32495\
        );

    \I__8000\ : Span4Mux_v
    port map (
            O => \N__32538\,
            I => \N__32495\
        );

    \I__7999\ : Span4Mux_v
    port map (
            O => \N__32533\,
            I => \N__32495\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__32524\,
            I => \N__32490\
        );

    \I__7997\ : Span4Mux_h
    port map (
            O => \N__32521\,
            I => \N__32490\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__32516\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__32513\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__32510\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7993\ : Odrv12
    port map (
            O => \N__32507\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7992\ : Odrv4
    port map (
            O => \N__32502\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7991\ : Odrv4
    port map (
            O => \N__32495\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7990\ : Odrv4
    port map (
            O => \N__32490\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__32475\,
            I => \N__32472\
        );

    \I__7988\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32469\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__32469\,
            I => \N__32466\
        );

    \I__7986\ : Odrv4
    port map (
            O => \N__32466\,
            I => \M_this_data_tmp_qZ0Z_21\
        );

    \I__7985\ : InMux
    port map (
            O => \N__32463\,
            I => \N__32444\
        );

    \I__7984\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32444\
        );

    \I__7983\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32444\
        );

    \I__7982\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32444\
        );

    \I__7981\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32421\
        );

    \I__7980\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32421\
        );

    \I__7979\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32414\
        );

    \I__7978\ : InMux
    port map (
            O => \N__32456\,
            I => \N__32414\
        );

    \I__7977\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32414\
        );

    \I__7976\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32409\
        );

    \I__7975\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32409\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__32444\,
            I => \N__32406\
        );

    \I__7973\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32403\
        );

    \I__7972\ : InMux
    port map (
            O => \N__32442\,
            I => \N__32394\
        );

    \I__7971\ : InMux
    port map (
            O => \N__32441\,
            I => \N__32394\
        );

    \I__7970\ : InMux
    port map (
            O => \N__32440\,
            I => \N__32394\
        );

    \I__7969\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32394\
        );

    \I__7968\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32385\
        );

    \I__7967\ : InMux
    port map (
            O => \N__32437\,
            I => \N__32385\
        );

    \I__7966\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32385\
        );

    \I__7965\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32385\
        );

    \I__7964\ : InMux
    port map (
            O => \N__32434\,
            I => \N__32378\
        );

    \I__7963\ : InMux
    port map (
            O => \N__32433\,
            I => \N__32378\
        );

    \I__7962\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32368\
        );

    \I__7961\ : InMux
    port map (
            O => \N__32431\,
            I => \N__32368\
        );

    \I__7960\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32359\
        );

    \I__7959\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32359\
        );

    \I__7958\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32359\
        );

    \I__7957\ : InMux
    port map (
            O => \N__32427\,
            I => \N__32359\
        );

    \I__7956\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32356\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__32421\,
            I => \N__32349\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__32414\,
            I => \N__32349\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32349\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__32406\,
            I => \N__32340\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__32403\,
            I => \N__32340\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__32394\,
            I => \N__32340\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__32385\,
            I => \N__32340\
        );

    \I__7948\ : CascadeMux
    port map (
            O => \N__32384\,
            I => \N__32337\
        );

    \I__7947\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32332\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__32378\,
            I => \N__32329\
        );

    \I__7945\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32326\
        );

    \I__7944\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32323\
        );

    \I__7943\ : InMux
    port map (
            O => \N__32375\,
            I => \N__32320\
        );

    \I__7942\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32315\
        );

    \I__7941\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32315\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32310\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__32359\,
            I => \N__32310\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__32356\,
            I => \N__32303\
        );

    \I__7937\ : Span4Mux_v
    port map (
            O => \N__32349\,
            I => \N__32303\
        );

    \I__7936\ : Span4Mux_v
    port map (
            O => \N__32340\,
            I => \N__32303\
        );

    \I__7935\ : InMux
    port map (
            O => \N__32337\,
            I => \N__32296\
        );

    \I__7934\ : InMux
    port map (
            O => \N__32336\,
            I => \N__32296\
        );

    \I__7933\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32296\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__32332\,
            I => \N__32287\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__32329\,
            I => \N__32287\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__32326\,
            I => \N__32287\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__32323\,
            I => \N__32287\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__32320\,
            I => \N__32280\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__32315\,
            I => \N__32280\
        );

    \I__7926\ : Span4Mux_v
    port map (
            O => \N__32310\,
            I => \N__32280\
        );

    \I__7925\ : Span4Mux_v
    port map (
            O => \N__32303\,
            I => \N__32277\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32270\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__32287\,
            I => \N__32270\
        );

    \I__7922\ : Span4Mux_h
    port map (
            O => \N__32280\,
            I => \N__32270\
        );

    \I__7921\ : Odrv4
    port map (
            O => \N__32277\,
            I => \N_122_0\
        );

    \I__7920\ : Odrv4
    port map (
            O => \N__32270\,
            I => \N_122_0\
        );

    \I__7919\ : InMux
    port map (
            O => \N__32265\,
            I => \N__32262\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__32262\,
            I => \M_this_oam_ram_write_data_21\
        );

    \I__7917\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32256\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__32256\,
            I => \N__32252\
        );

    \I__7915\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32249\
        );

    \I__7914\ : Span12Mux_s11_v
    port map (
            O => \N__32252\,
            I => \N__32246\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__32249\,
            I => \N__32243\
        );

    \I__7912\ : Span12Mux_v
    port map (
            O => \N__32246\,
            I => \N__32240\
        );

    \I__7911\ : Span4Mux_h
    port map (
            O => \N__32243\,
            I => \N__32237\
        );

    \I__7910\ : Odrv12
    port map (
            O => \N__32240\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__32237\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__7908\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32229\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__32229\,
            I => \N__32226\
        );

    \I__7906\ : Span4Mux_h
    port map (
            O => \N__32226\,
            I => \N__32222\
        );

    \I__7905\ : InMux
    port map (
            O => \N__32225\,
            I => \N__32219\
        );

    \I__7904\ : Span4Mux_h
    port map (
            O => \N__32222\,
            I => \N__32214\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__32219\,
            I => \N__32214\
        );

    \I__7902\ : Odrv4
    port map (
            O => \N__32214\,
            I => \M_this_oam_ram_read_data_5\
        );

    \I__7901\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32208\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32205\
        );

    \I__7899\ : Span4Mux_v
    port map (
            O => \N__32205\,
            I => \N__32202\
        );

    \I__7898\ : Sp12to4
    port map (
            O => \N__32202\,
            I => \N__32198\
        );

    \I__7897\ : CascadeMux
    port map (
            O => \N__32201\,
            I => \N__32195\
        );

    \I__7896\ : Span12Mux_h
    port map (
            O => \N__32198\,
            I => \N__32192\
        );

    \I__7895\ : InMux
    port map (
            O => \N__32195\,
            I => \N__32189\
        );

    \I__7894\ : Span12Mux_v
    port map (
            O => \N__32192\,
            I => \N__32186\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__32189\,
            I => \N__32183\
        );

    \I__7892\ : Odrv12
    port map (
            O => \N__32186\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__7891\ : Odrv4
    port map (
            O => \N__32183\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__7890\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32175\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__32175\,
            I => \N__32171\
        );

    \I__7888\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32168\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__32171\,
            I => \N__32165\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32162\
        );

    \I__7885\ : Odrv4
    port map (
            O => \N__32165\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__32162\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__7883\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32154\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__32154\,
            I => \N__32151\
        );

    \I__7881\ : Span4Mux_h
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__7880\ : Span4Mux_h
    port map (
            O => \N__32148\,
            I => \N__32145\
        );

    \I__7879\ : Odrv4
    port map (
            O => \N__32145\,
            I => \this_ppu.un9lto7Z0Z_4\
        );

    \I__7878\ : CascadeMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__7877\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32136\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__32136\,
            I => \N__32133\
        );

    \I__7875\ : Odrv4
    port map (
            O => \N__32133\,
            I => \M_this_data_tmp_qZ0Z_9\
        );

    \I__7874\ : InMux
    port map (
            O => \N__32130\,
            I => \N__32127\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__32127\,
            I => \N_741_0\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__32124\,
            I => \N__32121\
        );

    \I__7871\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32118\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__32118\,
            I => \N__32115\
        );

    \I__7869\ : Span4Mux_v
    port map (
            O => \N__32115\,
            I => \N__32112\
        );

    \I__7868\ : Span4Mux_h
    port map (
            O => \N__32112\,
            I => \N__32108\
        );

    \I__7867\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32105\
        );

    \I__7866\ : Span4Mux_h
    port map (
            O => \N__32108\,
            I => \N__32100\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__32105\,
            I => \N__32100\
        );

    \I__7864\ : Odrv4
    port map (
            O => \N__32100\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__7863\ : CascadeMux
    port map (
            O => \N__32097\,
            I => \this_ppu.un1_oam_data_c2_cascade_\
        );

    \I__7862\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32091\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__32091\,
            I => \N__32088\
        );

    \I__7860\ : Span4Mux_v
    port map (
            O => \N__32088\,
            I => \N__32085\
        );

    \I__7859\ : Span4Mux_h
    port map (
            O => \N__32085\,
            I => \N__32082\
        );

    \I__7858\ : Odrv4
    port map (
            O => \N__32082\,
            I => \this_ppu.un1_M_vaddress_q_3_7\
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__32079\,
            I => \N__32076\
        );

    \I__7856\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32073\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__32073\,
            I => \N__32070\
        );

    \I__7854\ : Odrv4
    port map (
            O => \N__32070\,
            I => \M_this_data_tmp_qZ0Z_13\
        );

    \I__7853\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32064\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__32064\,
            I => \M_this_oam_ram_write_data_13\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__32061\,
            I => \N__32058\
        );

    \I__7850\ : InMux
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__32055\,
            I => \N__32052\
        );

    \I__7848\ : Span4Mux_v
    port map (
            O => \N__32052\,
            I => \N__32049\
        );

    \I__7847\ : Span4Mux_h
    port map (
            O => \N__32049\,
            I => \N__32046\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__32046\,
            I => \M_this_data_tmp_qZ0Z_15\
        );

    \I__7845\ : InMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__32040\,
            I => \M_this_oam_ram_write_data_15\
        );

    \I__7843\ : CEMux
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__32034\,
            I => \N__32030\
        );

    \I__7841\ : CEMux
    port map (
            O => \N__32033\,
            I => \N__32027\
        );

    \I__7840\ : Span4Mux_v
    port map (
            O => \N__32030\,
            I => \N__32024\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__32021\
        );

    \I__7838\ : Span4Mux_h
    port map (
            O => \N__32024\,
            I => \N__32018\
        );

    \I__7837\ : Span4Mux_h
    port map (
            O => \N__32021\,
            I => \N__32015\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__32018\,
            I => \N_123_0\
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__32015\,
            I => \N_123_0\
        );

    \I__7834\ : InMux
    port map (
            O => \N__32010\,
            I => \N__32006\
        );

    \I__7833\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32003\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__32006\,
            I => \N__32000\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__32003\,
            I => \N__31997\
        );

    \I__7830\ : Span12Mux_h
    port map (
            O => \N__32000\,
            I => \N__31994\
        );

    \I__7829\ : Span4Mux_h
    port map (
            O => \N__31997\,
            I => \N__31991\
        );

    \I__7828\ : Odrv12
    port map (
            O => \N__31994\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__7827\ : Odrv4
    port map (
            O => \N__31991\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__31986\,
            I => \N__31983\
        );

    \I__7825\ : InMux
    port map (
            O => \N__31983\,
            I => \N__31980\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__31980\,
            I => \N__31977\
        );

    \I__7823\ : Span4Mux_h
    port map (
            O => \N__31977\,
            I => \N__31974\
        );

    \I__7822\ : Span4Mux_v
    port map (
            O => \N__31974\,
            I => \N__31970\
        );

    \I__7821\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31967\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__31970\,
            I => \N__31964\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__31967\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__31964\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__7817\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31955\
        );

    \I__7816\ : CascadeMux
    port map (
            O => \N__31958\,
            I => \N__31952\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__31955\,
            I => \N__31949\
        );

    \I__7814\ : InMux
    port map (
            O => \N__31952\,
            I => \N__31946\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__31949\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__31946\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__7811\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31938\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__31938\,
            I => \N__31935\
        );

    \I__7809\ : Span4Mux_v
    port map (
            O => \N__31935\,
            I => \N__31932\
        );

    \I__7808\ : Span4Mux_v
    port map (
            O => \N__31932\,
            I => \N__31929\
        );

    \I__7807\ : Span4Mux_v
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__7806\ : Span4Mux_h
    port map (
            O => \N__31926\,
            I => \N__31922\
        );

    \I__7805\ : InMux
    port map (
            O => \N__31925\,
            I => \N__31919\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__31922\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__31919\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__7802\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31911\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__31911\,
            I => \N__31908\
        );

    \I__7800\ : Span4Mux_h
    port map (
            O => \N__31908\,
            I => \N__31905\
        );

    \I__7799\ : Span4Mux_h
    port map (
            O => \N__31905\,
            I => \N__31902\
        );

    \I__7798\ : Odrv4
    port map (
            O => \N__31902\,
            I => \this_ppu.un9lto7Z0Z_5\
        );

    \I__7797\ : CascadeMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__7796\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31892\
        );

    \I__7795\ : CascadeMux
    port map (
            O => \N__31895\,
            I => \N__31889\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__31892\,
            I => \N__31886\
        );

    \I__7793\ : InMux
    port map (
            O => \N__31889\,
            I => \N__31883\
        );

    \I__7792\ : Span4Mux_h
    port map (
            O => \N__31886\,
            I => \N__31880\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__31883\,
            I => \N__31877\
        );

    \I__7790\ : Span4Mux_v
    port map (
            O => \N__31880\,
            I => \N__31874\
        );

    \I__7789\ : Span4Mux_h
    port map (
            O => \N__31877\,
            I => \N__31870\
        );

    \I__7788\ : Span4Mux_v
    port map (
            O => \N__31874\,
            I => \N__31867\
        );

    \I__7787\ : InMux
    port map (
            O => \N__31873\,
            I => \N__31864\
        );

    \I__7786\ : Span4Mux_v
    port map (
            O => \N__31870\,
            I => \N__31861\
        );

    \I__7785\ : Span4Mux_h
    port map (
            O => \N__31867\,
            I => \N__31858\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__31864\,
            I => \N__31853\
        );

    \I__7783\ : Span4Mux_h
    port map (
            O => \N__31861\,
            I => \N__31853\
        );

    \I__7782\ : Odrv4
    port map (
            O => \N__31858\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__7781\ : Odrv4
    port map (
            O => \N__31853\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__31848\,
            I => \N__31845\
        );

    \I__7779\ : InMux
    port map (
            O => \N__31845\,
            I => \N__31842\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__31842\,
            I => \N__31839\
        );

    \I__7777\ : Odrv12
    port map (
            O => \N__31839\,
            I => \M_this_oam_ram_read_data_i_17\
        );

    \I__7776\ : CascadeMux
    port map (
            O => \N__31836\,
            I => \N__31832\
        );

    \I__7775\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31829\
        );

    \I__7774\ : InMux
    port map (
            O => \N__31832\,
            I => \N__31826\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31820\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__31826\,
            I => \N__31820\
        );

    \I__7771\ : InMux
    port map (
            O => \N__31825\,
            I => \N__31817\
        );

    \I__7770\ : Span4Mux_h
    port map (
            O => \N__31820\,
            I => \N__31812\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__31817\,
            I => \N__31812\
        );

    \I__7768\ : Span4Mux_h
    port map (
            O => \N__31812\,
            I => \N__31809\
        );

    \I__7767\ : Odrv4
    port map (
            O => \N__31809\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__7766\ : InMux
    port map (
            O => \N__31806\,
            I => \this_ppu.un2_hscroll_cry_1\
        );

    \I__7765\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31800\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__31800\,
            I => \N__31797\
        );

    \I__7763\ : Odrv12
    port map (
            O => \N__31797\,
            I => \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\
        );

    \I__7762\ : CascadeMux
    port map (
            O => \N__31794\,
            I => \N__31791\
        );

    \I__7761\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31786\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__31790\,
            I => \N__31783\
        );

    \I__7759\ : InMux
    port map (
            O => \N__31789\,
            I => \N__31780\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__31786\,
            I => \N__31777\
        );

    \I__7757\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31774\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31771\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__31777\,
            I => \N__31766\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__31774\,
            I => \N__31766\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__31771\,
            I => \N__31761\
        );

    \I__7752\ : Span4Mux_h
    port map (
            O => \N__31766\,
            I => \N__31761\
        );

    \I__7751\ : Span4Mux_v
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__31758\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__31755\,
            I => \N__31752\
        );

    \I__7748\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31749\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__31749\,
            I => \M_this_oam_ram_read_data_i_9\
        );

    \I__7746\ : CascadeMux
    port map (
            O => \N__31746\,
            I => \N__31743\
        );

    \I__7745\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31737\
        );

    \I__7743\ : Odrv12
    port map (
            O => \N__31737\,
            I => \M_this_data_tmp_qZ0Z_1\
        );

    \I__7742\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__7740\ : Span4Mux_v
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__31725\,
            I => \N_747_0\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__31722\,
            I => \N__31719\
        );

    \I__7737\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__31716\,
            I => \M_this_data_tmp_qZ0Z_10\
        );

    \I__7735\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31710\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__7733\ : Odrv4
    port map (
            O => \N__31707\,
            I => \M_this_oam_ram_write_data_10\
        );

    \I__7732\ : InMux
    port map (
            O => \N__31704\,
            I => \N__31701\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__31701\,
            I => \N__31698\
        );

    \I__7730\ : Span4Mux_h
    port map (
            O => \N__31698\,
            I => \N__31695\
        );

    \I__7729\ : Span4Mux_h
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__7728\ : Span4Mux_h
    port map (
            O => \N__31692\,
            I => \N__31689\
        );

    \I__7727\ : Span4Mux_h
    port map (
            O => \N__31689\,
            I => \N__31686\
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__31686\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__31683\,
            I => \N__31679\
        );

    \I__7724\ : CascadeMux
    port map (
            O => \N__31682\,
            I => \N__31674\
        );

    \I__7723\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31668\
        );

    \I__7722\ : CascadeMux
    port map (
            O => \N__31678\,
            I => \N__31664\
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__31677\,
            I => \N__31660\
        );

    \I__7720\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31657\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__31673\,
            I => \N__31654\
        );

    \I__7718\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31649\
        );

    \I__7717\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31646\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31643\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__31667\,
            I => \N__31639\
        );

    \I__7714\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31636\
        );

    \I__7713\ : CascadeMux
    port map (
            O => \N__31663\,
            I => \N__31633\
        );

    \I__7712\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31630\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__31657\,
            I => \N__31627\
        );

    \I__7710\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31624\
        );

    \I__7709\ : CascadeMux
    port map (
            O => \N__31653\,
            I => \N__31621\
        );

    \I__7708\ : CascadeMux
    port map (
            O => \N__31652\,
            I => \N__31618\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__31649\,
            I => \N__31615\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__31646\,
            I => \N__31612\
        );

    \I__7705\ : Span4Mux_h
    port map (
            O => \N__31643\,
            I => \N__31609\
        );

    \I__7704\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31604\
        );

    \I__7703\ : InMux
    port map (
            O => \N__31639\,
            I => \N__31604\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__31636\,
            I => \N__31601\
        );

    \I__7701\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31598\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__31630\,
            I => \N__31595\
        );

    \I__7699\ : Span4Mux_h
    port map (
            O => \N__31627\,
            I => \N__31592\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__31624\,
            I => \N__31589\
        );

    \I__7697\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31586\
        );

    \I__7696\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31583\
        );

    \I__7695\ : Span4Mux_v
    port map (
            O => \N__31615\,
            I => \N__31579\
        );

    \I__7694\ : Span4Mux_v
    port map (
            O => \N__31612\,
            I => \N__31571\
        );

    \I__7693\ : Span4Mux_h
    port map (
            O => \N__31609\,
            I => \N__31571\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__31604\,
            I => \N__31571\
        );

    \I__7691\ : Span4Mux_h
    port map (
            O => \N__31601\,
            I => \N__31566\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__31598\,
            I => \N__31566\
        );

    \I__7689\ : Span4Mux_h
    port map (
            O => \N__31595\,
            I => \N__31563\
        );

    \I__7688\ : Span4Mux_v
    port map (
            O => \N__31592\,
            I => \N__31556\
        );

    \I__7687\ : Span4Mux_h
    port map (
            O => \N__31589\,
            I => \N__31556\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31556\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__31583\,
            I => \N__31553\
        );

    \I__7684\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31549\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__31579\,
            I => \N__31546\
        );

    \I__7682\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31543\
        );

    \I__7681\ : Span4Mux_v
    port map (
            O => \N__31571\,
            I => \N__31536\
        );

    \I__7680\ : Span4Mux_h
    port map (
            O => \N__31566\,
            I => \N__31536\
        );

    \I__7679\ : Span4Mux_h
    port map (
            O => \N__31563\,
            I => \N__31536\
        );

    \I__7678\ : Span4Mux_v
    port map (
            O => \N__31556\,
            I => \N__31531\
        );

    \I__7677\ : Span4Mux_h
    port map (
            O => \N__31553\,
            I => \N__31531\
        );

    \I__7676\ : InMux
    port map (
            O => \N__31552\,
            I => \N__31528\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__31549\,
            I => \N__31525\
        );

    \I__7674\ : Span4Mux_v
    port map (
            O => \N__31546\,
            I => \N__31520\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__31543\,
            I => \N__31520\
        );

    \I__7672\ : Span4Mux_v
    port map (
            O => \N__31536\,
            I => \N__31517\
        );

    \I__7671\ : Span4Mux_h
    port map (
            O => \N__31531\,
            I => \N__31512\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__31528\,
            I => \N__31512\
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__31525\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7668\ : Odrv4
    port map (
            O => \N__31520\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7667\ : Odrv4
    port map (
            O => \N__31517\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__31512\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__7665\ : CascadeMux
    port map (
            O => \N__31503\,
            I => \N__31496\
        );

    \I__7664\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31493\
        );

    \I__7663\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31489\
        );

    \I__7662\ : InMux
    port map (
            O => \N__31500\,
            I => \N__31486\
        );

    \I__7661\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31483\
        );

    \I__7660\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31474\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__31493\,
            I => \N__31471\
        );

    \I__7658\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31468\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__31489\,
            I => \N__31465\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__31486\,
            I => \N__31461\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31458\
        );

    \I__7654\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31454\
        );

    \I__7653\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31449\
        );

    \I__7652\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31446\
        );

    \I__7651\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31441\
        );

    \I__7650\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31441\
        );

    \I__7649\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31438\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__31474\,
            I => \N__31434\
        );

    \I__7647\ : Span4Mux_h
    port map (
            O => \N__31471\,
            I => \N__31429\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__31468\,
            I => \N__31429\
        );

    \I__7645\ : Span4Mux_v
    port map (
            O => \N__31465\,
            I => \N__31426\
        );

    \I__7644\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31423\
        );

    \I__7643\ : Span4Mux_h
    port map (
            O => \N__31461\,
            I => \N__31418\
        );

    \I__7642\ : Span4Mux_h
    port map (
            O => \N__31458\,
            I => \N__31418\
        );

    \I__7641\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31415\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__31454\,
            I => \N__31412\
        );

    \I__7639\ : InMux
    port map (
            O => \N__31453\,
            I => \N__31407\
        );

    \I__7638\ : InMux
    port map (
            O => \N__31452\,
            I => \N__31407\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__31449\,
            I => \N__31404\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__31446\,
            I => \N__31399\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__31441\,
            I => \N__31399\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__31438\,
            I => \N__31396\
        );

    \I__7633\ : InMux
    port map (
            O => \N__31437\,
            I => \N__31393\
        );

    \I__7632\ : Span4Mux_h
    port map (
            O => \N__31434\,
            I => \N__31388\
        );

    \I__7631\ : Span4Mux_h
    port map (
            O => \N__31429\,
            I => \N__31388\
        );

    \I__7630\ : Sp12to4
    port map (
            O => \N__31426\,
            I => \N__31383\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__31423\,
            I => \N__31383\
        );

    \I__7628\ : Sp12to4
    port map (
            O => \N__31418\,
            I => \N__31378\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__31415\,
            I => \N__31378\
        );

    \I__7626\ : Span4Mux_h
    port map (
            O => \N__31412\,
            I => \N__31375\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__31407\,
            I => \N__31372\
        );

    \I__7624\ : Span4Mux_v
    port map (
            O => \N__31404\,
            I => \N__31367\
        );

    \I__7623\ : Span4Mux_v
    port map (
            O => \N__31399\,
            I => \N__31367\
        );

    \I__7622\ : Span4Mux_h
    port map (
            O => \N__31396\,
            I => \N__31364\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__31393\,
            I => \N__31361\
        );

    \I__7620\ : Sp12to4
    port map (
            O => \N__31388\,
            I => \N__31356\
        );

    \I__7619\ : Span12Mux_h
    port map (
            O => \N__31383\,
            I => \N__31356\
        );

    \I__7618\ : Span12Mux_v
    port map (
            O => \N__31378\,
            I => \N__31353\
        );

    \I__7617\ : Span4Mux_h
    port map (
            O => \N__31375\,
            I => \N__31346\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__31372\,
            I => \N__31346\
        );

    \I__7615\ : Span4Mux_v
    port map (
            O => \N__31367\,
            I => \N__31346\
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__31364\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7613\ : Odrv12
    port map (
            O => \N__31361\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7612\ : Odrv12
    port map (
            O => \N__31356\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7611\ : Odrv12
    port map (
            O => \N__31353\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7610\ : Odrv4
    port map (
            O => \N__31346\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__7609\ : CascadeMux
    port map (
            O => \N__31335\,
            I => \N__31331\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__31334\,
            I => \N__31326\
        );

    \I__7607\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31322\
        );

    \I__7606\ : CascadeMux
    port map (
            O => \N__31330\,
            I => \N__31319\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__31329\,
            I => \N__31316\
        );

    \I__7604\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31311\
        );

    \I__7603\ : CascadeMux
    port map (
            O => \N__31325\,
            I => \N__31308\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__31322\,
            I => \N__31304\
        );

    \I__7601\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31301\
        );

    \I__7600\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31298\
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__31315\,
            I => \N__31295\
        );

    \I__7598\ : CascadeMux
    port map (
            O => \N__31314\,
            I => \N__31292\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__31311\,
            I => \N__31288\
        );

    \I__7596\ : InMux
    port map (
            O => \N__31308\,
            I => \N__31285\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__31307\,
            I => \N__31282\
        );

    \I__7594\ : Span4Mux_h
    port map (
            O => \N__31304\,
            I => \N__31278\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__31301\,
            I => \N__31275\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__31298\,
            I => \N__31272\
        );

    \I__7591\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31269\
        );

    \I__7590\ : InMux
    port map (
            O => \N__31292\,
            I => \N__31266\
        );

    \I__7589\ : CascadeMux
    port map (
            O => \N__31291\,
            I => \N__31263\
        );

    \I__7588\ : Span4Mux_h
    port map (
            O => \N__31288\,
            I => \N__31258\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__31285\,
            I => \N__31255\
        );

    \I__7586\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31252\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__31281\,
            I => \N__31249\
        );

    \I__7584\ : Span4Mux_v
    port map (
            O => \N__31278\,
            I => \N__31243\
        );

    \I__7583\ : Span4Mux_h
    port map (
            O => \N__31275\,
            I => \N__31243\
        );

    \I__7582\ : Span4Mux_v
    port map (
            O => \N__31272\,
            I => \N__31240\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31237\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__31266\,
            I => \N__31234\
        );

    \I__7579\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31231\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__31262\,
            I => \N__31228\
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__31261\,
            I => \N__31224\
        );

    \I__7576\ : Span4Mux_v
    port map (
            O => \N__31258\,
            I => \N__31219\
        );

    \I__7575\ : Span4Mux_h
    port map (
            O => \N__31255\,
            I => \N__31219\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31216\
        );

    \I__7573\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31213\
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__31248\,
            I => \N__31210\
        );

    \I__7571\ : Span4Mux_v
    port map (
            O => \N__31243\,
            I => \N__31203\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__31240\,
            I => \N__31203\
        );

    \I__7569\ : Span4Mux_h
    port map (
            O => \N__31237\,
            I => \N__31203\
        );

    \I__7568\ : Span4Mux_h
    port map (
            O => \N__31234\,
            I => \N__31200\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__31231\,
            I => \N__31197\
        );

    \I__7566\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31194\
        );

    \I__7565\ : CascadeMux
    port map (
            O => \N__31227\,
            I => \N__31191\
        );

    \I__7564\ : InMux
    port map (
            O => \N__31224\,
            I => \N__31187\
        );

    \I__7563\ : Span4Mux_v
    port map (
            O => \N__31219\,
            I => \N__31182\
        );

    \I__7562\ : Span4Mux_h
    port map (
            O => \N__31216\,
            I => \N__31182\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__31213\,
            I => \N__31179\
        );

    \I__7560\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31176\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__31203\,
            I => \N__31173\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__31200\,
            I => \N__31168\
        );

    \I__7557\ : Span4Mux_h
    port map (
            O => \N__31197\,
            I => \N__31168\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31165\
        );

    \I__7555\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31162\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__31190\,
            I => \N__31159\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__31187\,
            I => \N__31156\
        );

    \I__7552\ : Span4Mux_v
    port map (
            O => \N__31182\,
            I => \N__31151\
        );

    \I__7551\ : Span4Mux_h
    port map (
            O => \N__31179\,
            I => \N__31151\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__31176\,
            I => \N__31148\
        );

    \I__7549\ : Span4Mux_h
    port map (
            O => \N__31173\,
            I => \N__31145\
        );

    \I__7548\ : Span4Mux_v
    port map (
            O => \N__31168\,
            I => \N__31140\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__31165\,
            I => \N__31140\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__31162\,
            I => \N__31137\
        );

    \I__7545\ : InMux
    port map (
            O => \N__31159\,
            I => \N__31134\
        );

    \I__7544\ : Span12Mux_h
    port map (
            O => \N__31156\,
            I => \N__31130\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__31151\,
            I => \N__31125\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__31148\,
            I => \N__31125\
        );

    \I__7541\ : Span4Mux_h
    port map (
            O => \N__31145\,
            I => \N__31118\
        );

    \I__7540\ : Span4Mux_v
    port map (
            O => \N__31140\,
            I => \N__31118\
        );

    \I__7539\ : Span4Mux_h
    port map (
            O => \N__31137\,
            I => \N__31118\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31115\
        );

    \I__7537\ : CascadeMux
    port map (
            O => \N__31133\,
            I => \N__31112\
        );

    \I__7536\ : Span12Mux_v
    port map (
            O => \N__31130\,
            I => \N__31109\
        );

    \I__7535\ : Span4Mux_v
    port map (
            O => \N__31125\,
            I => \N__31106\
        );

    \I__7534\ : Span4Mux_v
    port map (
            O => \N__31118\,
            I => \N__31101\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__31115\,
            I => \N__31101\
        );

    \I__7532\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31098\
        );

    \I__7531\ : Odrv12
    port map (
            O => \N__31109\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__31106\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__7529\ : Odrv4
    port map (
            O => \N__31101\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__31098\,
            I => \M_this_ppu_sprites_addr_9\
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__7526\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31083\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__31080\,
            I => \N__31077\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__31077\,
            I => \M_this_data_tmp_qZ0Z_12\
        );

    \I__7522\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31071\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__31071\,
            I => \N_740_0\
        );

    \I__7520\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31064\
        );

    \I__7519\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31060\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__31064\,
            I => \N__31057\
        );

    \I__7517\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31054\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__31060\,
            I => \N__31051\
        );

    \I__7515\ : Span4Mux_h
    port map (
            O => \N__31057\,
            I => \N__31047\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__31042\
        );

    \I__7513\ : Span4Mux_h
    port map (
            O => \N__31051\,
            I => \N__31042\
        );

    \I__7512\ : InMux
    port map (
            O => \N__31050\,
            I => \N__31039\
        );

    \I__7511\ : Span4Mux_h
    port map (
            O => \N__31047\,
            I => \N__31036\
        );

    \I__7510\ : Span4Mux_h
    port map (
            O => \N__31042\,
            I => \N__31033\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__31039\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7508\ : Odrv4
    port map (
            O => \N__31036\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7507\ : Odrv4
    port map (
            O => \N__31033\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__7506\ : CascadeMux
    port map (
            O => \N__31026\,
            I => \N__31022\
        );

    \I__7505\ : InMux
    port map (
            O => \N__31025\,
            I => \N__31018\
        );

    \I__7504\ : InMux
    port map (
            O => \N__31022\,
            I => \N__31013\
        );

    \I__7503\ : InMux
    port map (
            O => \N__31021\,
            I => \N__31013\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__31018\,
            I => \N__31009\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__31013\,
            I => \N__31006\
        );

    \I__7500\ : InMux
    port map (
            O => \N__31012\,
            I => \N__31003\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__31009\,
            I => \N__30999\
        );

    \I__7498\ : Span4Mux_h
    port map (
            O => \N__31006\,
            I => \N__30994\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__31003\,
            I => \N__30994\
        );

    \I__7496\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30991\
        );

    \I__7495\ : Span4Mux_h
    port map (
            O => \N__30999\,
            I => \N__30988\
        );

    \I__7494\ : Span4Mux_h
    port map (
            O => \N__30994\,
            I => \N__30985\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__30991\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__30988\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__30985\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__7490\ : CascadeMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__7489\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30971\
        );

    \I__7488\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30967\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__30971\,
            I => \N__30964\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__30970\,
            I => \N__30961\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__30967\,
            I => \N__30956\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__30964\,
            I => \N__30956\
        );

    \I__7483\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30953\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__30956\,
            I => \N__30950\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__30953\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__30950\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__7479\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30937\
        );

    \I__7478\ : InMux
    port map (
            O => \N__30944\,
            I => \N__30937\
        );

    \I__7477\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30934\
        );

    \I__7476\ : InMux
    port map (
            O => \N__30942\,
            I => \N__30931\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__30937\,
            I => \N__30927\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__30934\,
            I => \N__30922\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__30931\,
            I => \N__30922\
        );

    \I__7472\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30919\
        );

    \I__7471\ : Span4Mux_v
    port map (
            O => \N__30927\,
            I => \N__30915\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__30922\,
            I => \N__30910\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__30919\,
            I => \N__30910\
        );

    \I__7468\ : InMux
    port map (
            O => \N__30918\,
            I => \N__30907\
        );

    \I__7467\ : Span4Mux_h
    port map (
            O => \N__30915\,
            I => \N__30902\
        );

    \I__7466\ : Span4Mux_v
    port map (
            O => \N__30910\,
            I => \N__30902\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__30907\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__30902\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__7463\ : CascadeMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__7462\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30891\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__7460\ : Span12Mux_v
    port map (
            O => \N__30888\,
            I => \N__30885\
        );

    \I__7459\ : Odrv12
    port map (
            O => \N__30885\,
            I => \this_ppu.un1_M_haddress_q_2_6\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__30882\,
            I => \N__30879\
        );

    \I__7457\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30876\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__30876\,
            I => \N__30873\
        );

    \I__7455\ : Span4Mux_v
    port map (
            O => \N__30873\,
            I => \N__30870\
        );

    \I__7454\ : Odrv4
    port map (
            O => \N__30870\,
            I => \M_this_data_tmp_qZ0Z_19\
        );

    \I__7453\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__30864\,
            I => \N__30861\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__7450\ : Odrv4
    port map (
            O => \N__30858\,
            I => \M_this_oam_ram_write_data_19\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__30855\,
            I => \N__30852\
        );

    \I__7448\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30849\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__30849\,
            I => \N__30846\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__30846\,
            I => \N__30843\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__30843\,
            I => \N__30837\
        );

    \I__7444\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30834\
        );

    \I__7443\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30831\
        );

    \I__7442\ : InMux
    port map (
            O => \N__30840\,
            I => \N__30828\
        );

    \I__7441\ : Span4Mux_h
    port map (
            O => \N__30837\,
            I => \N__30825\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__30834\,
            I => \N__30818\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__30831\,
            I => \N__30813\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__30828\,
            I => \N__30813\
        );

    \I__7437\ : Sp12to4
    port map (
            O => \N__30825\,
            I => \N__30809\
        );

    \I__7436\ : InMux
    port map (
            O => \N__30824\,
            I => \N__30802\
        );

    \I__7435\ : InMux
    port map (
            O => \N__30823\,
            I => \N__30802\
        );

    \I__7434\ : InMux
    port map (
            O => \N__30822\,
            I => \N__30802\
        );

    \I__7433\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30799\
        );

    \I__7432\ : Span4Mux_v
    port map (
            O => \N__30818\,
            I => \N__30794\
        );

    \I__7431\ : Span4Mux_h
    port map (
            O => \N__30813\,
            I => \N__30794\
        );

    \I__7430\ : InMux
    port map (
            O => \N__30812\,
            I => \N__30791\
        );

    \I__7429\ : Odrv12
    port map (
            O => \N__30809\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__30802\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__30799\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__30794\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__30791\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__7424\ : CascadeMux
    port map (
            O => \N__30780\,
            I => \N__30775\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__30779\,
            I => \N__30772\
        );

    \I__7422\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30769\
        );

    \I__7421\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30766\
        );

    \I__7420\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30762\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__30769\,
            I => \N__30759\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__30766\,
            I => \N__30756\
        );

    \I__7417\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30753\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__30762\,
            I => \N__30750\
        );

    \I__7415\ : Span4Mux_h
    port map (
            O => \N__30759\,
            I => \N__30747\
        );

    \I__7414\ : Span4Mux_h
    port map (
            O => \N__30756\,
            I => \N__30744\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__30753\,
            I => \N__30741\
        );

    \I__7412\ : Span4Mux_h
    port map (
            O => \N__30750\,
            I => \N__30738\
        );

    \I__7411\ : Span4Mux_v
    port map (
            O => \N__30747\,
            I => \N__30735\
        );

    \I__7410\ : Sp12to4
    port map (
            O => \N__30744\,
            I => \N__30732\
        );

    \I__7409\ : Span4Mux_v
    port map (
            O => \N__30741\,
            I => \N__30729\
        );

    \I__7408\ : Span4Mux_v
    port map (
            O => \N__30738\,
            I => \N__30726\
        );

    \I__7407\ : Span4Mux_v
    port map (
            O => \N__30735\,
            I => \N__30723\
        );

    \I__7406\ : Span12Mux_v
    port map (
            O => \N__30732\,
            I => \N__30720\
        );

    \I__7405\ : Span4Mux_v
    port map (
            O => \N__30729\,
            I => \N__30715\
        );

    \I__7404\ : Span4Mux_h
    port map (
            O => \N__30726\,
            I => \N__30715\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__30723\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__7402\ : Odrv12
    port map (
            O => \N__30720\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__30715\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__7400\ : CascadeMux
    port map (
            O => \N__30708\,
            I => \N__30705\
        );

    \I__7399\ : InMux
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__30702\,
            I => \this_ppu.M_this_oam_ram_read_data_i_16\
        );

    \I__7397\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30696\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__30696\,
            I => \N__30691\
        );

    \I__7395\ : CascadeMux
    port map (
            O => \N__30695\,
            I => \N__30687\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__30694\,
            I => \N__30684\
        );

    \I__7393\ : Span4Mux_v
    port map (
            O => \N__30691\,
            I => \N__30680\
        );

    \I__7392\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30677\
        );

    \I__7391\ : InMux
    port map (
            O => \N__30687\,
            I => \N__30671\
        );

    \I__7390\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30671\
        );

    \I__7389\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30668\
        );

    \I__7388\ : Sp12to4
    port map (
            O => \N__30680\,
            I => \N__30663\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__30677\,
            I => \N__30663\
        );

    \I__7386\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30660\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__30671\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__30668\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7383\ : Odrv12
    port map (
            O => \N__30663\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__30660\,
            I => \this_ppu.M_vaddress_qZ0Z_1\
        );

    \I__7381\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30648\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__30648\,
            I => \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\
        );

    \I__7379\ : InMux
    port map (
            O => \N__30645\,
            I => \this_ppu.un2_vscroll_cry_0\
        );

    \I__7378\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__7376\ : Span4Mux_v
    port map (
            O => \N__30636\,
            I => \N__30628\
        );

    \I__7375\ : InMux
    port map (
            O => \N__30635\,
            I => \N__30625\
        );

    \I__7374\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30617\
        );

    \I__7373\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30617\
        );

    \I__7372\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30617\
        );

    \I__7371\ : InMux
    port map (
            O => \N__30631\,
            I => \N__30614\
        );

    \I__7370\ : Sp12to4
    port map (
            O => \N__30628\,
            I => \N__30609\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__30625\,
            I => \N__30609\
        );

    \I__7368\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30606\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__30617\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__30614\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7365\ : Odrv12
    port map (
            O => \N__30609\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__30606\,
            I => \this_ppu.M_vaddress_qZ0Z_2\
        );

    \I__7363\ : CascadeMux
    port map (
            O => \N__30597\,
            I => \N__30594\
        );

    \I__7362\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__30591\,
            I => \N__30586\
        );

    \I__7360\ : CascadeMux
    port map (
            O => \N__30590\,
            I => \N__30583\
        );

    \I__7359\ : InMux
    port map (
            O => \N__30589\,
            I => \N__30580\
        );

    \I__7358\ : Span4Mux_v
    port map (
            O => \N__30586\,
            I => \N__30577\
        );

    \I__7357\ : InMux
    port map (
            O => \N__30583\,
            I => \N__30574\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__30580\,
            I => \N__30571\
        );

    \I__7355\ : Sp12to4
    port map (
            O => \N__30577\,
            I => \N__30566\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__30574\,
            I => \N__30566\
        );

    \I__7353\ : Span12Mux_v
    port map (
            O => \N__30571\,
            I => \N__30563\
        );

    \I__7352\ : Span12Mux_h
    port map (
            O => \N__30566\,
            I => \N__30560\
        );

    \I__7351\ : Odrv12
    port map (
            O => \N__30563\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__7350\ : Odrv12
    port map (
            O => \N__30560\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__7349\ : InMux
    port map (
            O => \N__30555\,
            I => \this_ppu.un2_vscroll_cry_1\
        );

    \I__7348\ : InMux
    port map (
            O => \N__30552\,
            I => \N__30549\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__30549\,
            I => \N__30546\
        );

    \I__7346\ : Odrv4
    port map (
            O => \N__30546\,
            I => \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\
        );

    \I__7345\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30537\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__7342\ : Span4Mux_v
    port map (
            O => \N__30534\,
            I => \N__30531\
        );

    \I__7341\ : Span4Mux_h
    port map (
            O => \N__30531\,
            I => \N__30528\
        );

    \I__7340\ : Sp12to4
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__7339\ : Span12Mux_h
    port map (
            O => \N__30525\,
            I => \N__30522\
        );

    \I__7338\ : Odrv12
    port map (
            O => \N__30522\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__7337\ : CascadeMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__7336\ : InMux
    port map (
            O => \N__30516\,
            I => \N__30511\
        );

    \I__7335\ : CascadeMux
    port map (
            O => \N__30515\,
            I => \N__30508\
        );

    \I__7334\ : CascadeMux
    port map (
            O => \N__30514\,
            I => \N__30504\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__30511\,
            I => \N__30501\
        );

    \I__7332\ : InMux
    port map (
            O => \N__30508\,
            I => \N__30498\
        );

    \I__7331\ : CascadeMux
    port map (
            O => \N__30507\,
            I => \N__30495\
        );

    \I__7330\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30490\
        );

    \I__7329\ : Span4Mux_h
    port map (
            O => \N__30501\,
            I => \N__30485\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__30498\,
            I => \N__30485\
        );

    \I__7327\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30482\
        );

    \I__7326\ : CascadeMux
    port map (
            O => \N__30494\,
            I => \N__30479\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__30493\,
            I => \N__30476\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__30490\,
            I => \N__30471\
        );

    \I__7323\ : Span4Mux_v
    port map (
            O => \N__30485\,
            I => \N__30466\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__30482\,
            I => \N__30466\
        );

    \I__7321\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30463\
        );

    \I__7320\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30460\
        );

    \I__7319\ : CascadeMux
    port map (
            O => \N__30475\,
            I => \N__30457\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__30474\,
            I => \N__30454\
        );

    \I__7317\ : Span4Mux_h
    port map (
            O => \N__30471\,
            I => \N__30449\
        );

    \I__7316\ : Span4Mux_v
    port map (
            O => \N__30466\,
            I => \N__30444\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__30463\,
            I => \N__30444\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__30460\,
            I => \N__30441\
        );

    \I__7313\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30438\
        );

    \I__7312\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30435\
        );

    \I__7311\ : CascadeMux
    port map (
            O => \N__30453\,
            I => \N__30432\
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__30452\,
            I => \N__30429\
        );

    \I__7309\ : Span4Mux_v
    port map (
            O => \N__30449\,
            I => \N__30420\
        );

    \I__7308\ : Span4Mux_h
    port map (
            O => \N__30444\,
            I => \N__30420\
        );

    \I__7307\ : Span4Mux_s1_v
    port map (
            O => \N__30441\,
            I => \N__30413\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30413\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__30435\,
            I => \N__30413\
        );

    \I__7304\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30410\
        );

    \I__7303\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30407\
        );

    \I__7302\ : CascadeMux
    port map (
            O => \N__30428\,
            I => \N__30404\
        );

    \I__7301\ : CascadeMux
    port map (
            O => \N__30427\,
            I => \N__30401\
        );

    \I__7300\ : CascadeMux
    port map (
            O => \N__30426\,
            I => \N__30398\
        );

    \I__7299\ : CascadeMux
    port map (
            O => \N__30425\,
            I => \N__30395\
        );

    \I__7298\ : Span4Mux_h
    port map (
            O => \N__30420\,
            I => \N__30391\
        );

    \I__7297\ : Span4Mux_v
    port map (
            O => \N__30413\,
            I => \N__30386\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__30410\,
            I => \N__30386\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30383\
        );

    \I__7294\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30380\
        );

    \I__7293\ : InMux
    port map (
            O => \N__30401\,
            I => \N__30377\
        );

    \I__7292\ : InMux
    port map (
            O => \N__30398\,
            I => \N__30374\
        );

    \I__7291\ : InMux
    port map (
            O => \N__30395\,
            I => \N__30371\
        );

    \I__7290\ : CascadeMux
    port map (
            O => \N__30394\,
            I => \N__30368\
        );

    \I__7289\ : Span4Mux_h
    port map (
            O => \N__30391\,
            I => \N__30364\
        );

    \I__7288\ : Span4Mux_v
    port map (
            O => \N__30386\,
            I => \N__30355\
        );

    \I__7287\ : Span4Mux_v
    port map (
            O => \N__30383\,
            I => \N__30355\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__30380\,
            I => \N__30355\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__30377\,
            I => \N__30355\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__30374\,
            I => \N__30350\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__30371\,
            I => \N__30350\
        );

    \I__7282\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30347\
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__30367\,
            I => \N__30344\
        );

    \I__7280\ : Span4Mux_h
    port map (
            O => \N__30364\,
            I => \N__30341\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__30355\,
            I => \N__30334\
        );

    \I__7278\ : Span4Mux_v
    port map (
            O => \N__30350\,
            I => \N__30334\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30334\
        );

    \I__7276\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30331\
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__30341\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__30334\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__30331\,
            I => \M_this_ppu_sprites_addr_10\
        );

    \I__7272\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30321\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__30321\,
            I => \N__30314\
        );

    \I__7270\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30311\
        );

    \I__7269\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30308\
        );

    \I__7268\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30303\
        );

    \I__7267\ : InMux
    port map (
            O => \N__30317\,
            I => \N__30303\
        );

    \I__7266\ : Span4Mux_v
    port map (
            O => \N__30314\,
            I => \N__30296\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__30311\,
            I => \N__30296\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__30308\,
            I => \N__30296\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__30303\,
            I => \N__30290\
        );

    \I__7262\ : Span4Mux_v
    port map (
            O => \N__30296\,
            I => \N__30287\
        );

    \I__7261\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30284\
        );

    \I__7260\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30281\
        );

    \I__7259\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30276\
        );

    \I__7258\ : Span4Mux_h
    port map (
            O => \N__30290\,
            I => \N__30273\
        );

    \I__7257\ : Sp12to4
    port map (
            O => \N__30287\,
            I => \N__30268\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__30284\,
            I => \N__30268\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__30281\,
            I => \N__30265\
        );

    \I__7254\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30262\
        );

    \I__7253\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30259\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__30276\,
            I => \N__30256\
        );

    \I__7251\ : Odrv4
    port map (
            O => \N__30273\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7250\ : Odrv12
    port map (
            O => \N__30268\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7249\ : Odrv4
    port map (
            O => \N__30265\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__30262\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__30259\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__30256\,
            I => \M_this_sprites_address_qZ0Z_11\
        );

    \I__7245\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30235\
        );

    \I__7244\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30232\
        );

    \I__7243\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30229\
        );

    \I__7242\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30226\
        );

    \I__7241\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30221\
        );

    \I__7240\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30221\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__30235\,
            I => \N__30216\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__30232\,
            I => \N__30213\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__30229\,
            I => \N__30208\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__30226\,
            I => \N__30208\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__30221\,
            I => \N__30205\
        );

    \I__7234\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30202\
        );

    \I__7233\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30199\
        );

    \I__7232\ : Span4Mux_h
    port map (
            O => \N__30216\,
            I => \N__30194\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__30213\,
            I => \N__30189\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__30208\,
            I => \N__30189\
        );

    \I__7229\ : Span12Mux_h
    port map (
            O => \N__30205\,
            I => \N__30184\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__30202\,
            I => \N__30184\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__30199\,
            I => \N__30181\
        );

    \I__7226\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30178\
        );

    \I__7225\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30175\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__30194\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7223\ : Odrv4
    port map (
            O => \N__30189\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7222\ : Odrv12
    port map (
            O => \N__30184\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__30181\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__30178\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__30175\,
            I => \M_this_sprites_address_qZ0Z_12\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__30162\,
            I => \N__30154\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__30161\,
            I => \N__30151\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__30160\,
            I => \N__30148\
        );

    \I__7215\ : CascadeMux
    port map (
            O => \N__30159\,
            I => \N__30145\
        );

    \I__7214\ : CascadeMux
    port map (
            O => \N__30158\,
            I => \N__30141\
        );

    \I__7213\ : CascadeMux
    port map (
            O => \N__30157\,
            I => \N__30138\
        );

    \I__7212\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30133\
        );

    \I__7211\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30133\
        );

    \I__7210\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30130\
        );

    \I__7209\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30127\
        );

    \I__7208\ : CascadeMux
    port map (
            O => \N__30144\,
            I => \N__30124\
        );

    \I__7207\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30120\
        );

    \I__7206\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30117\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__30133\,
            I => \N__30114\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__30130\,
            I => \N__30109\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30109\
        );

    \I__7202\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30106\
        );

    \I__7201\ : CascadeMux
    port map (
            O => \N__30123\,
            I => \N__30103\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__30120\,
            I => \N__30099\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__30117\,
            I => \N__30096\
        );

    \I__7198\ : Span4Mux_v
    port map (
            O => \N__30114\,
            I => \N__30093\
        );

    \I__7197\ : Span4Mux_v
    port map (
            O => \N__30109\,
            I => \N__30088\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__30106\,
            I => \N__30088\
        );

    \I__7195\ : InMux
    port map (
            O => \N__30103\,
            I => \N__30085\
        );

    \I__7194\ : InMux
    port map (
            O => \N__30102\,
            I => \N__30081\
        );

    \I__7193\ : Span4Mux_h
    port map (
            O => \N__30099\,
            I => \N__30076\
        );

    \I__7192\ : Span4Mux_h
    port map (
            O => \N__30096\,
            I => \N__30076\
        );

    \I__7191\ : Span4Mux_h
    port map (
            O => \N__30093\,
            I => \N__30071\
        );

    \I__7190\ : Span4Mux_h
    port map (
            O => \N__30088\,
            I => \N__30071\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__30085\,
            I => \N__30068\
        );

    \I__7188\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30065\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__30081\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__30076\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7185\ : Odrv4
    port map (
            O => \N__30071\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__30068\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__30065\,
            I => \M_this_sprites_address_qZ0Z_13\
        );

    \I__7182\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30044\
        );

    \I__7181\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30041\
        );

    \I__7180\ : InMux
    port map (
            O => \N__30052\,
            I => \N__30038\
        );

    \I__7179\ : InMux
    port map (
            O => \N__30051\,
            I => \N__30035\
        );

    \I__7178\ : InMux
    port map (
            O => \N__30050\,
            I => \N__30032\
        );

    \I__7177\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30029\
        );

    \I__7176\ : InMux
    port map (
            O => \N__30048\,
            I => \N__30024\
        );

    \I__7175\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30024\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__30044\,
            I => \N__30021\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__30041\,
            I => \N__30018\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__30038\,
            I => \N__30015\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__30035\,
            I => \N__30010\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__30010\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__30029\,
            I => \N__30007\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__30004\
        );

    \I__7167\ : Span4Mux_v
    port map (
            O => \N__30021\,
            I => \N__29999\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__30018\,
            I => \N__29999\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__30015\,
            I => \N__29990\
        );

    \I__7164\ : Span4Mux_v
    port map (
            O => \N__30010\,
            I => \N__29990\
        );

    \I__7163\ : Span4Mux_h
    port map (
            O => \N__30007\,
            I => \N__29990\
        );

    \I__7162\ : Span4Mux_h
    port map (
            O => \N__30004\,
            I => \N__29990\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__29999\,
            I => \N_23_0\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__29990\,
            I => \N_23_0\
        );

    \I__7159\ : CEMux
    port map (
            O => \N__29985\,
            I => \N__29981\
        );

    \I__7158\ : CEMux
    port map (
            O => \N__29984\,
            I => \N__29978\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__29981\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__29978\,
            I => \this_sprites_ram.mem_WE_2\
        );

    \I__7155\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29970\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29966\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \N__29962\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__29966\,
            I => \N__29958\
        );

    \I__7151\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29955\
        );

    \I__7150\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29952\
        );

    \I__7149\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29944\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__29958\,
            I => \N__29939\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__29955\,
            I => \N__29939\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29936\
        );

    \I__7145\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29931\
        );

    \I__7144\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29931\
        );

    \I__7143\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29924\
        );

    \I__7142\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29924\
        );

    \I__7141\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29924\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__29944\,
            I => \N__29921\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__29939\,
            I => \N__29918\
        );

    \I__7138\ : Span12Mux_h
    port map (
            O => \N__29936\,
            I => \N__29915\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29906\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__29924\,
            I => \N__29906\
        );

    \I__7135\ : Span4Mux_v
    port map (
            O => \N__29921\,
            I => \N__29906\
        );

    \I__7134\ : Span4Mux_v
    port map (
            O => \N__29918\,
            I => \N__29906\
        );

    \I__7133\ : Odrv12
    port map (
            O => \N__29915\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__29906\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__29901\,
            I => \N__29898\
        );

    \I__7130\ : InMux
    port map (
            O => \N__29898\,
            I => \N__29892\
        );

    \I__7129\ : CascadeMux
    port map (
            O => \N__29897\,
            I => \N__29889\
        );

    \I__7128\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29886\
        );

    \I__7127\ : InMux
    port map (
            O => \N__29895\,
            I => \N__29883\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__29892\,
            I => \N__29880\
        );

    \I__7125\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29877\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__29886\,
            I => \N__29874\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29871\
        );

    \I__7122\ : Span4Mux_h
    port map (
            O => \N__29880\,
            I => \N__29866\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__29877\,
            I => \N__29866\
        );

    \I__7120\ : Span12Mux_h
    port map (
            O => \N__29874\,
            I => \N__29863\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__29871\,
            I => \N__29858\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__29866\,
            I => \N__29858\
        );

    \I__7117\ : Span12Mux_v
    port map (
            O => \N__29863\,
            I => \N__29855\
        );

    \I__7116\ : Span4Mux_v
    port map (
            O => \N__29858\,
            I => \N__29852\
        );

    \I__7115\ : Odrv12
    port map (
            O => \N__29855\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__29852\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__7113\ : CascadeMux
    port map (
            O => \N__29847\,
            I => \N__29844\
        );

    \I__7112\ : InMux
    port map (
            O => \N__29844\,
            I => \N__29841\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__29841\,
            I => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\
        );

    \I__7110\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29833\
        );

    \I__7109\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29830\
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__29836\,
            I => \N__29827\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__29833\,
            I => \N__29821\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__29830\,
            I => \N__29821\
        );

    \I__7105\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29817\
        );

    \I__7104\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29814\
        );

    \I__7103\ : Span4Mux_h
    port map (
            O => \N__29821\,
            I => \N__29811\
        );

    \I__7102\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29808\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__29817\,
            I => \N__29805\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__29814\,
            I => \N__29801\
        );

    \I__7099\ : Span4Mux_h
    port map (
            O => \N__29811\,
            I => \N__29796\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__29808\,
            I => \N__29796\
        );

    \I__7097\ : Sp12to4
    port map (
            O => \N__29805\,
            I => \N__29793\
        );

    \I__7096\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29789\
        );

    \I__7095\ : Span4Mux_v
    port map (
            O => \N__29801\,
            I => \N__29784\
        );

    \I__7094\ : Span4Mux_v
    port map (
            O => \N__29796\,
            I => \N__29784\
        );

    \I__7093\ : Span12Mux_s10_v
    port map (
            O => \N__29793\,
            I => \N__29781\
        );

    \I__7092\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29778\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__29789\,
            I => \N__29773\
        );

    \I__7090\ : Span4Mux_v
    port map (
            O => \N__29784\,
            I => \N__29773\
        );

    \I__7089\ : Odrv12
    port map (
            O => \N__29781\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__29778\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__29773\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__7086\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29763\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__29763\,
            I => \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\
        );

    \I__7084\ : InMux
    port map (
            O => \N__29760\,
            I => \this_ppu.un2_hscroll_cry_0\
        );

    \I__7083\ : CascadeMux
    port map (
            O => \N__29757\,
            I => \N__29754\
        );

    \I__7082\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29750\
        );

    \I__7081\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29747\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__29750\,
            I => \N__29744\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__29747\,
            I => \N__29738\
        );

    \I__7078\ : Span4Mux_v
    port map (
            O => \N__29744\,
            I => \N__29735\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__29743\,
            I => \N__29731\
        );

    \I__7076\ : CascadeMux
    port map (
            O => \N__29742\,
            I => \N__29728\
        );

    \I__7075\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29723\
        );

    \I__7074\ : Sp12to4
    port map (
            O => \N__29738\,
            I => \N__29720\
        );

    \I__7073\ : Sp12to4
    port map (
            O => \N__29735\,
            I => \N__29717\
        );

    \I__7072\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29714\
        );

    \I__7071\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29707\
        );

    \I__7070\ : InMux
    port map (
            O => \N__29728\,
            I => \N__29707\
        );

    \I__7069\ : InMux
    port map (
            O => \N__29727\,
            I => \N__29707\
        );

    \I__7068\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29704\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29699\
        );

    \I__7066\ : Span12Mux_v
    port map (
            O => \N__29720\,
            I => \N__29699\
        );

    \I__7065\ : Span12Mux_h
    port map (
            O => \N__29717\,
            I => \N__29694\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__29714\,
            I => \N__29694\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__29707\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__29704\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7061\ : Odrv12
    port map (
            O => \N__29699\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__29694\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__7059\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29682\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__29682\,
            I => \N__29679\
        );

    \I__7057\ : Odrv4
    port map (
            O => \N__29679\,
            I => \M_this_oam_ram_write_data_30\
        );

    \I__7056\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29673\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__29673\,
            I => \this_sprites_ram.mem_out_bus5_1\
        );

    \I__7054\ : InMux
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__29667\,
            I => \N__29664\
        );

    \I__7052\ : Span4Mux_v
    port map (
            O => \N__29664\,
            I => \N__29661\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__29661\,
            I => \this_sprites_ram.mem_out_bus1_1\
        );

    \I__7050\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29653\
        );

    \I__7049\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29643\
        );

    \I__7048\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29643\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__29653\,
            I => \N__29640\
        );

    \I__7046\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29637\
        );

    \I__7045\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29634\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__29650\,
            I => \N__29624\
        );

    \I__7043\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29618\
        );

    \I__7042\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29618\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__29643\,
            I => \N__29611\
        );

    \I__7040\ : Span4Mux_v
    port map (
            O => \N__29640\,
            I => \N__29611\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__29637\,
            I => \N__29611\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29608\
        );

    \I__7037\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29605\
        );

    \I__7036\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29600\
        );

    \I__7035\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29600\
        );

    \I__7034\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29597\
        );

    \I__7033\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29594\
        );

    \I__7032\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29591\
        );

    \I__7031\ : InMux
    port map (
            O => \N__29627\,
            I => \N__29584\
        );

    \I__7030\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29584\
        );

    \I__7029\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29584\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__29618\,
            I => \N__29581\
        );

    \I__7027\ : Span4Mux_h
    port map (
            O => \N__29611\,
            I => \N__29574\
        );

    \I__7026\ : Span4Mux_v
    port map (
            O => \N__29608\,
            I => \N__29574\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__29605\,
            I => \N__29574\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__29600\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__29597\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__29594\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__29591\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__29584\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__29581\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7018\ : Odrv4
    port map (
            O => \N__29574\,
            I => \this_sprites_ram.mem_radregZ0Z_13\
        );

    \I__7017\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29556\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__29553\,
            I => \N__29550\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__29550\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\
        );

    \I__7013\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__7012\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29539\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__29543\,
            I => \N__29536\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__29542\,
            I => \N__29532\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__29539\,
            I => \N__29529\
        );

    \I__7008\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29526\
        );

    \I__7007\ : CascadeMux
    port map (
            O => \N__29535\,
            I => \N__29523\
        );

    \I__7006\ : InMux
    port map (
            O => \N__29532\,
            I => \N__29516\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__29529\,
            I => \N__29511\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29511\
        );

    \I__7003\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29508\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__29522\,
            I => \N__29504\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__29521\,
            I => \N__29500\
        );

    \I__7000\ : CascadeMux
    port map (
            O => \N__29520\,
            I => \N__29496\
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__29519\,
            I => \N__29493\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__29516\,
            I => \N__29484\
        );

    \I__6997\ : Span4Mux_v
    port map (
            O => \N__29511\,
            I => \N__29484\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__29508\,
            I => \N__29484\
        );

    \I__6995\ : CascadeMux
    port map (
            O => \N__29507\,
            I => \N__29481\
        );

    \I__6994\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29478\
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__29503\,
            I => \N__29475\
        );

    \I__6992\ : InMux
    port map (
            O => \N__29500\,
            I => \N__29471\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__29499\,
            I => \N__29468\
        );

    \I__6990\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29465\
        );

    \I__6989\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29462\
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__29492\,
            I => \N__29459\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__29491\,
            I => \N__29456\
        );

    \I__6986\ : Span4Mux_v
    port map (
            O => \N__29484\,
            I => \N__29452\
        );

    \I__6985\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29449\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__29478\,
            I => \N__29446\
        );

    \I__6983\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29443\
        );

    \I__6982\ : CascadeMux
    port map (
            O => \N__29474\,
            I => \N__29440\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__29471\,
            I => \N__29437\
        );

    \I__6980\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29434\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29429\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29429\
        );

    \I__6977\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29426\
        );

    \I__6976\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29423\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__29455\,
            I => \N__29420\
        );

    \I__6974\ : Sp12to4
    port map (
            O => \N__29452\,
            I => \N__29414\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__29449\,
            I => \N__29414\
        );

    \I__6972\ : Span4Mux_s3_v
    port map (
            O => \N__29446\,
            I => \N__29409\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__29443\,
            I => \N__29409\
        );

    \I__6970\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29406\
        );

    \I__6969\ : Span4Mux_v
    port map (
            O => \N__29437\,
            I => \N__29401\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__29434\,
            I => \N__29401\
        );

    \I__6967\ : Span4Mux_v
    port map (
            O => \N__29429\,
            I => \N__29394\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__29426\,
            I => \N__29394\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__29423\,
            I => \N__29394\
        );

    \I__6964\ : InMux
    port map (
            O => \N__29420\,
            I => \N__29391\
        );

    \I__6963\ : CascadeMux
    port map (
            O => \N__29419\,
            I => \N__29388\
        );

    \I__6962\ : Span12Mux_h
    port map (
            O => \N__29414\,
            I => \N__29385\
        );

    \I__6961\ : Span4Mux_v
    port map (
            O => \N__29409\,
            I => \N__29380\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__29406\,
            I => \N__29380\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__29401\,
            I => \N__29373\
        );

    \I__6958\ : Span4Mux_v
    port map (
            O => \N__29394\,
            I => \N__29373\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__29391\,
            I => \N__29373\
        );

    \I__6956\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29370\
        );

    \I__6955\ : Odrv12
    port map (
            O => \N__29385\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__29380\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__29373\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__29370\,
            I => \M_this_ppu_sprites_addr_2\
        );

    \I__6951\ : CEMux
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__29358\,
            I => \N__29355\
        );

    \I__6949\ : Span4Mux_v
    port map (
            O => \N__29355\,
            I => \N__29351\
        );

    \I__6948\ : CEMux
    port map (
            O => \N__29354\,
            I => \N__29348\
        );

    \I__6947\ : Odrv4
    port map (
            O => \N__29351\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__29348\,
            I => \this_sprites_ram.mem_WE_4\
        );

    \I__6945\ : CEMux
    port map (
            O => \N__29343\,
            I => \N__29339\
        );

    \I__6944\ : CEMux
    port map (
            O => \N__29342\,
            I => \N__29336\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29331\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__29336\,
            I => \N__29331\
        );

    \I__6941\ : Span4Mux_v
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__29328\,
            I => \this_sprites_ram.mem_WE_12\
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__29325\,
            I => \N__29320\
        );

    \I__6938\ : CascadeMux
    port map (
            O => \N__29324\,
            I => \N__29317\
        );

    \I__6937\ : CascadeMux
    port map (
            O => \N__29323\,
            I => \N__29312\
        );

    \I__6936\ : InMux
    port map (
            O => \N__29320\,
            I => \N__29309\
        );

    \I__6935\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29306\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__29316\,
            I => \N__29303\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__29315\,
            I => \N__29300\
        );

    \I__6932\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29294\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__29309\,
            I => \N__29291\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__29306\,
            I => \N__29288\
        );

    \I__6929\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29285\
        );

    \I__6928\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29281\
        );

    \I__6927\ : CascadeMux
    port map (
            O => \N__29299\,
            I => \N__29278\
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__29298\,
            I => \N__29274\
        );

    \I__6925\ : CascadeMux
    port map (
            O => \N__29297\,
            I => \N__29269\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__29294\,
            I => \N__29265\
        );

    \I__6923\ : Span4Mux_v
    port map (
            O => \N__29291\,
            I => \N__29258\
        );

    \I__6922\ : Span4Mux_h
    port map (
            O => \N__29288\,
            I => \N__29258\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29258\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__29284\,
            I => \N__29255\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__29281\,
            I => \N__29252\
        );

    \I__6918\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29249\
        );

    \I__6917\ : CascadeMux
    port map (
            O => \N__29277\,
            I => \N__29246\
        );

    \I__6916\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29243\
        );

    \I__6915\ : CascadeMux
    port map (
            O => \N__29273\,
            I => \N__29240\
        );

    \I__6914\ : CascadeMux
    port map (
            O => \N__29272\,
            I => \N__29237\
        );

    \I__6913\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29233\
        );

    \I__6912\ : CascadeMux
    port map (
            O => \N__29268\,
            I => \N__29230\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__29265\,
            I => \N__29224\
        );

    \I__6910\ : Span4Mux_v
    port map (
            O => \N__29258\,
            I => \N__29224\
        );

    \I__6909\ : InMux
    port map (
            O => \N__29255\,
            I => \N__29221\
        );

    \I__6908\ : Span4Mux_s3_v
    port map (
            O => \N__29252\,
            I => \N__29216\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__29249\,
            I => \N__29216\
        );

    \I__6906\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29213\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__29243\,
            I => \N__29210\
        );

    \I__6904\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29207\
        );

    \I__6903\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29204\
        );

    \I__6902\ : CascadeMux
    port map (
            O => \N__29236\,
            I => \N__29201\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29198\
        );

    \I__6900\ : InMux
    port map (
            O => \N__29230\,
            I => \N__29195\
        );

    \I__6899\ : CascadeMux
    port map (
            O => \N__29229\,
            I => \N__29192\
        );

    \I__6898\ : Sp12to4
    port map (
            O => \N__29224\,
            I => \N__29188\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29185\
        );

    \I__6896\ : Span4Mux_v
    port map (
            O => \N__29216\,
            I => \N__29180\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__29213\,
            I => \N__29180\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__29210\,
            I => \N__29173\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__29207\,
            I => \N__29173\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__29204\,
            I => \N__29173\
        );

    \I__6891\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29170\
        );

    \I__6890\ : Span4Mux_v
    port map (
            O => \N__29198\,
            I => \N__29165\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29165\
        );

    \I__6888\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29162\
        );

    \I__6887\ : CascadeMux
    port map (
            O => \N__29191\,
            I => \N__29159\
        );

    \I__6886\ : Span12Mux_h
    port map (
            O => \N__29188\,
            I => \N__29156\
        );

    \I__6885\ : Span12Mux_h
    port map (
            O => \N__29185\,
            I => \N__29153\
        );

    \I__6884\ : Span4Mux_v
    port map (
            O => \N__29180\,
            I => \N__29146\
        );

    \I__6883\ : Span4Mux_v
    port map (
            O => \N__29173\,
            I => \N__29146\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__29170\,
            I => \N__29146\
        );

    \I__6881\ : Span4Mux_v
    port map (
            O => \N__29165\,
            I => \N__29141\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__29162\,
            I => \N__29141\
        );

    \I__6879\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29138\
        );

    \I__6878\ : Odrv12
    port map (
            O => \N__29156\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6877\ : Odrv12
    port map (
            O => \N__29153\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__29146\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__29141\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__29138\,
            I => \M_this_ppu_sprites_addr_5\
        );

    \I__6873\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29122\
        );

    \I__6872\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29117\
        );

    \I__6871\ : InMux
    port map (
            O => \N__29125\,
            I => \N__29117\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__29122\,
            I => \N__29106\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__29117\,
            I => \N__29106\
        );

    \I__6868\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29101\
        );

    \I__6867\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29101\
        );

    \I__6866\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29098\
        );

    \I__6865\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29095\
        );

    \I__6864\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29092\
        );

    \I__6863\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29088\
        );

    \I__6862\ : Span4Mux_v
    port map (
            O => \N__29106\,
            I => \N__29078\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__29101\,
            I => \N__29078\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29078\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__29095\,
            I => \N__29078\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__29092\,
            I => \N__29075\
        );

    \I__6857\ : InMux
    port map (
            O => \N__29091\,
            I => \N__29072\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__29088\,
            I => \N__29068\
        );

    \I__6855\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29065\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__29078\,
            I => \N__29062\
        );

    \I__6853\ : Span4Mux_h
    port map (
            O => \N__29075\,
            I => \N__29057\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__29072\,
            I => \N__29057\
        );

    \I__6851\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29054\
        );

    \I__6850\ : Odrv12
    port map (
            O => \N__29068\,
            I => \N_809\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N_809\
        );

    \I__6848\ : Odrv4
    port map (
            O => \N__29062\,
            I => \N_809\
        );

    \I__6847\ : Odrv4
    port map (
            O => \N__29057\,
            I => \N_809\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__29054\,
            I => \N_809\
        );

    \I__6845\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__29040\,
            I => \N__29037\
        );

    \I__6843\ : Span4Mux_v
    port map (
            O => \N__29037\,
            I => \N__29034\
        );

    \I__6842\ : Odrv4
    port map (
            O => \N__29034\,
            I => \M_this_sprites_address_q_RNO_0Z0Z_5\
        );

    \I__6841\ : CascadeMux
    port map (
            O => \N__29031\,
            I => \N__29028\
        );

    \I__6840\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__29025\,
            I => \N_595\
        );

    \I__6838\ : CascadeMux
    port map (
            O => \N__29022\,
            I => \N__29013\
        );

    \I__6837\ : CascadeMux
    port map (
            O => \N__29021\,
            I => \N__29004\
        );

    \I__6836\ : CascadeMux
    port map (
            O => \N__29020\,
            I => \N__29000\
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__29019\,
            I => \N__28996\
        );

    \I__6834\ : InMux
    port map (
            O => \N__29018\,
            I => \N__28986\
        );

    \I__6833\ : InMux
    port map (
            O => \N__29017\,
            I => \N__28986\
        );

    \I__6832\ : InMux
    port map (
            O => \N__29016\,
            I => \N__28986\
        );

    \I__6831\ : InMux
    port map (
            O => \N__29013\,
            I => \N__28983\
        );

    \I__6830\ : InMux
    port map (
            O => \N__29012\,
            I => \N__28980\
        );

    \I__6829\ : InMux
    port map (
            O => \N__29011\,
            I => \N__28973\
        );

    \I__6828\ : InMux
    port map (
            O => \N__29010\,
            I => \N__28973\
        );

    \I__6827\ : InMux
    port map (
            O => \N__29009\,
            I => \N__28973\
        );

    \I__6826\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28968\
        );

    \I__6825\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28968\
        );

    \I__6824\ : InMux
    port map (
            O => \N__29004\,
            I => \N__28963\
        );

    \I__6823\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28963\
        );

    \I__6822\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28956\
        );

    \I__6821\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28956\
        );

    \I__6820\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28956\
        );

    \I__6819\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28951\
        );

    \I__6818\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28951\
        );

    \I__6817\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28948\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__28986\,
            I => \N__28943\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__28983\,
            I => \N__28938\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__28980\,
            I => \N__28933\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__28973\,
            I => \N__28933\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__28968\,
            I => \N__28928\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__28963\,
            I => \N__28928\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28921\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28921\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__28948\,
            I => \N__28921\
        );

    \I__6807\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28918\
        );

    \I__6806\ : CascadeMux
    port map (
            O => \N__28946\,
            I => \N__28915\
        );

    \I__6805\ : Span4Mux_v
    port map (
            O => \N__28943\,
            I => \N__28911\
        );

    \I__6804\ : InMux
    port map (
            O => \N__28942\,
            I => \N__28908\
        );

    \I__6803\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28905\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__28938\,
            I => \N__28894\
        );

    \I__6801\ : Span4Mux_h
    port map (
            O => \N__28933\,
            I => \N__28894\
        );

    \I__6800\ : Span4Mux_v
    port map (
            O => \N__28928\,
            I => \N__28894\
        );

    \I__6799\ : Span4Mux_v
    port map (
            O => \N__28921\,
            I => \N__28894\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__28918\,
            I => \N__28894\
        );

    \I__6797\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28891\
        );

    \I__6796\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28888\
        );

    \I__6795\ : Sp12to4
    port map (
            O => \N__28911\,
            I => \N__28881\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__28908\,
            I => \N__28881\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28881\
        );

    \I__6792\ : Span4Mux_h
    port map (
            O => \N__28894\,
            I => \N__28878\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N_383_0\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__28888\,
            I => \N_383_0\
        );

    \I__6789\ : Odrv12
    port map (
            O => \N__28881\,
            I => \N_383_0\
        );

    \I__6788\ : Odrv4
    port map (
            O => \N__28878\,
            I => \N_383_0\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__28869\,
            I => \N__28865\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__28868\,
            I => \N__28862\
        );

    \I__6785\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28855\
        );

    \I__6784\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28852\
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__28861\,
            I => \N__28849\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__28860\,
            I => \N__28846\
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__28859\,
            I => \N__28842\
        );

    \I__6780\ : CascadeMux
    port map (
            O => \N__28858\,
            I => \N__28839\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__28855\,
            I => \N__28834\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__28852\,
            I => \N__28831\
        );

    \I__6777\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28828\
        );

    \I__6776\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28825\
        );

    \I__6775\ : CascadeMux
    port map (
            O => \N__28845\,
            I => \N__28821\
        );

    \I__6774\ : InMux
    port map (
            O => \N__28842\,
            I => \N__28816\
        );

    \I__6773\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28813\
        );

    \I__6772\ : CascadeMux
    port map (
            O => \N__28838\,
            I => \N__28810\
        );

    \I__6771\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \N__28807\
        );

    \I__6770\ : Span4Mux_v
    port map (
            O => \N__28834\,
            I => \N__28798\
        );

    \I__6769\ : Span4Mux_h
    port map (
            O => \N__28831\,
            I => \N__28798\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28798\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__28825\,
            I => \N__28795\
        );

    \I__6766\ : CascadeMux
    port map (
            O => \N__28824\,
            I => \N__28792\
        );

    \I__6765\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28789\
        );

    \I__6764\ : CascadeMux
    port map (
            O => \N__28820\,
            I => \N__28786\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__28819\,
            I => \N__28783\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28778\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__28813\,
            I => \N__28778\
        );

    \I__6760\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28775\
        );

    \I__6759\ : InMux
    port map (
            O => \N__28807\,
            I => \N__28772\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__28806\,
            I => \N__28769\
        );

    \I__6757\ : CascadeMux
    port map (
            O => \N__28805\,
            I => \N__28766\
        );

    \I__6756\ : Span4Mux_v
    port map (
            O => \N__28798\,
            I => \N__28759\
        );

    \I__6755\ : Span4Mux_v
    port map (
            O => \N__28795\,
            I => \N__28759\
        );

    \I__6754\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28756\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28753\
        );

    \I__6752\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28750\
        );

    \I__6751\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28747\
        );

    \I__6750\ : Span4Mux_v
    port map (
            O => \N__28778\,
            I => \N__28740\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__28775\,
            I => \N__28740\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__28772\,
            I => \N__28740\
        );

    \I__6747\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28737\
        );

    \I__6746\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28734\
        );

    \I__6745\ : CascadeMux
    port map (
            O => \N__28765\,
            I => \N__28731\
        );

    \I__6744\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28727\
        );

    \I__6743\ : Sp12to4
    port map (
            O => \N__28759\,
            I => \N__28722\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__28756\,
            I => \N__28722\
        );

    \I__6741\ : Span4Mux_v
    port map (
            O => \N__28753\,
            I => \N__28715\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28715\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__28747\,
            I => \N__28715\
        );

    \I__6738\ : Span4Mux_v
    port map (
            O => \N__28740\,
            I => \N__28708\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__28737\,
            I => \N__28708\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__28734\,
            I => \N__28708\
        );

    \I__6735\ : InMux
    port map (
            O => \N__28731\,
            I => \N__28705\
        );

    \I__6734\ : CascadeMux
    port map (
            O => \N__28730\,
            I => \N__28702\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28698\
        );

    \I__6732\ : Span12Mux_h
    port map (
            O => \N__28722\,
            I => \N__28695\
        );

    \I__6731\ : Span4Mux_v
    port map (
            O => \N__28715\,
            I => \N__28688\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__28708\,
            I => \N__28688\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28688\
        );

    \I__6728\ : InMux
    port map (
            O => \N__28702\,
            I => \N__28685\
        );

    \I__6727\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28682\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__28698\,
            I => \N__28679\
        );

    \I__6725\ : Odrv12
    port map (
            O => \N__28695\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6724\ : Odrv4
    port map (
            O => \N__28688\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__28685\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__28682\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__28679\,
            I => \M_this_sprites_address_qZ0Z_5\
        );

    \I__6720\ : SRMux
    port map (
            O => \N__28668\,
            I => \N__28632\
        );

    \I__6719\ : SRMux
    port map (
            O => \N__28667\,
            I => \N__28632\
        );

    \I__6718\ : SRMux
    port map (
            O => \N__28666\,
            I => \N__28632\
        );

    \I__6717\ : SRMux
    port map (
            O => \N__28665\,
            I => \N__28632\
        );

    \I__6716\ : SRMux
    port map (
            O => \N__28664\,
            I => \N__28632\
        );

    \I__6715\ : SRMux
    port map (
            O => \N__28663\,
            I => \N__28632\
        );

    \I__6714\ : SRMux
    port map (
            O => \N__28662\,
            I => \N__28632\
        );

    \I__6713\ : SRMux
    port map (
            O => \N__28661\,
            I => \N__28632\
        );

    \I__6712\ : SRMux
    port map (
            O => \N__28660\,
            I => \N__28632\
        );

    \I__6711\ : SRMux
    port map (
            O => \N__28659\,
            I => \N__28632\
        );

    \I__6710\ : SRMux
    port map (
            O => \N__28658\,
            I => \N__28632\
        );

    \I__6709\ : SRMux
    port map (
            O => \N__28657\,
            I => \N__28632\
        );

    \I__6708\ : GlobalMux
    port map (
            O => \N__28632\,
            I => \N__28629\
        );

    \I__6707\ : gio2CtrlBuf
    port map (
            O => \N__28629\,
            I => \N_515_g\
        );

    \I__6706\ : CEMux
    port map (
            O => \N__28626\,
            I => \N__28622\
        );

    \I__6705\ : CEMux
    port map (
            O => \N__28625\,
            I => \N__28619\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__28622\,
            I => \N__28614\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__28619\,
            I => \N__28614\
        );

    \I__6702\ : Span4Mux_v
    port map (
            O => \N__28614\,
            I => \N__28611\
        );

    \I__6701\ : Odrv4
    port map (
            O => \N__28611\,
            I => \this_sprites_ram.mem_WE_0\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__6699\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28600\
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__28604\,
            I => \N__28597\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__28603\,
            I => \N__28594\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__28600\,
            I => \N__28588\
        );

    \I__6695\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28585\
        );

    \I__6694\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28582\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__28593\,
            I => \N__28579\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__28592\,
            I => \N__28575\
        );

    \I__6691\ : CascadeMux
    port map (
            O => \N__28591\,
            I => \N__28571\
        );

    \I__6690\ : Span4Mux_h
    port map (
            O => \N__28588\,
            I => \N__28565\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28565\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__28582\,
            I => \N__28562\
        );

    \I__6687\ : InMux
    port map (
            O => \N__28579\,
            I => \N__28559\
        );

    \I__6686\ : CascadeMux
    port map (
            O => \N__28578\,
            I => \N__28556\
        );

    \I__6685\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28551\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__28574\,
            I => \N__28548\
        );

    \I__6683\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28544\
        );

    \I__6682\ : CascadeMux
    port map (
            O => \N__28570\,
            I => \N__28541\
        );

    \I__6681\ : Span4Mux_v
    port map (
            O => \N__28565\,
            I => \N__28533\
        );

    \I__6680\ : Span4Mux_h
    port map (
            O => \N__28562\,
            I => \N__28533\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__28559\,
            I => \N__28533\
        );

    \I__6678\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28530\
        );

    \I__6677\ : CascadeMux
    port map (
            O => \N__28555\,
            I => \N__28527\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__28554\,
            I => \N__28524\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__28551\,
            I => \N__28521\
        );

    \I__6674\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28518\
        );

    \I__6673\ : CascadeMux
    port map (
            O => \N__28547\,
            I => \N__28515\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__28544\,
            I => \N__28511\
        );

    \I__6671\ : InMux
    port map (
            O => \N__28541\,
            I => \N__28508\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__28540\,
            I => \N__28505\
        );

    \I__6669\ : Span4Mux_v
    port map (
            O => \N__28533\,
            I => \N__28501\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__28530\,
            I => \N__28498\
        );

    \I__6667\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28495\
        );

    \I__6666\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28492\
        );

    \I__6665\ : Span4Mux_v
    port map (
            O => \N__28521\,
            I => \N__28487\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__28518\,
            I => \N__28487\
        );

    \I__6663\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28484\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__28514\,
            I => \N__28481\
        );

    \I__6661\ : Span4Mux_s3_v
    port map (
            O => \N__28511\,
            I => \N__28476\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__28508\,
            I => \N__28476\
        );

    \I__6659\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28473\
        );

    \I__6658\ : CascadeMux
    port map (
            O => \N__28504\,
            I => \N__28470\
        );

    \I__6657\ : Sp12to4
    port map (
            O => \N__28501\,
            I => \N__28466\
        );

    \I__6656\ : Sp12to4
    port map (
            O => \N__28498\,
            I => \N__28463\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__28495\,
            I => \N__28458\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__28492\,
            I => \N__28458\
        );

    \I__6653\ : Span4Mux_v
    port map (
            O => \N__28487\,
            I => \N__28453\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28453\
        );

    \I__6651\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28450\
        );

    \I__6650\ : Span4Mux_v
    port map (
            O => \N__28476\,
            I => \N__28445\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__28473\,
            I => \N__28445\
        );

    \I__6648\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28442\
        );

    \I__6647\ : CascadeMux
    port map (
            O => \N__28469\,
            I => \N__28439\
        );

    \I__6646\ : Span12Mux_h
    port map (
            O => \N__28466\,
            I => \N__28436\
        );

    \I__6645\ : Span12Mux_h
    port map (
            O => \N__28463\,
            I => \N__28433\
        );

    \I__6644\ : Span4Mux_v
    port map (
            O => \N__28458\,
            I => \N__28426\
        );

    \I__6643\ : Span4Mux_v
    port map (
            O => \N__28453\,
            I => \N__28426\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__28450\,
            I => \N__28426\
        );

    \I__6641\ : Span4Mux_v
    port map (
            O => \N__28445\,
            I => \N__28421\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__28442\,
            I => \N__28421\
        );

    \I__6639\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28418\
        );

    \I__6638\ : Odrv12
    port map (
            O => \N__28436\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__6637\ : Odrv12
    port map (
            O => \N__28433\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__28426\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__6635\ : Odrv4
    port map (
            O => \N__28421\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__28418\,
            I => \M_this_ppu_sprites_addr_4\
        );

    \I__6633\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__28404\,
            I => \N__28401\
        );

    \I__6631\ : Span4Mux_v
    port map (
            O => \N__28401\,
            I => \N__28398\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__28398\,
            I => \N_32_0\
        );

    \I__6629\ : CascadeMux
    port map (
            O => \N__28395\,
            I => \N__28392\
        );

    \I__6628\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28389\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28386\
        );

    \I__6626\ : Odrv4
    port map (
            O => \N__28386\,
            I => \M_this_data_tmp_qZ0Z_11\
        );

    \I__6625\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28380\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__28380\,
            I => \N__28377\
        );

    \I__6623\ : Odrv4
    port map (
            O => \N__28377\,
            I => \M_this_oam_ram_write_data_11\
        );

    \I__6622\ : CascadeMux
    port map (
            O => \N__28374\,
            I => \N__28371\
        );

    \I__6621\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__6619\ : Odrv4
    port map (
            O => \N__28365\,
            I => \M_this_data_tmp_qZ0Z_0\
        );

    \I__6618\ : InMux
    port map (
            O => \N__28362\,
            I => \N__28359\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__28359\,
            I => \N__28356\
        );

    \I__6616\ : Span4Mux_h
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__28353\,
            I => \N_748_0\
        );

    \I__6614\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28347\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__6612\ : Span4Mux_v
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__28341\,
            I => \N_44_0\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__28338\,
            I => \N__28335\
        );

    \I__6609\ : InMux
    port map (
            O => \N__28335\,
            I => \N__28332\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__28332\,
            I => \M_this_data_tmp_qZ0Z_17\
        );

    \I__6607\ : CEMux
    port map (
            O => \N__28329\,
            I => \N__28322\
        );

    \I__6606\ : CEMux
    port map (
            O => \N__28328\,
            I => \N__28319\
        );

    \I__6605\ : CEMux
    port map (
            O => \N__28327\,
            I => \N__28316\
        );

    \I__6604\ : CEMux
    port map (
            O => \N__28326\,
            I => \N__28313\
        );

    \I__6603\ : CEMux
    port map (
            O => \N__28325\,
            I => \N__28310\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__28322\,
            I => \N__28307\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__28319\,
            I => \N__28304\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__28316\,
            I => \N__28301\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__28313\,
            I => \N__28298\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__28310\,
            I => \N__28295\
        );

    \I__6597\ : Span4Mux_v
    port map (
            O => \N__28307\,
            I => \N__28292\
        );

    \I__6596\ : Span4Mux_v
    port map (
            O => \N__28304\,
            I => \N__28289\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__28301\,
            I => \N__28286\
        );

    \I__6594\ : Span4Mux_h
    port map (
            O => \N__28298\,
            I => \N__28283\
        );

    \I__6593\ : Span4Mux_v
    port map (
            O => \N__28295\,
            I => \N__28280\
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__28292\,
            I => \N_1174_0\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__28289\,
            I => \N_1174_0\
        );

    \I__6590\ : Odrv4
    port map (
            O => \N__28286\,
            I => \N_1174_0\
        );

    \I__6589\ : Odrv4
    port map (
            O => \N__28283\,
            I => \N_1174_0\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__28280\,
            I => \N_1174_0\
        );

    \I__6587\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__28266\,
            I => \N__28263\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__28263\,
            I => \M_this_data_tmp_qZ0Z_23\
        );

    \I__6584\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28254\
        );

    \I__6582\ : Span4Mux_h
    port map (
            O => \N__28254\,
            I => \N__28251\
        );

    \I__6581\ : Odrv4
    port map (
            O => \N__28251\,
            I => \M_this_oam_ram_write_data_23\
        );

    \I__6580\ : CascadeMux
    port map (
            O => \N__28248\,
            I => \N__28245\
        );

    \I__6579\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28242\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__28242\,
            I => \M_this_data_tmp_qZ0Z_20\
        );

    \I__6577\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28236\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__28233\,
            I => \N__28230\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__28230\,
            I => \N_42_0\
        );

    \I__6573\ : CascadeMux
    port map (
            O => \N__28227\,
            I => \N__28224\
        );

    \I__6572\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28221\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__28221\,
            I => \M_this_data_tmp_qZ0Z_8\
        );

    \I__6570\ : CEMux
    port map (
            O => \N__28218\,
            I => \N__28214\
        );

    \I__6569\ : CEMux
    port map (
            O => \N__28217\,
            I => \N__28210\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__28214\,
            I => \N__28207\
        );

    \I__6567\ : CEMux
    port map (
            O => \N__28213\,
            I => \N__28204\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28201\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__28207\,
            I => \N__28198\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28195\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__28201\,
            I => \N__28192\
        );

    \I__6562\ : Span4Mux_h
    port map (
            O => \N__28198\,
            I => \N__28187\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__28195\,
            I => \N__28187\
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__28192\,
            I => \N_1182_0\
        );

    \I__6559\ : Odrv4
    port map (
            O => \N__28187\,
            I => \N_1182_0\
        );

    \I__6558\ : CascadeMux
    port map (
            O => \N__28182\,
            I => \N__28179\
        );

    \I__6557\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28176\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__28176\,
            I => \M_this_data_tmp_qZ0Z_3\
        );

    \I__6555\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__6553\ : Span4Mux_h
    port map (
            O => \N__28167\,
            I => \N__28164\
        );

    \I__6552\ : Odrv4
    port map (
            O => \N__28164\,
            I => \N_745_0\
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__28161\,
            I => \N__28158\
        );

    \I__6550\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28155\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__28152\,
            I => \M_this_data_tmp_qZ0Z_14\
        );

    \I__6547\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28146\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__28146\,
            I => \N__28143\
        );

    \I__6545\ : Span4Mux_h
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__28140\,
            I => \N_739_0\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__6542\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__28131\,
            I => \N__28128\
        );

    \I__6540\ : Odrv4
    port map (
            O => \N__28128\,
            I => \M_this_data_tmp_qZ0Z_5\
        );

    \I__6539\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__28122\,
            I => \N__28119\
        );

    \I__6537\ : Span4Mux_h
    port map (
            O => \N__28119\,
            I => \N__28116\
        );

    \I__6536\ : Odrv4
    port map (
            O => \N__28116\,
            I => \N_743_0\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__28113\,
            I => \N_101_cascade_\
        );

    \I__6534\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28107\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__28107\,
            I => \N__28104\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__28104\,
            I => \M_this_sprites_address_q_RNO_0Z0Z_6\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__28101\,
            I => \N__28095\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__28100\,
            I => \N__28092\
        );

    \I__6529\ : CascadeMux
    port map (
            O => \N__28099\,
            I => \N__28087\
        );

    \I__6528\ : CascadeMux
    port map (
            O => \N__28098\,
            I => \N__28080\
        );

    \I__6527\ : InMux
    port map (
            O => \N__28095\,
            I => \N__28075\
        );

    \I__6526\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28072\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__28091\,
            I => \N__28069\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__28090\,
            I => \N__28066\
        );

    \I__6523\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28061\
        );

    \I__6522\ : CascadeMux
    port map (
            O => \N__28086\,
            I => \N__28058\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__28085\,
            I => \N__28055\
        );

    \I__6520\ : CascadeMux
    port map (
            O => \N__28084\,
            I => \N__28052\
        );

    \I__6519\ : CascadeMux
    port map (
            O => \N__28083\,
            I => \N__28049\
        );

    \I__6518\ : InMux
    port map (
            O => \N__28080\,
            I => \N__28046\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__28079\,
            I => \N__28043\
        );

    \I__6516\ : CascadeMux
    port map (
            O => \N__28078\,
            I => \N__28040\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__28075\,
            I => \N__28036\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__28072\,
            I => \N__28033\
        );

    \I__6513\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28030\
        );

    \I__6512\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28027\
        );

    \I__6511\ : CascadeMux
    port map (
            O => \N__28065\,
            I => \N__28024\
        );

    \I__6510\ : CascadeMux
    port map (
            O => \N__28064\,
            I => \N__28021\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__28061\,
            I => \N__28017\
        );

    \I__6508\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28014\
        );

    \I__6507\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28011\
        );

    \I__6506\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28008\
        );

    \I__6505\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28005\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__28002\
        );

    \I__6503\ : InMux
    port map (
            O => \N__28043\,
            I => \N__27999\
        );

    \I__6502\ : InMux
    port map (
            O => \N__28040\,
            I => \N__27996\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__28039\,
            I => \N__27993\
        );

    \I__6500\ : Span4Mux_v
    port map (
            O => \N__28036\,
            I => \N__27984\
        );

    \I__6499\ : Span4Mux_v
    port map (
            O => \N__28033\,
            I => \N__27984\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__28030\,
            I => \N__27984\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__28027\,
            I => \N__27984\
        );

    \I__6496\ : InMux
    port map (
            O => \N__28024\,
            I => \N__27981\
        );

    \I__6495\ : InMux
    port map (
            O => \N__28021\,
            I => \N__27978\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__28020\,
            I => \N__27975\
        );

    \I__6493\ : Span4Mux_v
    port map (
            O => \N__28017\,
            I => \N__27968\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__28014\,
            I => \N__27968\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__28011\,
            I => \N__27968\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__28008\,
            I => \N__27963\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__28005\,
            I => \N__27963\
        );

    \I__6488\ : Span4Mux_v
    port map (
            O => \N__28002\,
            I => \N__27956\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__27999\,
            I => \N__27956\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__27996\,
            I => \N__27956\
        );

    \I__6485\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27953\
        );

    \I__6484\ : Span4Mux_v
    port map (
            O => \N__27984\,
            I => \N__27946\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__27981\,
            I => \N__27946\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__27978\,
            I => \N__27946\
        );

    \I__6481\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27943\
        );

    \I__6480\ : Span4Mux_v
    port map (
            O => \N__27968\,
            I => \N__27938\
        );

    \I__6479\ : Span4Mux_v
    port map (
            O => \N__27963\,
            I => \N__27938\
        );

    \I__6478\ : Span4Mux_v
    port map (
            O => \N__27956\,
            I => \N__27929\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__27953\,
            I => \N__27929\
        );

    \I__6476\ : Span4Mux_v
    port map (
            O => \N__27946\,
            I => \N__27929\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__27943\,
            I => \N__27929\
        );

    \I__6474\ : Sp12to4
    port map (
            O => \N__27938\,
            I => \N__27925\
        );

    \I__6473\ : Span4Mux_v
    port map (
            O => \N__27929\,
            I => \N__27922\
        );

    \I__6472\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27918\
        );

    \I__6471\ : Span12Mux_h
    port map (
            O => \N__27925\,
            I => \N__27915\
        );

    \I__6470\ : Sp12to4
    port map (
            O => \N__27922\,
            I => \N__27912\
        );

    \I__6469\ : InMux
    port map (
            O => \N__27921\,
            I => \N__27909\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__27918\,
            I => \N__27906\
        );

    \I__6467\ : Odrv12
    port map (
            O => \N__27915\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__6466\ : Odrv12
    port map (
            O => \N__27912\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__27909\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__27906\,
            I => \M_this_sprites_address_qZ0Z_6\
        );

    \I__6463\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27894\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__27894\,
            I => \this_vga_signals.M_this_sprites_address_q_3_bmZ0Z_1\
        );

    \I__6461\ : CascadeMux
    port map (
            O => \N__27891\,
            I => \N__27881\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__27890\,
            I => \N__27878\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__27889\,
            I => \N__27873\
        );

    \I__6458\ : CascadeMux
    port map (
            O => \N__27888\,
            I => \N__27868\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__27887\,
            I => \N__27865\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__27886\,
            I => \N__27862\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__27885\,
            I => \N__27859\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__27884\,
            I => \N__27856\
        );

    \I__6453\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27852\
        );

    \I__6452\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27849\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__27877\,
            I => \N__27846\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__27876\,
            I => \N__27843\
        );

    \I__6449\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27839\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__27872\,
            I => \N__27836\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__27871\,
            I => \N__27833\
        );

    \I__6446\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27828\
        );

    \I__6445\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27825\
        );

    \I__6444\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27822\
        );

    \I__6443\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27819\
        );

    \I__6442\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27816\
        );

    \I__6441\ : CascadeMux
    port map (
            O => \N__27855\,
            I => \N__27813\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__27852\,
            I => \N__27810\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__27849\,
            I => \N__27807\
        );

    \I__6438\ : InMux
    port map (
            O => \N__27846\,
            I => \N__27804\
        );

    \I__6437\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27801\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__27842\,
            I => \N__27798\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__27839\,
            I => \N__27795\
        );

    \I__6434\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27792\
        );

    \I__6433\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27789\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__27832\,
            I => \N__27786\
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__27831\,
            I => \N__27783\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27776\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__27825\,
            I => \N__27776\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27776\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27771\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__27816\,
            I => \N__27771\
        );

    \I__6425\ : InMux
    port map (
            O => \N__27813\,
            I => \N__27767\
        );

    \I__6424\ : Span4Mux_v
    port map (
            O => \N__27810\,
            I => \N__27757\
        );

    \I__6423\ : Span4Mux_v
    port map (
            O => \N__27807\,
            I => \N__27757\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__27804\,
            I => \N__27757\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__27801\,
            I => \N__27757\
        );

    \I__6420\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27754\
        );

    \I__6419\ : Span4Mux_v
    port map (
            O => \N__27795\,
            I => \N__27747\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__27792\,
            I => \N__27747\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27747\
        );

    \I__6416\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27744\
        );

    \I__6415\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27741\
        );

    \I__6414\ : Span12Mux_v
    port map (
            O => \N__27776\,
            I => \N__27735\
        );

    \I__6413\ : Span12Mux_v
    port map (
            O => \N__27771\,
            I => \N__27735\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__27770\,
            I => \N__27732\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__27767\,
            I => \N__27729\
        );

    \I__6410\ : InMux
    port map (
            O => \N__27766\,
            I => \N__27726\
        );

    \I__6409\ : Span4Mux_v
    port map (
            O => \N__27757\,
            I => \N__27721\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__27754\,
            I => \N__27721\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__27747\,
            I => \N__27714\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__27744\,
            I => \N__27714\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27714\
        );

    \I__6404\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27711\
        );

    \I__6403\ : Span12Mux_h
    port map (
            O => \N__27735\,
            I => \N__27708\
        );

    \I__6402\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27705\
        );

    \I__6401\ : Span4Mux_h
    port map (
            O => \N__27729\,
            I => \N__27700\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27700\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__27721\,
            I => \N__27693\
        );

    \I__6398\ : Span4Mux_v
    port map (
            O => \N__27714\,
            I => \N__27693\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__27711\,
            I => \N__27693\
        );

    \I__6396\ : Odrv12
    port map (
            O => \N__27708\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__27705\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__6394\ : Odrv4
    port map (
            O => \N__27700\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__27693\,
            I => \M_this_sprites_address_qZ0Z_1\
        );

    \I__6392\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27673\
        );

    \I__6391\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27670\
        );

    \I__6390\ : InMux
    port map (
            O => \N__27682\,
            I => \N__27663\
        );

    \I__6389\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27658\
        );

    \I__6388\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27658\
        );

    \I__6387\ : InMux
    port map (
            O => \N__27679\,
            I => \N__27653\
        );

    \I__6386\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27653\
        );

    \I__6385\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27648\
        );

    \I__6384\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27648\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__27673\,
            I => \N__27643\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__27670\,
            I => \N__27643\
        );

    \I__6381\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27640\
        );

    \I__6380\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27637\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__27667\,
            I => \N__27633\
        );

    \I__6378\ : CascadeMux
    port map (
            O => \N__27666\,
            I => \N__27629\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__27663\,
            I => \N__27626\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__27658\,
            I => \N__27622\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__27653\,
            I => \N__27611\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__27648\,
            I => \N__27611\
        );

    \I__6373\ : Span4Mux_v
    port map (
            O => \N__27643\,
            I => \N__27611\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__27640\,
            I => \N__27611\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__27637\,
            I => \N__27611\
        );

    \I__6370\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27608\
        );

    \I__6369\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27604\
        );

    \I__6368\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27601\
        );

    \I__6367\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27598\
        );

    \I__6366\ : Span4Mux_v
    port map (
            O => \N__27626\,
            I => \N__27595\
        );

    \I__6365\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27592\
        );

    \I__6364\ : Span4Mux_v
    port map (
            O => \N__27622\,
            I => \N__27585\
        );

    \I__6363\ : Span4Mux_h
    port map (
            O => \N__27611\,
            I => \N__27585\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27585\
        );

    \I__6361\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27581\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27570\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__27601\,
            I => \N__27570\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__27598\,
            I => \N__27570\
        );

    \I__6357\ : Sp12to4
    port map (
            O => \N__27595\,
            I => \N__27570\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__27592\,
            I => \N__27570\
        );

    \I__6355\ : Span4Mux_h
    port map (
            O => \N__27585\,
            I => \N__27567\
        );

    \I__6354\ : InMux
    port map (
            O => \N__27584\,
            I => \N__27564\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__27581\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6352\ : Odrv12
    port map (
            O => \N__27570\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6351\ : Odrv4
    port map (
            O => \N__27567\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__27564\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__6349\ : InMux
    port map (
            O => \N__27555\,
            I => \N__27539\
        );

    \I__6348\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27533\
        );

    \I__6347\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27528\
        );

    \I__6346\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27528\
        );

    \I__6345\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27522\
        );

    \I__6344\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27522\
        );

    \I__6343\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27515\
        );

    \I__6342\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27511\
        );

    \I__6341\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27506\
        );

    \I__6340\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27506\
        );

    \I__6339\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27498\
        );

    \I__6338\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27498\
        );

    \I__6337\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27493\
        );

    \I__6336\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27493\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__27539\,
            I => \N__27490\
        );

    \I__6334\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27487\
        );

    \I__6333\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27484\
        );

    \I__6332\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27481\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__27533\,
            I => \N__27478\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27475\
        );

    \I__6329\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27472\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__27522\,
            I => \N__27469\
        );

    \I__6327\ : InMux
    port map (
            O => \N__27521\,
            I => \N__27466\
        );

    \I__6326\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27461\
        );

    \I__6325\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27461\
        );

    \I__6324\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27454\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__27515\,
            I => \N__27451\
        );

    \I__6322\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27448\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__27511\,
            I => \N__27443\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27443\
        );

    \I__6319\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27440\
        );

    \I__6318\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27435\
        );

    \I__6317\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27435\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__27498\,
            I => \N__27426\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__27493\,
            I => \N__27426\
        );

    \I__6314\ : Span4Mux_v
    port map (
            O => \N__27490\,
            I => \N__27426\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__27487\,
            I => \N__27426\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__27484\,
            I => \N__27423\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__27481\,
            I => \N__27420\
        );

    \I__6310\ : Span4Mux_h
    port map (
            O => \N__27478\,
            I => \N__27409\
        );

    \I__6309\ : Span4Mux_v
    port map (
            O => \N__27475\,
            I => \N__27409\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__27472\,
            I => \N__27409\
        );

    \I__6307\ : Span4Mux_v
    port map (
            O => \N__27469\,
            I => \N__27406\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__27466\,
            I => \N__27401\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__27461\,
            I => \N__27401\
        );

    \I__6304\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27394\
        );

    \I__6303\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27394\
        );

    \I__6302\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27394\
        );

    \I__6301\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27391\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27378\
        );

    \I__6299\ : Span4Mux_h
    port map (
            O => \N__27451\,
            I => \N__27378\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__27448\,
            I => \N__27378\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__27443\,
            I => \N__27378\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__27440\,
            I => \N__27378\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__27435\,
            I => \N__27378\
        );

    \I__6294\ : Span4Mux_h
    port map (
            O => \N__27426\,
            I => \N__27371\
        );

    \I__6293\ : Span4Mux_h
    port map (
            O => \N__27423\,
            I => \N__27371\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__27420\,
            I => \N__27371\
        );

    \I__6291\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27362\
        );

    \I__6290\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27362\
        );

    \I__6289\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27362\
        );

    \I__6288\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27362\
        );

    \I__6287\ : Odrv4
    port map (
            O => \N__27409\,
            I => \N_87_0\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__27406\,
            I => \N_87_0\
        );

    \I__6285\ : Odrv12
    port map (
            O => \N__27401\,
            I => \N_87_0\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__27394\,
            I => \N_87_0\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__27391\,
            I => \N_87_0\
        );

    \I__6282\ : Odrv4
    port map (
            O => \N__27378\,
            I => \N_87_0\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__27371\,
            I => \N_87_0\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N_87_0\
        );

    \I__6279\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27339\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__27339\,
            I => \this_vga_signals.M_this_sprites_address_q_3_amZ0Z_1\
        );

    \I__6276\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27333\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__27333\,
            I => \N__27330\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__27330\,
            I => \N__27324\
        );

    \I__6273\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27319\
        );

    \I__6272\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27319\
        );

    \I__6271\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27316\
        );

    \I__6270\ : Odrv4
    port map (
            O => \N__27324\,
            I => \this_vga_signals.un1_M_this_state_q_3_0_i_0_0\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__27319\,
            I => \this_vga_signals.un1_M_this_state_q_3_0_i_0_0\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__27316\,
            I => \this_vga_signals.un1_M_this_state_q_3_0_i_0_0\
        );

    \I__6267\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27306\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__27306\,
            I => \N__27302\
        );

    \I__6265\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27299\
        );

    \I__6264\ : Span4Mux_h
    port map (
            O => \N__27302\,
            I => \N__27293\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__27299\,
            I => \N__27290\
        );

    \I__6262\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27283\
        );

    \I__6261\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27283\
        );

    \I__6260\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27283\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__27293\,
            I => \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__27290\,
            I => \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__27283\,
            I => \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2\
        );

    \I__6256\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27270\
        );

    \I__6255\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27266\
        );

    \I__6254\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27263\
        );

    \I__6253\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27259\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__27270\,
            I => \N__27256\
        );

    \I__6251\ : InMux
    port map (
            O => \N__27269\,
            I => \N__27253\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27246\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27246\
        );

    \I__6248\ : InMux
    port map (
            O => \N__27262\,
            I => \N__27243\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__27259\,
            I => \N__27240\
        );

    \I__6246\ : Span4Mux_h
    port map (
            O => \N__27256\,
            I => \N__27237\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__27253\,
            I => \N__27234\
        );

    \I__6244\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27231\
        );

    \I__6243\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27228\
        );

    \I__6242\ : Span12Mux_v
    port map (
            O => \N__27246\,
            I => \N__27223\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__27243\,
            I => \N__27223\
        );

    \I__6240\ : Span12Mux_h
    port map (
            O => \N__27240\,
            I => \N__27220\
        );

    \I__6239\ : Span4Mux_v
    port map (
            O => \N__27237\,
            I => \N__27217\
        );

    \I__6238\ : Span4Mux_h
    port map (
            O => \N__27234\,
            I => \N__27214\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__27231\,
            I => \N__27211\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__27228\,
            I => \N__27208\
        );

    \I__6235\ : Span12Mux_h
    port map (
            O => \N__27223\,
            I => \N__27203\
        );

    \I__6234\ : Span12Mux_v
    port map (
            O => \N__27220\,
            I => \N__27203\
        );

    \I__6233\ : Span4Mux_v
    port map (
            O => \N__27217\,
            I => \N__27200\
        );

    \I__6232\ : Span4Mux_v
    port map (
            O => \N__27214\,
            I => \N__27193\
        );

    \I__6231\ : Span4Mux_h
    port map (
            O => \N__27211\,
            I => \N__27193\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__27208\,
            I => \N__27193\
        );

    \I__6229\ : Odrv12
    port map (
            O => \N__27203\,
            I => \M_this_sprites_ram_write_data_iv_i_i_3\
        );

    \I__6228\ : Odrv4
    port map (
            O => \N__27200\,
            I => \M_this_sprites_ram_write_data_iv_i_i_3\
        );

    \I__6227\ : Odrv4
    port map (
            O => \N__27193\,
            I => \M_this_sprites_ram_write_data_iv_i_i_3\
        );

    \I__6226\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__27183\,
            I => \this_ppu.un2_vscroll_axb_0\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27176\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__27179\,
            I => \N__27173\
        );

    \I__6222\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27168\
        );

    \I__6221\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27165\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__27172\,
            I => \N__27162\
        );

    \I__6219\ : CascadeMux
    port map (
            O => \N__27171\,
            I => \N__27156\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__27168\,
            I => \N__27151\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__27165\,
            I => \N__27151\
        );

    \I__6216\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27148\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__27161\,
            I => \N__27145\
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__27160\,
            I => \N__27141\
        );

    \I__6213\ : CascadeMux
    port map (
            O => \N__27159\,
            I => \N__27138\
        );

    \I__6212\ : InMux
    port map (
            O => \N__27156\,
            I => \N__27134\
        );

    \I__6211\ : Span4Mux_s2_v
    port map (
            O => \N__27151\,
            I => \N__27129\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__27148\,
            I => \N__27129\
        );

    \I__6209\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27126\
        );

    \I__6208\ : CascadeMux
    port map (
            O => \N__27144\,
            I => \N__27123\
        );

    \I__6207\ : InMux
    port map (
            O => \N__27141\,
            I => \N__27119\
        );

    \I__6206\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27116\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__27137\,
            I => \N__27113\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__27134\,
            I => \N__27110\
        );

    \I__6203\ : Span4Mux_v
    port map (
            O => \N__27129\,
            I => \N__27105\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__27126\,
            I => \N__27105\
        );

    \I__6201\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27102\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__27122\,
            I => \N__27099\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__27119\,
            I => \N__27094\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__27116\,
            I => \N__27091\
        );

    \I__6197\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27088\
        );

    \I__6196\ : Span4Mux_h
    port map (
            O => \N__27110\,
            I => \N__27085\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__27105\,
            I => \N__27080\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__27102\,
            I => \N__27080\
        );

    \I__6193\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27077\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__27098\,
            I => \N__27074\
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__27097\,
            I => \N__27070\
        );

    \I__6190\ : Span4Mux_h
    port map (
            O => \N__27094\,
            I => \N__27067\
        );

    \I__6189\ : Span4Mux_v
    port map (
            O => \N__27091\,
            I => \N__27062\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__27088\,
            I => \N__27062\
        );

    \I__6187\ : Span4Mux_h
    port map (
            O => \N__27085\,
            I => \N__27058\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__27080\,
            I => \N__27053\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__27077\,
            I => \N__27053\
        );

    \I__6184\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27050\
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__27073\,
            I => \N__27047\
        );

    \I__6182\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27043\
        );

    \I__6181\ : Span4Mux_v
    port map (
            O => \N__27067\,
            I => \N__27038\
        );

    \I__6180\ : Span4Mux_h
    port map (
            O => \N__27062\,
            I => \N__27038\
        );

    \I__6179\ : CascadeMux
    port map (
            O => \N__27061\,
            I => \N__27035\
        );

    \I__6178\ : Span4Mux_h
    port map (
            O => \N__27058\,
            I => \N__27032\
        );

    \I__6177\ : Span4Mux_h
    port map (
            O => \N__27053\,
            I => \N__27027\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__27050\,
            I => \N__27027\
        );

    \I__6175\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27024\
        );

    \I__6174\ : CascadeMux
    port map (
            O => \N__27046\,
            I => \N__27021\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__27043\,
            I => \N__27017\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__27038\,
            I => \N__27014\
        );

    \I__6171\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27011\
        );

    \I__6170\ : Span4Mux_h
    port map (
            O => \N__27032\,
            I => \N__27004\
        );

    \I__6169\ : Span4Mux_v
    port map (
            O => \N__27027\,
            I => \N__27004\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27004\
        );

    \I__6167\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27001\
        );

    \I__6166\ : CascadeMux
    port map (
            O => \N__27020\,
            I => \N__26998\
        );

    \I__6165\ : Span12Mux_h
    port map (
            O => \N__27017\,
            I => \N__26995\
        );

    \I__6164\ : Sp12to4
    port map (
            O => \N__27014\,
            I => \N__26992\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__27011\,
            I => \N__26989\
        );

    \I__6162\ : Span4Mux_h
    port map (
            O => \N__27004\,
            I => \N__26984\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__27001\,
            I => \N__26984\
        );

    \I__6160\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26981\
        );

    \I__6159\ : Span12Mux_v
    port map (
            O => \N__26995\,
            I => \N__26978\
        );

    \I__6158\ : Span12Mux_h
    port map (
            O => \N__26992\,
            I => \N__26975\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__26989\,
            I => \N__26968\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__26984\,
            I => \N__26968\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__26981\,
            I => \N__26968\
        );

    \I__6154\ : Odrv12
    port map (
            O => \N__26978\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__6153\ : Odrv12
    port map (
            O => \N__26975\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__6152\ : Odrv4
    port map (
            O => \N__26968\,
            I => \M_this_ppu_sprites_addr_1\
        );

    \I__6151\ : CascadeMux
    port map (
            O => \N__26961\,
            I => \N__26958\
        );

    \I__6150\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26955\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__26955\,
            I => \M_this_data_tmp_qZ0Z_4\
        );

    \I__6148\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26949\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__26949\,
            I => \N__26946\
        );

    \I__6146\ : Span4Mux_v
    port map (
            O => \N__26946\,
            I => \N__26943\
        );

    \I__6145\ : Odrv4
    port map (
            O => \N__26943\,
            I => \N_744_0\
        );

    \I__6144\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__26934\,
            I => \M_this_data_tmp_qZ0Z_7\
        );

    \I__6141\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26928\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26925\
        );

    \I__6139\ : Span4Mux_h
    port map (
            O => \N__26925\,
            I => \N__26922\
        );

    \I__6138\ : Odrv4
    port map (
            O => \N__26922\,
            I => \N_56_0\
        );

    \I__6137\ : CascadeMux
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__6136\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26913\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__26913\,
            I => \M_this_data_tmp_qZ0Z_16\
        );

    \I__6134\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26907\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__6132\ : Span4Mux_h
    port map (
            O => \N__26904\,
            I => \N__26901\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__26901\,
            I => \N_738_0\
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__6129\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__26892\,
            I => \M_this_data_tmp_qZ0Z_22\
        );

    \I__6127\ : InMux
    port map (
            O => \N__26889\,
            I => \N__26886\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26883\
        );

    \I__6125\ : Span4Mux_h
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__6124\ : Odrv4
    port map (
            O => \N__26880\,
            I => \N_40_0\
        );

    \I__6123\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26874\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__26874\,
            I => \N__26871\
        );

    \I__6121\ : Span4Mux_h
    port map (
            O => \N__26871\,
            I => \N__26868\
        );

    \I__6120\ : Span4Mux_v
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__6119\ : Odrv4
    port map (
            O => \N__26865\,
            I => \this_sprites_ram.mem_out_bus6_0\
        );

    \I__6118\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__6116\ : Span4Mux_v
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__26853\,
            I => \this_sprites_ram.mem_out_bus2_0\
        );

    \I__6114\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__26847\,
            I => \N__26844\
        );

    \I__6112\ : Odrv12
    port map (
            O => \N__26844\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__26841\,
            I => \N__26838\
        );

    \I__6110\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__26835\,
            I => \N_102\
        );

    \I__6108\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__26829\,
            I => \N__26826\
        );

    \I__6106\ : Odrv4
    port map (
            O => \N__26826\,
            I => \M_this_sprites_address_q_RNO_0Z0Z_4\
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__26823\,
            I => \N__26817\
        );

    \I__6104\ : CascadeMux
    port map (
            O => \N__26822\,
            I => \N__26812\
        );

    \I__6103\ : CascadeMux
    port map (
            O => \N__26821\,
            I => \N__26805\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__26820\,
            I => \N__26802\
        );

    \I__6101\ : InMux
    port map (
            O => \N__26817\,
            I => \N__26797\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__26816\,
            I => \N__26794\
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__26815\,
            I => \N__26791\
        );

    \I__6098\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26787\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__26811\,
            I => \N__26784\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__26810\,
            I => \N__26781\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__26809\,
            I => \N__26778\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__26808\,
            I => \N__26775\
        );

    \I__6093\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26772\
        );

    \I__6092\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26769\
        );

    \I__6091\ : CascadeMux
    port map (
            O => \N__26801\,
            I => \N__26766\
        );

    \I__6090\ : CascadeMux
    port map (
            O => \N__26800\,
            I => \N__26763\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__26797\,
            I => \N__26760\
        );

    \I__6088\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26757\
        );

    \I__6087\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26754\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__26790\,
            I => \N__26751\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__26787\,
            I => \N__26745\
        );

    \I__6084\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26742\
        );

    \I__6083\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26739\
        );

    \I__6082\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26736\
        );

    \I__6081\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26733\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__26772\,
            I => \N__26728\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__26769\,
            I => \N__26728\
        );

    \I__6078\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26725\
        );

    \I__6077\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26722\
        );

    \I__6076\ : Span4Mux_v
    port map (
            O => \N__26760\,
            I => \N__26715\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__26757\,
            I => \N__26715\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26715\
        );

    \I__6073\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26712\
        );

    \I__6072\ : CascadeMux
    port map (
            O => \N__26750\,
            I => \N__26709\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__26749\,
            I => \N__26706\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__26748\,
            I => \N__26703\
        );

    \I__6069\ : Span4Mux_v
    port map (
            O => \N__26745\,
            I => \N__26698\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26698\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__26739\,
            I => \N__26695\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26690\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__26733\,
            I => \N__26690\
        );

    \I__6064\ : Span4Mux_v
    port map (
            O => \N__26728\,
            I => \N__26683\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__26725\,
            I => \N__26683\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__26722\,
            I => \N__26683\
        );

    \I__6061\ : Span4Mux_v
    port map (
            O => \N__26715\,
            I => \N__26678\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__26712\,
            I => \N__26678\
        );

    \I__6059\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26675\
        );

    \I__6058\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26672\
        );

    \I__6057\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26669\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__26698\,
            I => \N__26662\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__26695\,
            I => \N__26662\
        );

    \I__6054\ : Span4Mux_v
    port map (
            O => \N__26690\,
            I => \N__26662\
        );

    \I__6053\ : Span4Mux_v
    port map (
            O => \N__26683\,
            I => \N__26655\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__26678\,
            I => \N__26655\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__26675\,
            I => \N__26655\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__26672\,
            I => \N__26651\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__26669\,
            I => \N__26648\
        );

    \I__6048\ : Sp12to4
    port map (
            O => \N__26662\,
            I => \N__26644\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__26655\,
            I => \N__26641\
        );

    \I__6046\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26638\
        );

    \I__6045\ : Span4Mux_h
    port map (
            O => \N__26651\,
            I => \N__26633\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__26648\,
            I => \N__26633\
        );

    \I__6043\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26630\
        );

    \I__6042\ : Span12Mux_h
    port map (
            O => \N__26644\,
            I => \N__26623\
        );

    \I__6041\ : Sp12to4
    port map (
            O => \N__26641\,
            I => \N__26623\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__26638\,
            I => \N__26623\
        );

    \I__6039\ : Odrv4
    port map (
            O => \N__26633\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__26630\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__6037\ : Odrv12
    port map (
            O => \N__26623\,
            I => \M_this_sprites_address_qZ0Z_4\
        );

    \I__6036\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__6034\ : Span4Mux_h
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__6033\ : Sp12to4
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__6032\ : Span12Mux_v
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__6031\ : Odrv12
    port map (
            O => \N__26601\,
            I => port_address_in_3
        );

    \I__6030\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__6028\ : Span12Mux_v
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__6027\ : Odrv12
    port map (
            O => \N__26589\,
            I => port_address_in_2
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__26586\,
            I => \N__26583\
        );

    \I__6025\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__26580\,
            I => \N__26577\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__26574\,
            I => \N__26571\
        );

    \I__6021\ : Sp12to4
    port map (
            O => \N__26571\,
            I => \N__26568\
        );

    \I__6020\ : Span12Mux_h
    port map (
            O => \N__26568\,
            I => \N__26564\
        );

    \I__6019\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26561\
        );

    \I__6018\ : Odrv12
    port map (
            O => \N__26564\,
            I => port_rw_in
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__26561\,
            I => port_rw_in
        );

    \I__6016\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26553\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__26553\,
            I => \N__26550\
        );

    \I__6014\ : Span4Mux_v
    port map (
            O => \N__26550\,
            I => \N__26547\
        );

    \I__6013\ : Sp12to4
    port map (
            O => \N__26547\,
            I => \N__26544\
        );

    \I__6012\ : Odrv12
    port map (
            O => \N__26544\,
            I => port_address_in_6
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__26541\,
            I => \N__26537\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__26540\,
            I => \N__26534\
        );

    \I__6009\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26529\
        );

    \I__6008\ : InMux
    port map (
            O => \N__26534\,
            I => \N__26529\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__26529\,
            I => \N__26526\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__26526\,
            I => \N__26523\
        );

    \I__6005\ : Span4Mux_h
    port map (
            O => \N__26523\,
            I => \N__26520\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__26520\,
            I => \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_4_0\
        );

    \I__6003\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26514\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__26511\,
            I => \N__26508\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__26508\,
            I => \N_54_0\
        );

    \I__5999\ : InMux
    port map (
            O => \N__26505\,
            I => \N__26502\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__26502\,
            I => \this_ppu.un1_oam_data_1_c2\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__26499\,
            I => \N__26493\
        );

    \I__5996\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26484\
        );

    \I__5995\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26484\
        );

    \I__5994\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26484\
        );

    \I__5993\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26480\
        );

    \I__5992\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26475\
        );

    \I__5991\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26475\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__26484\,
            I => \N__26472\
        );

    \I__5989\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26469\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__26480\,
            I => \N__26466\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__26475\,
            I => \N__26463\
        );

    \I__5986\ : Span4Mux_h
    port map (
            O => \N__26472\,
            I => \N__26458\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__26469\,
            I => \N__26458\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__26466\,
            I => \N__26455\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__26463\,
            I => \N__26450\
        );

    \I__5982\ : Span4Mux_v
    port map (
            O => \N__26458\,
            I => \N__26450\
        );

    \I__5981\ : Odrv4
    port map (
            O => \N__26455\,
            I => \N_163\
        );

    \I__5980\ : Odrv4
    port map (
            O => \N__26450\,
            I => \N_163\
        );

    \I__5979\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__26442\,
            I => \N__26438\
        );

    \I__5977\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26434\
        );

    \I__5976\ : Span4Mux_v
    port map (
            O => \N__26438\,
            I => \N__26431\
        );

    \I__5975\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26428\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__26434\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__26431\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__26428\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__5971\ : CascadeMux
    port map (
            O => \N__26421\,
            I => \N__26418\
        );

    \I__5970\ : CascadeBuf
    port map (
            O => \N__26418\,
            I => \N__26415\
        );

    \I__5969\ : CascadeMux
    port map (
            O => \N__26415\,
            I => \N__26412\
        );

    \I__5968\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26408\
        );

    \I__5967\ : InMux
    port map (
            O => \N__26411\,
            I => \N__26403\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__26408\,
            I => \N__26400\
        );

    \I__5965\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26397\
        );

    \I__5964\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26394\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__26403\,
            I => \N__26389\
        );

    \I__5962\ : Span12Mux_s11_v
    port map (
            O => \N__26400\,
            I => \N__26389\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__26397\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__26394\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5959\ : Odrv12
    port map (
            O => \N__26389\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__5958\ : CEMux
    port map (
            O => \N__26382\,
            I => \N__26378\
        );

    \I__5957\ : CEMux
    port map (
            O => \N__26381\,
            I => \N__26375\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__26378\,
            I => \N__26371\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26368\
        );

    \I__5954\ : CEMux
    port map (
            O => \N__26374\,
            I => \N__26365\
        );

    \I__5953\ : Span4Mux_v
    port map (
            O => \N__26371\,
            I => \N__26358\
        );

    \I__5952\ : Span4Mux_v
    port map (
            O => \N__26368\,
            I => \N__26358\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__26365\,
            I => \N__26358\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__26358\,
            I => \N__26355\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__26355\,
            I => \N_1190_0\
        );

    \I__5948\ : CascadeMux
    port map (
            O => \N__26352\,
            I => \N__26349\
        );

    \I__5947\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26346\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__26346\,
            I => \M_this_data_tmp_qZ0Z_6\
        );

    \I__5945\ : InMux
    port map (
            O => \N__26343\,
            I => \N__26340\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__5943\ : Span4Mux_h
    port map (
            O => \N__26337\,
            I => \N__26334\
        );

    \I__5942\ : Odrv4
    port map (
            O => \N__26334\,
            I => \N_742_0\
        );

    \I__5941\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26328\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__26328\,
            I => \N__26325\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__26325\,
            I => \N__26322\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__26322\,
            I => \N__26319\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__26319\,
            I => \N_34_0\
        );

    \I__5936\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26313\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__26313\,
            I => \M_this_sprites_address_q_RNO_0Z0Z_2\
        );

    \I__5934\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26305\
        );

    \I__5933\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26302\
        );

    \I__5932\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26299\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__26305\,
            I => \N__26293\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__26302\,
            I => \N__26293\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__26299\,
            I => \N__26290\
        );

    \I__5928\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26287\
        );

    \I__5927\ : Span4Mux_h
    port map (
            O => \N__26293\,
            I => \N__26282\
        );

    \I__5926\ : Span4Mux_v
    port map (
            O => \N__26290\,
            I => \N__26279\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26276\
        );

    \I__5924\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26273\
        );

    \I__5923\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26270\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__26282\,
            I => \N_813\
        );

    \I__5921\ : Odrv4
    port map (
            O => \N__26279\,
            I => \N_813\
        );

    \I__5920\ : Odrv12
    port map (
            O => \N__26276\,
            I => \N_813\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__26273\,
            I => \N_813\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N_813\
        );

    \I__5917\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26256\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__26256\,
            I => \N__26253\
        );

    \I__5915\ : Span4Mux_v
    port map (
            O => \N__26253\,
            I => \N__26250\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__26250\,
            I => \N_799\
        );

    \I__5913\ : CascadeMux
    port map (
            O => \N__26247\,
            I => \M_this_sprites_address_qc_11_0_cascade_\
        );

    \I__5912\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26241\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__26241\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_9\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \N__26234\
        );

    \I__5909\ : CascadeMux
    port map (
            O => \N__26237\,
            I => \N__26231\
        );

    \I__5908\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26224\
        );

    \I__5907\ : InMux
    port map (
            O => \N__26231\,
            I => \N__26221\
        );

    \I__5906\ : CascadeMux
    port map (
            O => \N__26230\,
            I => \N__26218\
        );

    \I__5905\ : CascadeMux
    port map (
            O => \N__26229\,
            I => \N__26215\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__26228\,
            I => \N__26212\
        );

    \I__5903\ : CascadeMux
    port map (
            O => \N__26227\,
            I => \N__26209\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__26224\,
            I => \N__26204\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__26221\,
            I => \N__26201\
        );

    \I__5900\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26198\
        );

    \I__5899\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26195\
        );

    \I__5898\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26192\
        );

    \I__5897\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26189\
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__26208\,
            I => \N__26186\
        );

    \I__5895\ : CascadeMux
    port map (
            O => \N__26207\,
            I => \N__26183\
        );

    \I__5894\ : Span4Mux_v
    port map (
            O => \N__26204\,
            I => \N__26172\
        );

    \I__5893\ : Span4Mux_h
    port map (
            O => \N__26201\,
            I => \N__26172\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__26198\,
            I => \N__26172\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__26195\,
            I => \N__26169\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__26192\,
            I => \N__26166\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__26189\,
            I => \N__26163\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26160\
        );

    \I__5887\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26157\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__26182\,
            I => \N__26154\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__26181\,
            I => \N__26151\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__26180\,
            I => \N__26147\
        );

    \I__5883\ : CascadeMux
    port map (
            O => \N__26179\,
            I => \N__26144\
        );

    \I__5882\ : Span4Mux_v
    port map (
            O => \N__26172\,
            I => \N__26134\
        );

    \I__5881\ : Span4Mux_v
    port map (
            O => \N__26169\,
            I => \N__26134\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__26166\,
            I => \N__26134\
        );

    \I__5879\ : Span4Mux_s1_v
    port map (
            O => \N__26163\,
            I => \N__26129\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__26160\,
            I => \N__26129\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26126\
        );

    \I__5876\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26123\
        );

    \I__5875\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26120\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__26150\,
            I => \N__26117\
        );

    \I__5873\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26114\
        );

    \I__5872\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26111\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__26143\,
            I => \N__26108\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__26142\,
            I => \N__26105\
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__26141\,
            I => \N__26102\
        );

    \I__5868\ : Span4Mux_h
    port map (
            O => \N__26134\,
            I => \N__26099\
        );

    \I__5867\ : Span4Mux_v
    port map (
            O => \N__26129\,
            I => \N__26092\
        );

    \I__5866\ : Span4Mux_h
    port map (
            O => \N__26126\,
            I => \N__26092\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__26123\,
            I => \N__26092\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__26120\,
            I => \N__26089\
        );

    \I__5863\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26086\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__26114\,
            I => \N__26081\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26081\
        );

    \I__5860\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26078\
        );

    \I__5859\ : InMux
    port map (
            O => \N__26105\,
            I => \N__26075\
        );

    \I__5858\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26072\
        );

    \I__5857\ : Span4Mux_h
    port map (
            O => \N__26099\,
            I => \N__26069\
        );

    \I__5856\ : Span4Mux_v
    port map (
            O => \N__26092\,
            I => \N__26062\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__26089\,
            I => \N__26062\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__26086\,
            I => \N__26062\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__26081\,
            I => \N__26055\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__26078\,
            I => \N__26055\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__26075\,
            I => \N__26055\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__26072\,
            I => \N__26052\
        );

    \I__5849\ : Span4Mux_h
    port map (
            O => \N__26069\,
            I => \N__26041\
        );

    \I__5848\ : Span4Mux_v
    port map (
            O => \N__26062\,
            I => \N__26041\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__26055\,
            I => \N__26041\
        );

    \I__5846\ : Span4Mux_h
    port map (
            O => \N__26052\,
            I => \N__26041\
        );

    \I__5845\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26038\
        );

    \I__5844\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26035\
        );

    \I__5843\ : Odrv4
    port map (
            O => \N__26041\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__26038\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__26035\,
            I => \M_this_sprites_address_qZ0Z_9\
        );

    \I__5840\ : InMux
    port map (
            O => \N__26028\,
            I => \N__26025\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__26025\,
            I => \M_this_sprites_address_q_RNO_0Z0Z_3\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__26022\,
            I => \N__26015\
        );

    \I__5837\ : CascadeMux
    port map (
            O => \N__26021\,
            I => \N__26012\
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__26020\,
            I => \N__26009\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__26019\,
            I => \N__26001\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__26018\,
            I => \N__25997\
        );

    \I__5833\ : InMux
    port map (
            O => \N__26015\,
            I => \N__25994\
        );

    \I__5832\ : InMux
    port map (
            O => \N__26012\,
            I => \N__25991\
        );

    \I__5831\ : InMux
    port map (
            O => \N__26009\,
            I => \N__25988\
        );

    \I__5830\ : CascadeMux
    port map (
            O => \N__26008\,
            I => \N__25985\
        );

    \I__5829\ : CascadeMux
    port map (
            O => \N__26007\,
            I => \N__25978\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__26006\,
            I => \N__25974\
        );

    \I__5827\ : CascadeMux
    port map (
            O => \N__26005\,
            I => \N__25971\
        );

    \I__5826\ : CascadeMux
    port map (
            O => \N__26004\,
            I => \N__25968\
        );

    \I__5825\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25965\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__26000\,
            I => \N__25962\
        );

    \I__5823\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25959\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__25994\,
            I => \N__25956\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25953\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25950\
        );

    \I__5819\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25947\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__25984\,
            I => \N__25944\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__25983\,
            I => \N__25941\
        );

    \I__5816\ : CascadeMux
    port map (
            O => \N__25982\,
            I => \N__25938\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__25981\,
            I => \N__25935\
        );

    \I__5814\ : InMux
    port map (
            O => \N__25978\,
            I => \N__25932\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__25977\,
            I => \N__25929\
        );

    \I__5812\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25926\
        );

    \I__5811\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25923\
        );

    \I__5810\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25920\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__25965\,
            I => \N__25917\
        );

    \I__5808\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25914\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__25959\,
            I => \N__25911\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__25956\,
            I => \N__25902\
        );

    \I__5805\ : Span4Mux_v
    port map (
            O => \N__25953\,
            I => \N__25902\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__25950\,
            I => \N__25902\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25902\
        );

    \I__5802\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25899\
        );

    \I__5801\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25896\
        );

    \I__5800\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25893\
        );

    \I__5799\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25890\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__25932\,
            I => \N__25887\
        );

    \I__5797\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25884\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__25926\,
            I => \N__25881\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__25923\,
            I => \N__25878\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__25920\,
            I => \N__25875\
        );

    \I__5793\ : Span4Mux_h
    port map (
            O => \N__25917\,
            I => \N__25871\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__25914\,
            I => \N__25868\
        );

    \I__5791\ : Span4Mux_h
    port map (
            O => \N__25911\,
            I => \N__25863\
        );

    \I__5790\ : Span4Mux_v
    port map (
            O => \N__25902\,
            I => \N__25863\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__25899\,
            I => \N__25858\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__25896\,
            I => \N__25858\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__25893\,
            I => \N__25851\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__25890\,
            I => \N__25851\
        );

    \I__5785\ : Span4Mux_v
    port map (
            O => \N__25887\,
            I => \N__25851\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__25884\,
            I => \N__25848\
        );

    \I__5783\ : Sp12to4
    port map (
            O => \N__25881\,
            I => \N__25845\
        );

    \I__5782\ : Span4Mux_h
    port map (
            O => \N__25878\,
            I => \N__25840\
        );

    \I__5781\ : Span4Mux_h
    port map (
            O => \N__25875\,
            I => \N__25840\
        );

    \I__5780\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25837\
        );

    \I__5779\ : Sp12to4
    port map (
            O => \N__25871\,
            I => \N__25832\
        );

    \I__5778\ : Span12Mux_s8_h
    port map (
            O => \N__25868\,
            I => \N__25832\
        );

    \I__5777\ : Span4Mux_h
    port map (
            O => \N__25863\,
            I => \N__25829\
        );

    \I__5776\ : Span4Mux_v
    port map (
            O => \N__25858\,
            I => \N__25823\
        );

    \I__5775\ : Span4Mux_v
    port map (
            O => \N__25851\,
            I => \N__25823\
        );

    \I__5774\ : Span12Mux_s10_h
    port map (
            O => \N__25848\,
            I => \N__25816\
        );

    \I__5773\ : Span12Mux_s10_h
    port map (
            O => \N__25845\,
            I => \N__25816\
        );

    \I__5772\ : Sp12to4
    port map (
            O => \N__25840\,
            I => \N__25816\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__25837\,
            I => \N__25813\
        );

    \I__5770\ : Span12Mux_v
    port map (
            O => \N__25832\,
            I => \N__25808\
        );

    \I__5769\ : Sp12to4
    port map (
            O => \N__25829\,
            I => \N__25808\
        );

    \I__5768\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25805\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__25823\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5766\ : Odrv12
    port map (
            O => \N__25816\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5765\ : Odrv4
    port map (
            O => \N__25813\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5764\ : Odrv12
    port map (
            O => \N__25808\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__25805\,
            I => \M_this_sprites_address_qZ0Z_3\
        );

    \I__5762\ : CascadeMux
    port map (
            O => \N__25794\,
            I => \N__25791\
        );

    \I__5761\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25788\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__25788\,
            I => \N_50\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__25785\,
            I => \N__25780\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__25784\,
            I => \N__25777\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__25783\,
            I => \N__25773\
        );

    \I__5756\ : InMux
    port map (
            O => \N__25780\,
            I => \N__25768\
        );

    \I__5755\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25765\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__25776\,
            I => \N__25762\
        );

    \I__5753\ : InMux
    port map (
            O => \N__25773\,
            I => \N__25758\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__25772\,
            I => \N__25755\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__25771\,
            I => \N__25752\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25746\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__25765\,
            I => \N__25746\
        );

    \I__5748\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25743\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__25761\,
            I => \N__25740\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25736\
        );

    \I__5745\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25733\
        );

    \I__5744\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25730\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__25751\,
            I => \N__25727\
        );

    \I__5742\ : Span4Mux_s2_v
    port map (
            O => \N__25746\,
            I => \N__25720\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__25743\,
            I => \N__25720\
        );

    \I__5740\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25717\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__25739\,
            I => \N__25714\
        );

    \I__5738\ : Span4Mux_h
    port map (
            O => \N__25736\,
            I => \N__25708\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__25733\,
            I => \N__25708\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__25730\,
            I => \N__25705\
        );

    \I__5735\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25702\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__25726\,
            I => \N__25698\
        );

    \I__5733\ : CascadeMux
    port map (
            O => \N__25725\,
            I => \N__25695\
        );

    \I__5732\ : Span4Mux_v
    port map (
            O => \N__25720\,
            I => \N__25689\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__25717\,
            I => \N__25689\
        );

    \I__5730\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25686\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__25713\,
            I => \N__25683\
        );

    \I__5728\ : Span4Mux_v
    port map (
            O => \N__25708\,
            I => \N__25675\
        );

    \I__5727\ : Span4Mux_h
    port map (
            O => \N__25705\,
            I => \N__25675\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__25702\,
            I => \N__25675\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__25701\,
            I => \N__25672\
        );

    \I__5724\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25669\
        );

    \I__5723\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25666\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__25694\,
            I => \N__25663\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__25689\,
            I => \N__25658\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25658\
        );

    \I__5719\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25655\
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__25682\,
            I => \N__25652\
        );

    \I__5717\ : Span4Mux_v
    port map (
            O => \N__25675\,
            I => \N__25648\
        );

    \I__5716\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25645\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25642\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__25666\,
            I => \N__25639\
        );

    \I__5713\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25636\
        );

    \I__5712\ : Span4Mux_v
    port map (
            O => \N__25658\,
            I => \N__25631\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__25655\,
            I => \N__25631\
        );

    \I__5710\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25628\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__25651\,
            I => \N__25625\
        );

    \I__5708\ : Sp12to4
    port map (
            O => \N__25648\,
            I => \N__25620\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__25645\,
            I => \N__25620\
        );

    \I__5706\ : Span4Mux_v
    port map (
            O => \N__25642\,
            I => \N__25613\
        );

    \I__5705\ : Span4Mux_h
    port map (
            O => \N__25639\,
            I => \N__25613\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25613\
        );

    \I__5703\ : Span4Mux_h
    port map (
            O => \N__25631\,
            I => \N__25608\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__25628\,
            I => \N__25608\
        );

    \I__5701\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25605\
        );

    \I__5700\ : Span12Mux_h
    port map (
            O => \N__25620\,
            I => \N__25602\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__25613\,
            I => \N__25595\
        );

    \I__5698\ : Span4Mux_v
    port map (
            O => \N__25608\,
            I => \N__25595\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__25605\,
            I => \N__25595\
        );

    \I__5696\ : Odrv12
    port map (
            O => \N__25602\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__25595\,
            I => \M_this_ppu_sprites_addr_3\
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__25590\,
            I => \N__25585\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__25589\,
            I => \N__25581\
        );

    \I__5692\ : CascadeMux
    port map (
            O => \N__25588\,
            I => \N__25578\
        );

    \I__5691\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25573\
        );

    \I__5690\ : CascadeMux
    port map (
            O => \N__25584\,
            I => \N__25570\
        );

    \I__5689\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25566\
        );

    \I__5688\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25563\
        );

    \I__5687\ : CascadeMux
    port map (
            O => \N__25577\,
            I => \N__25560\
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__25576\,
            I => \N__25557\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__25573\,
            I => \N__25554\
        );

    \I__5684\ : InMux
    port map (
            O => \N__25570\,
            I => \N__25551\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__25569\,
            I => \N__25548\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__25566\,
            I => \N__25541\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__25563\,
            I => \N__25538\
        );

    \I__5680\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25535\
        );

    \I__5679\ : InMux
    port map (
            O => \N__25557\,
            I => \N__25532\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__25554\,
            I => \N__25526\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__25551\,
            I => \N__25526\
        );

    \I__5676\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25523\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__25547\,
            I => \N__25520\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__25546\,
            I => \N__25516\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__25545\,
            I => \N__25513\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__25544\,
            I => \N__25508\
        );

    \I__5671\ : Span4Mux_v
    port map (
            O => \N__25541\,
            I => \N__25501\
        );

    \I__5670\ : Span4Mux_h
    port map (
            O => \N__25538\,
            I => \N__25501\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__25535\,
            I => \N__25501\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__25532\,
            I => \N__25498\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__25531\,
            I => \N__25495\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__25526\,
            I => \N__25490\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__25523\,
            I => \N__25490\
        );

    \I__5664\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25487\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__25519\,
            I => \N__25484\
        );

    \I__5662\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25481\
        );

    \I__5661\ : InMux
    port map (
            O => \N__25513\,
            I => \N__25478\
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__25512\,
            I => \N__25475\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__25511\,
            I => \N__25472\
        );

    \I__5658\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25468\
        );

    \I__5657\ : Span4Mux_v
    port map (
            O => \N__25501\,
            I => \N__25463\
        );

    \I__5656\ : Span4Mux_v
    port map (
            O => \N__25498\,
            I => \N__25463\
        );

    \I__5655\ : InMux
    port map (
            O => \N__25495\,
            I => \N__25460\
        );

    \I__5654\ : Span4Mux_v
    port map (
            O => \N__25490\,
            I => \N__25455\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25455\
        );

    \I__5652\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25452\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__25481\,
            I => \N__25449\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__25478\,
            I => \N__25446\
        );

    \I__5649\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25443\
        );

    \I__5648\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25440\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__25471\,
            I => \N__25437\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__25468\,
            I => \N__25434\
        );

    \I__5645\ : Sp12to4
    port map (
            O => \N__25463\,
            I => \N__25429\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__25460\,
            I => \N__25429\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__25455\,
            I => \N__25424\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__25452\,
            I => \N__25424\
        );

    \I__5641\ : Span4Mux_v
    port map (
            O => \N__25449\,
            I => \N__25415\
        );

    \I__5640\ : Span4Mux_v
    port map (
            O => \N__25446\,
            I => \N__25415\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25415\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__25440\,
            I => \N__25415\
        );

    \I__5637\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25412\
        );

    \I__5636\ : Span12Mux_s10_h
    port map (
            O => \N__25434\,
            I => \N__25407\
        );

    \I__5635\ : Span12Mux_h
    port map (
            O => \N__25429\,
            I => \N__25404\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__25424\,
            I => \N__25397\
        );

    \I__5633\ : Span4Mux_v
    port map (
            O => \N__25415\,
            I => \N__25397\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25397\
        );

    \I__5631\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25394\
        );

    \I__5630\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25391\
        );

    \I__5629\ : Odrv12
    port map (
            O => \N__25407\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5628\ : Odrv12
    port map (
            O => \N__25404\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__25397\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__25394\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__25391\,
            I => \M_this_sprites_address_qZ0Z_2\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__25380\,
            I => \N__25377\
        );

    \I__5623\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__25374\,
            I => \N_103\
        );

    \I__5621\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25367\
        );

    \I__5620\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25363\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__25367\,
            I => \N__25359\
        );

    \I__5618\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25356\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__25363\,
            I => \N__25353\
        );

    \I__5616\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25350\
        );

    \I__5615\ : Span4Mux_v
    port map (
            O => \N__25359\,
            I => \N__25343\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__25356\,
            I => \N__25343\
        );

    \I__5613\ : Span4Mux_s3_v
    port map (
            O => \N__25353\,
            I => \N__25337\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__25350\,
            I => \N__25337\
        );

    \I__5611\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25334\
        );

    \I__5610\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25331\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__25343\,
            I => \N__25327\
        );

    \I__5608\ : InMux
    port map (
            O => \N__25342\,
            I => \N__25324\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__25337\,
            I => \N__25317\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__25334\,
            I => \N__25317\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__25331\,
            I => \N__25317\
        );

    \I__5604\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25314\
        );

    \I__5603\ : Sp12to4
    port map (
            O => \N__25327\,
            I => \N__25311\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__25324\,
            I => \N__25308\
        );

    \I__5601\ : Span4Mux_v
    port map (
            O => \N__25317\,
            I => \N__25303\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25303\
        );

    \I__5599\ : Span12Mux_h
    port map (
            O => \N__25311\,
            I => \N__25300\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__25308\,
            I => \N__25295\
        );

    \I__5597\ : Span4Mux_v
    port map (
            O => \N__25303\,
            I => \N__25295\
        );

    \I__5596\ : Odrv12
    port map (
            O => \N__25300\,
            I => \M_this_sprites_ram_write_data_iv_i_i_1\
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__25295\,
            I => \M_this_sprites_ram_write_data_iv_i_i_1\
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__25290\,
            I => \N__25287\
        );

    \I__5593\ : InMux
    port map (
            O => \N__25287\,
            I => \N__25284\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__25284\,
            I => \N__25281\
        );

    \I__5591\ : Odrv4
    port map (
            O => \N__25281\,
            I => \M_this_data_tmp_qZ0Z_2\
        );

    \I__5590\ : InMux
    port map (
            O => \N__25278\,
            I => \N__25275\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__25275\,
            I => \N__25272\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__25269\,
            I => \N__25266\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__25266\,
            I => \N_746_0\
        );

    \I__5585\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25260\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__25260\,
            I => \N__25257\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__25257\,
            I => \N__25254\
        );

    \I__5582\ : Odrv4
    port map (
            O => \N__25254\,
            I => \M_this_oam_ram_write_data_28\
        );

    \I__5581\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__25248\,
            I => \N__25241\
        );

    \I__5579\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25238\
        );

    \I__5578\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25235\
        );

    \I__5577\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25229\
        );

    \I__5576\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25226\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__25241\,
            I => \N__25222\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__25238\,
            I => \N__25217\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__25235\,
            I => \N__25217\
        );

    \I__5572\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25210\
        );

    \I__5571\ : InMux
    port map (
            O => \N__25233\,
            I => \N__25210\
        );

    \I__5570\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25210\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__25229\,
            I => \N__25205\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__25226\,
            I => \N__25205\
        );

    \I__5567\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25202\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__25222\,
            I => \N__25199\
        );

    \I__5565\ : Span4Mux_v
    port map (
            O => \N__25217\,
            I => \N__25194\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__25210\,
            I => \N__25194\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__25205\,
            I => \N__25191\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__25202\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__25199\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__25194\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__25191\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__5558\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__25179\,
            I => \un1_M_this_sprites_address_q_cry_0_THRU_CO\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__25176\,
            I => \N__25173\
        );

    \I__5555\ : InMux
    port map (
            O => \N__25173\,
            I => \N__25165\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__25172\,
            I => \N__25162\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__25171\,
            I => \N__25159\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__25170\,
            I => \N__25152\
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__25169\,
            I => \N__25149\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__25168\,
            I => \N__25146\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__25165\,
            I => \N__25143\
        );

    \I__5548\ : InMux
    port map (
            O => \N__25162\,
            I => \N__25140\
        );

    \I__5547\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25137\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__25158\,
            I => \N__25134\
        );

    \I__5545\ : CascadeMux
    port map (
            O => \N__25157\,
            I => \N__25131\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__25156\,
            I => \N__25124\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__25155\,
            I => \N__25121\
        );

    \I__5542\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25118\
        );

    \I__5541\ : InMux
    port map (
            O => \N__25149\,
            I => \N__25115\
        );

    \I__5540\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25110\
        );

    \I__5539\ : Span4Mux_h
    port map (
            O => \N__25143\,
            I => \N__25103\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__25140\,
            I => \N__25103\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__25137\,
            I => \N__25103\
        );

    \I__5536\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25100\
        );

    \I__5535\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25097\
        );

    \I__5534\ : CascadeMux
    port map (
            O => \N__25130\,
            I => \N__25094\
        );

    \I__5533\ : CascadeMux
    port map (
            O => \N__25129\,
            I => \N__25091\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__25128\,
            I => \N__25088\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__25127\,
            I => \N__25085\
        );

    \I__5530\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25082\
        );

    \I__5529\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25079\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__25118\,
            I => \N__25076\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25073\
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__25114\,
            I => \N__25070\
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__25113\,
            I => \N__25067\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__25110\,
            I => \N__25064\
        );

    \I__5523\ : Span4Mux_v
    port map (
            O => \N__25103\,
            I => \N__25059\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25059\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__25097\,
            I => \N__25056\
        );

    \I__5520\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25053\
        );

    \I__5519\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25050\
        );

    \I__5518\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25047\
        );

    \I__5517\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25044\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__25082\,
            I => \N__25041\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25038\
        );

    \I__5514\ : Span4Mux_h
    port map (
            O => \N__25076\,
            I => \N__25033\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__25073\,
            I => \N__25033\
        );

    \I__5512\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25030\
        );

    \I__5511\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25027\
        );

    \I__5510\ : Span4Mux_h
    port map (
            O => \N__25064\,
            I => \N__25022\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__25059\,
            I => \N__25022\
        );

    \I__5508\ : Span4Mux_v
    port map (
            O => \N__25056\,
            I => \N__25019\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__25053\,
            I => \N__25013\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__25050\,
            I => \N__25013\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__25047\,
            I => \N__25008\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__25044\,
            I => \N__25008\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__25041\,
            I => \N__25005\
        );

    \I__5502\ : Span4Mux_h
    port map (
            O => \N__25038\,
            I => \N__25002\
        );

    \I__5501\ : Sp12to4
    port map (
            O => \N__25033\,
            I => \N__24998\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__24995\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__25027\,
            I => \N__24992\
        );

    \I__5498\ : Sp12to4
    port map (
            O => \N__25022\,
            I => \N__24989\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__25019\,
            I => \N__24986\
        );

    \I__5496\ : InMux
    port map (
            O => \N__25018\,
            I => \N__24983\
        );

    \I__5495\ : Span4Mux_v
    port map (
            O => \N__25013\,
            I => \N__24978\
        );

    \I__5494\ : Span4Mux_v
    port map (
            O => \N__25008\,
            I => \N__24978\
        );

    \I__5493\ : Span4Mux_v
    port map (
            O => \N__25005\,
            I => \N__24973\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__25002\,
            I => \N__24973\
        );

    \I__5491\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24970\
        );

    \I__5490\ : Span12Mux_v
    port map (
            O => \N__24998\,
            I => \N__24967\
        );

    \I__5489\ : Span12Mux_s11_h
    port map (
            O => \N__24995\,
            I => \N__24960\
        );

    \I__5488\ : Span12Mux_s11_h
    port map (
            O => \N__24992\,
            I => \N__24960\
        );

    \I__5487\ : Span12Mux_h
    port map (
            O => \N__24989\,
            I => \N__24960\
        );

    \I__5486\ : Span4Mux_v
    port map (
            O => \N__24986\,
            I => \N__24955\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__24983\,
            I => \N__24955\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__24978\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5483\ : Odrv4
    port map (
            O => \N__24973\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__24970\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5481\ : Odrv12
    port map (
            O => \N__24967\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5480\ : Odrv12
    port map (
            O => \N__24960\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__24955\,
            I => \M_this_sprites_address_qZ0Z_7\
        );

    \I__5478\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24939\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__24939\,
            I => \M_this_sprites_address_qc_9_0\
        );

    \I__5476\ : CascadeMux
    port map (
            O => \N__24936\,
            I => \N__24933\
        );

    \I__5475\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24930\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__24930\,
            I => \N__24927\
        );

    \I__5473\ : Odrv12
    port map (
            O => \N__24927\,
            I => \M_this_oam_ram_read_data_i_19\
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__24924\,
            I => \N__24921\
        );

    \I__5471\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24918\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__24918\,
            I => \N__24915\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__24915\,
            I => \M_this_oam_ram_read_data_i_11\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__5467\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24905\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__24908\,
            I => \N__24902\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__24905\,
            I => \N__24899\
        );

    \I__5464\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24896\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__24899\,
            I => \N__24891\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__24896\,
            I => \N__24891\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__24891\,
            I => \N__24888\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__24888\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__5459\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24882\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__24882\,
            I => \N__24879\
        );

    \I__5457\ : Odrv4
    port map (
            O => \N__24879\,
            I => \this_ppu.un1_M_haddress_q_2_7\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__24876\,
            I => \N__24873\
        );

    \I__5455\ : CascadeBuf
    port map (
            O => \N__24873\,
            I => \N__24870\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__24870\,
            I => \N__24867\
        );

    \I__5453\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__5451\ : Span4Mux_h
    port map (
            O => \N__24861\,
            I => \N__24857\
        );

    \I__5450\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24854\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__24857\,
            I => \N__24850\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__24854\,
            I => \N__24847\
        );

    \I__5447\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24844\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__24850\,
            I => \N__24841\
        );

    \I__5445\ : Odrv12
    port map (
            O => \N__24847\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__24844\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__24841\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__5442\ : InMux
    port map (
            O => \N__24834\,
            I => \N__24830\
        );

    \I__5441\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24827\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__24830\,
            I => \un1_M_this_oam_address_q_c4\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__24827\,
            I => \un1_M_this_oam_address_q_c4\
        );

    \I__5438\ : CascadeMux
    port map (
            O => \N__24822\,
            I => \N__24819\
        );

    \I__5437\ : CascadeBuf
    port map (
            O => \N__24819\,
            I => \N__24816\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__24816\,
            I => \N__24813\
        );

    \I__5435\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24810\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__24810\,
            I => \N__24806\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__24809\,
            I => \N__24803\
        );

    \I__5432\ : Span4Mux_v
    port map (
            O => \N__24806\,
            I => \N__24800\
        );

    \I__5431\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24797\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__24800\,
            I => \N__24794\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__24797\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__5428\ : Odrv4
    port map (
            O => \N__24794\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__5426\ : CascadeBuf
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__5425\ : CascadeMux
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__5424\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24776\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__24779\,
            I => \N__24773\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__24776\,
            I => \N__24769\
        );

    \I__5421\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24766\
        );

    \I__5420\ : InMux
    port map (
            O => \N__24772\,
            I => \N__24763\
        );

    \I__5419\ : Span12Mux_s11_v
    port map (
            O => \N__24769\,
            I => \N__24760\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__24766\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__24763\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5416\ : Odrv12
    port map (
            O => \N__24760\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__5415\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__24750\,
            I => \M_this_sprites_address_qc_2_1\
        );

    \I__5413\ : InMux
    port map (
            O => \N__24747\,
            I => \un1_M_this_sprites_address_q_cry_12\
        );

    \I__5412\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24741\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__24741\,
            I => \M_this_sprites_address_q_RNO_0Z0Z_12\
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__24738\,
            I => \N_807_cascade_\
        );

    \I__5409\ : InMux
    port map (
            O => \N__24735\,
            I => \N__24732\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__24732\,
            I => \N__24729\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__24729\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_7\
        );

    \I__5406\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__24723\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_8\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__24720\,
            I => \N_803_cascade_\
        );

    \I__5403\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__24714\,
            I => \M_this_sprites_address_qc_10_0\
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__5400\ : InMux
    port map (
            O => \N__24708\,
            I => \N__24702\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__24707\,
            I => \N__24699\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__24706\,
            I => \N__24695\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__24705\,
            I => \N__24692\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__24702\,
            I => \N__24686\
        );

    \I__5395\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24683\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__24698\,
            I => \N__24680\
        );

    \I__5393\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24674\
        );

    \I__5392\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24671\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__24691\,
            I => \N__24668\
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__24690\,
            I => \N__24665\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__24689\,
            I => \N__24662\
        );

    \I__5388\ : Span4Mux_s3_v
    port map (
            O => \N__24686\,
            I => \N__24657\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__24683\,
            I => \N__24657\
        );

    \I__5386\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24654\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__24679\,
            I => \N__24651\
        );

    \I__5384\ : CascadeMux
    port map (
            O => \N__24678\,
            I => \N__24647\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__24677\,
            I => \N__24644\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__24674\,
            I => \N__24637\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24637\
        );

    \I__5380\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24634\
        );

    \I__5379\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24631\
        );

    \I__5378\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24628\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__24657\,
            I => \N__24623\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__24654\,
            I => \N__24623\
        );

    \I__5375\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24620\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__24650\,
            I => \N__24617\
        );

    \I__5373\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24613\
        );

    \I__5372\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24610\
        );

    \I__5371\ : CascadeMux
    port map (
            O => \N__24643\,
            I => \N__24607\
        );

    \I__5370\ : CascadeMux
    port map (
            O => \N__24642\,
            I => \N__24604\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__24637\,
            I => \N__24596\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__24634\,
            I => \N__24596\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__24631\,
            I => \N__24596\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24593\
        );

    \I__5365\ : Span4Mux_v
    port map (
            O => \N__24623\,
            I => \N__24588\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__24620\,
            I => \N__24588\
        );

    \I__5363\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24585\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__24616\,
            I => \N__24582\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__24613\,
            I => \N__24579\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__24610\,
            I => \N__24576\
        );

    \I__5359\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24573\
        );

    \I__5358\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24570\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__24603\,
            I => \N__24567\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__24596\,
            I => \N__24562\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__24593\,
            I => \N__24562\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__24588\,
            I => \N__24557\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24557\
        );

    \I__5352\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24554\
        );

    \I__5351\ : Span4Mux_v
    port map (
            O => \N__24579\,
            I => \N__24547\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__24576\,
            I => \N__24547\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__24573\,
            I => \N__24547\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24544\
        );

    \I__5347\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24541\
        );

    \I__5346\ : Sp12to4
    port map (
            O => \N__24562\,
            I => \N__24538\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__24557\,
            I => \N__24533\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__24554\,
            I => \N__24533\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__24547\,
            I => \N__24526\
        );

    \I__5342\ : Span4Mux_v
    port map (
            O => \N__24544\,
            I => \N__24526\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__24541\,
            I => \N__24526\
        );

    \I__5340\ : Span12Mux_h
    port map (
            O => \N__24538\,
            I => \N__24521\
        );

    \I__5339\ : Span4Mux_h
    port map (
            O => \N__24533\,
            I => \N__24516\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__24526\,
            I => \N__24516\
        );

    \I__5337\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24513\
        );

    \I__5336\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24510\
        );

    \I__5335\ : Odrv12
    port map (
            O => \N__24521\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__24516\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__24513\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__24510\,
            I => \M_this_sprites_address_qZ0Z_8\
        );

    \I__5331\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24498\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__24498\,
            I => \N_602\
        );

    \I__5329\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24491\
        );

    \I__5328\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24486\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24480\
        );

    \I__5326\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24477\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__24489\,
            I => \N__24473\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__24486\,
            I => \N__24470\
        );

    \I__5323\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24465\
        );

    \I__5322\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24465\
        );

    \I__5321\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24462\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__24480\,
            I => \N__24457\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__24477\,
            I => \N__24457\
        );

    \I__5318\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24454\
        );

    \I__5317\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24451\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__24470\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__24465\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__24462\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5313\ : Odrv4
    port map (
            O => \N__24457\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__24454\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__24451\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__5310\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24434\
        );

    \I__5309\ : CascadeMux
    port map (
            O => \N__24437\,
            I => \N__24429\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__24434\,
            I => \N__24426\
        );

    \I__5307\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24423\
        );

    \I__5306\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24418\
        );

    \I__5305\ : InMux
    port map (
            O => \N__24429\,
            I => \N__24415\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__24426\,
            I => \N__24412\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__24423\,
            I => \N__24409\
        );

    \I__5302\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24404\
        );

    \I__5301\ : InMux
    port map (
            O => \N__24421\,
            I => \N__24404\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__24418\,
            I => \N__24399\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__24415\,
            I => \N__24399\
        );

    \I__5298\ : Span4Mux_h
    port map (
            O => \N__24412\,
            I => \N__24396\
        );

    \I__5297\ : Span4Mux_v
    port map (
            O => \N__24409\,
            I => \N__24393\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__24404\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5295\ : Odrv12
    port map (
            O => \N__24399\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__24396\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__24393\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__5292\ : InMux
    port map (
            O => \N__24384\,
            I => \un1_M_this_sprites_address_q_cry_3\
        );

    \I__5291\ : InMux
    port map (
            O => \N__24381\,
            I => \un1_M_this_sprites_address_q_cry_4\
        );

    \I__5290\ : InMux
    port map (
            O => \N__24378\,
            I => \un1_M_this_sprites_address_q_cry_5\
        );

    \I__5289\ : InMux
    port map (
            O => \N__24375\,
            I => \un1_M_this_sprites_address_q_cry_6\
        );

    \I__5288\ : InMux
    port map (
            O => \N__24372\,
            I => \bfn_21_14_0_\
        );

    \I__5287\ : InMux
    port map (
            O => \N__24369\,
            I => \un1_M_this_sprites_address_q_cry_8\
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__24366\,
            I => \N__24361\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__24365\,
            I => \N__24358\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__24364\,
            I => \N__24353\
        );

    \I__5283\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24350\
        );

    \I__5282\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24347\
        );

    \I__5281\ : CascadeMux
    port map (
            O => \N__24357\,
            I => \N__24344\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__24356\,
            I => \N__24340\
        );

    \I__5279\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24334\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__24350\,
            I => \N__24329\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__24347\,
            I => \N__24326\
        );

    \I__5276\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24323\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__24343\,
            I => \N__24320\
        );

    \I__5274\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24316\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__24339\,
            I => \N__24313\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__24338\,
            I => \N__24310\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__24337\,
            I => \N__24307\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__24334\,
            I => \N__24304\
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__24333\,
            I => \N__24301\
        );

    \I__5268\ : CascadeMux
    port map (
            O => \N__24332\,
            I => \N__24298\
        );

    \I__5267\ : Span4Mux_s3_v
    port map (
            O => \N__24329\,
            I => \N__24290\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__24326\,
            I => \N__24290\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__24323\,
            I => \N__24290\
        );

    \I__5264\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24287\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__24319\,
            I => \N__24284\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__24316\,
            I => \N__24280\
        );

    \I__5261\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24277\
        );

    \I__5260\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24274\
        );

    \I__5259\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24271\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__24304\,
            I => \N__24267\
        );

    \I__5257\ : InMux
    port map (
            O => \N__24301\,
            I => \N__24264\
        );

    \I__5256\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24261\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__24297\,
            I => \N__24258\
        );

    \I__5254\ : Span4Mux_v
    port map (
            O => \N__24290\,
            I => \N__24253\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__24287\,
            I => \N__24253\
        );

    \I__5252\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24250\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__24283\,
            I => \N__24247\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__24280\,
            I => \N__24242\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__24277\,
            I => \N__24242\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__24274\,
            I => \N__24237\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__24271\,
            I => \N__24237\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__24270\,
            I => \N__24234\
        );

    \I__5245\ : Span4Mux_h
    port map (
            O => \N__24267\,
            I => \N__24227\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__24264\,
            I => \N__24227\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__24261\,
            I => \N__24227\
        );

    \I__5242\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24224\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__24253\,
            I => \N__24219\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__24250\,
            I => \N__24219\
        );

    \I__5239\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24216\
        );

    \I__5238\ : Span4Mux_v
    port map (
            O => \N__24242\,
            I => \N__24210\
        );

    \I__5237\ : Span4Mux_v
    port map (
            O => \N__24237\,
            I => \N__24210\
        );

    \I__5236\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24207\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__24227\,
            I => \N__24198\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__24224\,
            I => \N__24198\
        );

    \I__5233\ : Span4Mux_v
    port map (
            O => \N__24219\,
            I => \N__24198\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__24216\,
            I => \N__24198\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__24215\,
            I => \N__24195\
        );

    \I__5230\ : Span4Mux_h
    port map (
            O => \N__24210\,
            I => \N__24191\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__24207\,
            I => \N__24188\
        );

    \I__5228\ : Span4Mux_v
    port map (
            O => \N__24198\,
            I => \N__24185\
        );

    \I__5227\ : InMux
    port map (
            O => \N__24195\,
            I => \N__24182\
        );

    \I__5226\ : InMux
    port map (
            O => \N__24194\,
            I => \N__24178\
        );

    \I__5225\ : Sp12to4
    port map (
            O => \N__24191\,
            I => \N__24173\
        );

    \I__5224\ : Span12Mux_s11_h
    port map (
            O => \N__24188\,
            I => \N__24173\
        );

    \I__5223\ : Sp12to4
    port map (
            O => \N__24185\,
            I => \N__24168\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__24182\,
            I => \N__24168\
        );

    \I__5221\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24165\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__24178\,
            I => \N__24162\
        );

    \I__5219\ : Odrv12
    port map (
            O => \N__24173\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5218\ : Odrv12
    port map (
            O => \N__24168\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__24165\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__24162\,
            I => \M_this_sprites_address_qZ0Z_10\
        );

    \I__5215\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24150\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__24150\,
            I => \N__24147\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__24147\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_10\
        );

    \I__5212\ : InMux
    port map (
            O => \N__24144\,
            I => \un1_M_this_sprites_address_q_cry_9\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24141\,
            I => \N__24138\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__24138\,
            I => \N__24135\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__24135\,
            I => \M_this_sprites_address_q_RNO_1Z0Z_11\
        );

    \I__5208\ : InMux
    port map (
            O => \N__24132\,
            I => \un1_M_this_sprites_address_q_cry_10\
        );

    \I__5207\ : InMux
    port map (
            O => \N__24129\,
            I => \un1_M_this_sprites_address_q_cry_11\
        );

    \I__5206\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24123\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__24123\,
            I => \N__24120\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__24120\,
            I => \N__24117\
        );

    \I__5203\ : Span4Mux_v
    port map (
            O => \N__24117\,
            I => \N__24114\
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__24114\,
            I => \this_sprites_ram.mem_out_bus6_1\
        );

    \I__5201\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24108\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24105\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__24105\,
            I => \N__24102\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__24102\,
            I => \this_sprites_ram.mem_out_bus2_1\
        );

    \I__5197\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24096\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__24096\,
            I => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\
        );

    \I__5195\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24090\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__24090\,
            I => \N__24087\
        );

    \I__5193\ : Span4Mux_v
    port map (
            O => \N__24087\,
            I => \N__24084\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__24084\,
            I => \this_sprites_ram.mem_out_bus5_2\
        );

    \I__5191\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24075\
        );

    \I__5189\ : Span4Mux_h
    port map (
            O => \N__24075\,
            I => \N__24072\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__24072\,
            I => \this_sprites_ram.mem_out_bus1_2\
        );

    \I__5187\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24066\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__24066\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__24063\,
            I => \N__24060\
        );

    \I__5184\ : InMux
    port map (
            O => \N__24060\,
            I => \N__24057\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24054\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__24054\,
            I => \N__24051\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__24051\,
            I => \this_sprites_ram.mem_out_bus5_0\
        );

    \I__5180\ : InMux
    port map (
            O => \N__24048\,
            I => \N__24045\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__24042\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__24042\,
            I => \N__24039\
        );

    \I__5177\ : Span4Mux_h
    port map (
            O => \N__24039\,
            I => \N__24036\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__24036\,
            I => \this_sprites_ram.mem_out_bus1_0\
        );

    \I__5175\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24030\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__24030\,
            I => \N__24027\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__24027\,
            I => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\
        );

    \I__5172\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24021\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__24021\,
            I => \M_this_sprites_address_qc_0_0\
        );

    \I__5170\ : CEMux
    port map (
            O => \N__24018\,
            I => \N__24014\
        );

    \I__5169\ : CEMux
    port map (
            O => \N__24017\,
            I => \N__24011\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__24014\,
            I => \N__24008\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24005\
        );

    \I__5166\ : Span4Mux_s3_v
    port map (
            O => \N__24008\,
            I => \N__24002\
        );

    \I__5165\ : Span4Mux_h
    port map (
            O => \N__24005\,
            I => \N__23999\
        );

    \I__5164\ : Span4Mux_v
    port map (
            O => \N__24002\,
            I => \N__23994\
        );

    \I__5163\ : Span4Mux_v
    port map (
            O => \N__23999\,
            I => \N__23994\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__23994\,
            I => \N__23991\
        );

    \I__5161\ : Odrv4
    port map (
            O => \N__23991\,
            I => \this_sprites_ram.mem_WE_14\
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__23988\,
            I => \N__23981\
        );

    \I__5159\ : CascadeMux
    port map (
            O => \N__23987\,
            I => \N__23978\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__23986\,
            I => \N__23973\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__23985\,
            I => \N__23968\
        );

    \I__5156\ : CascadeMux
    port map (
            O => \N__23984\,
            I => \N__23965\
        );

    \I__5155\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23960\
        );

    \I__5154\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23957\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__23977\,
            I => \N__23954\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__23976\,
            I => \N__23951\
        );

    \I__5151\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23945\
        );

    \I__5150\ : CascadeMux
    port map (
            O => \N__23972\,
            I => \N__23942\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__23971\,
            I => \N__23939\
        );

    \I__5148\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23935\
        );

    \I__5147\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23932\
        );

    \I__5146\ : CascadeMux
    port map (
            O => \N__23964\,
            I => \N__23929\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__23963\,
            I => \N__23926\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__23960\,
            I => \N__23920\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__23957\,
            I => \N__23920\
        );

    \I__5142\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23917\
        );

    \I__5141\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23914\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__23950\,
            I => \N__23911\
        );

    \I__5139\ : CascadeMux
    port map (
            O => \N__23949\,
            I => \N__23908\
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__23948\,
            I => \N__23905\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23902\
        );

    \I__5136\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23899\
        );

    \I__5135\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23896\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__23938\,
            I => \N__23893\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23890\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__23932\,
            I => \N__23887\
        );

    \I__5131\ : InMux
    port map (
            O => \N__23929\,
            I => \N__23884\
        );

    \I__5130\ : InMux
    port map (
            O => \N__23926\,
            I => \N__23881\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__23925\,
            I => \N__23878\
        );

    \I__5128\ : Span4Mux_v
    port map (
            O => \N__23920\,
            I => \N__23871\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__23917\,
            I => \N__23871\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__23914\,
            I => \N__23871\
        );

    \I__5125\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23868\
        );

    \I__5124\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23865\
        );

    \I__5123\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23862\
        );

    \I__5122\ : Span4Mux_v
    port map (
            O => \N__23902\,
            I => \N__23855\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__23899\,
            I => \N__23855\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__23896\,
            I => \N__23855\
        );

    \I__5119\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23852\
        );

    \I__5118\ : Span4Mux_v
    port map (
            O => \N__23890\,
            I => \N__23845\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__23887\,
            I => \N__23845\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__23884\,
            I => \N__23845\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__23881\,
            I => \N__23842\
        );

    \I__5114\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23839\
        );

    \I__5113\ : Span4Mux_v
    port map (
            O => \N__23871\,
            I => \N__23832\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__23868\,
            I => \N__23832\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__23865\,
            I => \N__23832\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__23862\,
            I => \N__23825\
        );

    \I__5109\ : Span4Mux_v
    port map (
            O => \N__23855\,
            I => \N__23825\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__23852\,
            I => \N__23825\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__23845\,
            I => \N__23819\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__23842\,
            I => \N__23819\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23816\
        );

    \I__5104\ : Span4Mux_v
    port map (
            O => \N__23832\,
            I => \N__23811\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__23825\,
            I => \N__23811\
        );

    \I__5102\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23808\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__23819\,
            I => \N__23805\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__23816\,
            I => \N__23802\
        );

    \I__5099\ : Span4Mux_h
    port map (
            O => \N__23811\,
            I => \N__23796\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__23808\,
            I => \N__23796\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__23805\,
            I => \N__23793\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__23802\,
            I => \N__23790\
        );

    \I__5095\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23787\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__23796\,
            I => \N__23784\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__23793\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5092\ : Odrv4
    port map (
            O => \N__23790\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__23787\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__23784\,
            I => \M_this_sprites_address_qZ0Z_0\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__23775\,
            I => \N__23771\
        );

    \I__5088\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23768\
        );

    \I__5087\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23765\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N_443_i\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__23765\,
            I => \N_443_i\
        );

    \I__5084\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23757\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__23757\,
            I => \N__23754\
        );

    \I__5082\ : Span4Mux_v
    port map (
            O => \N__23754\,
            I => \N__23751\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__23751\,
            I => \N__23748\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__23748\,
            I => \M_this_sprites_address_q_RNO_0Z0Z_0\
        );

    \I__5079\ : InMux
    port map (
            O => \N__23745\,
            I => \un1_M_this_sprites_address_q_cry_0\
        );

    \I__5078\ : InMux
    port map (
            O => \N__23742\,
            I => \un1_M_this_sprites_address_q_cry_1\
        );

    \I__5077\ : InMux
    port map (
            O => \N__23739\,
            I => \un1_M_this_sprites_address_q_cry_2\
        );

    \I__5076\ : InMux
    port map (
            O => \N__23736\,
            I => \bfn_20_20_0_\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__5074\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__23727\,
            I => \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__23724\,
            I => \N__23721\
        );

    \I__5071\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23718\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__23718\,
            I => \N__23715\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__23715\,
            I => \N__23712\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__23712\,
            I => \N__23709\
        );

    \I__5067\ : Span4Mux_h
    port map (
            O => \N__23709\,
            I => \N__23706\
        );

    \I__5066\ : Span4Mux_h
    port map (
            O => \N__23706\,
            I => \N__23703\
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__23703\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__23700\,
            I => \N__23692\
        );

    \I__5063\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23688\
        );

    \I__5062\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23685\
        );

    \I__5061\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23682\
        );

    \I__5060\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23678\
        );

    \I__5059\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23675\
        );

    \I__5058\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23670\
        );

    \I__5057\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23670\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__23688\,
            I => \N__23663\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__23685\,
            I => \N__23663\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__23682\,
            I => \N__23663\
        );

    \I__5053\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23660\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__23678\,
            I => \N__23653\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__23675\,
            I => \N__23653\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__23670\,
            I => \N__23653\
        );

    \I__5049\ : Sp12to4
    port map (
            O => \N__23663\,
            I => \N__23646\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23646\
        );

    \I__5047\ : Sp12to4
    port map (
            O => \N__23653\,
            I => \N__23646\
        );

    \I__5046\ : Odrv12
    port map (
            O => \N__23646\,
            I => \this_sprites_ram.mem_radregZ0Z_11\
        );

    \I__5045\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23640\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__23640\,
            I => \N__23635\
        );

    \I__5043\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23632\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__23638\,
            I => \N__23629\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__23635\,
            I => \N__23624\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__23632\,
            I => \N__23624\
        );

    \I__5039\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23621\
        );

    \I__5038\ : Span4Mux_v
    port map (
            O => \N__23624\,
            I => \N__23612\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__23621\,
            I => \N__23612\
        );

    \I__5036\ : CascadeMux
    port map (
            O => \N__23620\,
            I => \N__23609\
        );

    \I__5035\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23601\
        );

    \I__5034\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23601\
        );

    \I__5033\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23601\
        );

    \I__5032\ : Span4Mux_v
    port map (
            O => \N__23612\,
            I => \N__23598\
        );

    \I__5031\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23595\
        );

    \I__5030\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23592\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__23601\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__23598\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__23595\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__23592\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__5025\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23571\
        );

    \I__5024\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23571\
        );

    \I__5023\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23571\
        );

    \I__5022\ : InMux
    port map (
            O => \N__23580\,
            I => \N__23571\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__23571\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5020\ : InMux
    port map (
            O => \N__23568\,
            I => \N__23564\
        );

    \I__5019\ : InMux
    port map (
            O => \N__23567\,
            I => \N__23561\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__23564\,
            I => \N__23558\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__23561\,
            I => \this_ppu.M_this_ppu_vram_addr_i_7\
        );

    \I__5016\ : Odrv4
    port map (
            O => \N__23558\,
            I => \this_ppu.M_this_ppu_vram_addr_i_7\
        );

    \I__5015\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23549\
        );

    \I__5014\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23546\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23543\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__23546\,
            I => \this_ppu.M_vaddress_q_i_1\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__23543\,
            I => \this_ppu.M_vaddress_q_i_1\
        );

    \I__5010\ : InMux
    port map (
            O => \N__23538\,
            I => \N__23534\
        );

    \I__5009\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23531\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23528\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__23531\,
            I => \this_ppu.M_vaddress_q_i_2\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__23528\,
            I => \this_ppu.M_vaddress_q_i_2\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__23523\,
            I => \N__23520\
        );

    \I__5004\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23516\
        );

    \I__5003\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23513\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__23516\,
            I => \N__23510\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__23513\,
            I => \this_ppu.M_this_ppu_map_addr_i_5\
        );

    \I__5000\ : Odrv4
    port map (
            O => \N__23510\,
            I => \this_ppu.M_this_ppu_map_addr_i_5\
        );

    \I__4999\ : CascadeMux
    port map (
            O => \N__23505\,
            I => \N__23502\
        );

    \I__4998\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23498\
        );

    \I__4997\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23495\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23492\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__23495\,
            I => \this_ppu.M_this_ppu_map_addr_i_6\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__23492\,
            I => \this_ppu.M_this_ppu_map_addr_i_6\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__23487\,
            I => \N__23484\
        );

    \I__4992\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23480\
        );

    \I__4991\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23477\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__23480\,
            I => \N__23474\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__23477\,
            I => \this_ppu.M_this_ppu_map_addr_i_7\
        );

    \I__4988\ : Odrv4
    port map (
            O => \N__23474\,
            I => \this_ppu.M_this_ppu_map_addr_i_7\
        );

    \I__4987\ : CascadeMux
    port map (
            O => \N__23469\,
            I => \N__23466\
        );

    \I__4986\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23462\
        );

    \I__4985\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23459\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__23462\,
            I => \N__23456\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__23459\,
            I => \this_ppu.M_this_ppu_map_addr_i_8\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__23456\,
            I => \this_ppu.M_this_ppu_map_addr_i_8\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__23451\,
            I => \N__23447\
        );

    \I__4980\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23444\
        );

    \I__4979\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23441\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23438\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__23441\,
            I => \this_ppu.M_this_ppu_map_addr_i_9\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__23438\,
            I => \this_ppu.M_this_ppu_map_addr_i_9\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__23433\,
            I => \N__23425\
        );

    \I__4974\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23422\
        );

    \I__4973\ : InMux
    port map (
            O => \N__23431\,
            I => \N__23419\
        );

    \I__4972\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23416\
        );

    \I__4971\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23411\
        );

    \I__4970\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23411\
        );

    \I__4969\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23408\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__23422\,
            I => \N__23405\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23398\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__23416\,
            I => \N__23398\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__23411\,
            I => \N__23398\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__23408\,
            I => \N__23395\
        );

    \I__4963\ : Span4Mux_h
    port map (
            O => \N__23405\,
            I => \N__23392\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__23398\,
            I => \N__23389\
        );

    \I__4961\ : Odrv12
    port map (
            O => \N__23395\,
            I => \N_775_0\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__23392\,
            I => \N_775_0\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__23389\,
            I => \N_775_0\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__23382\,
            I => \N_775_0_cascade_\
        );

    \I__4957\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23376\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__23376\,
            I => \N__23373\
        );

    \I__4955\ : Span4Mux_h
    port map (
            O => \N__23373\,
            I => \N__23370\
        );

    \I__4954\ : Span4Mux_v
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__4953\ : Sp12to4
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__4952\ : Odrv12
    port map (
            O => \N__23364\,
            I => port_address_in_5
        );

    \I__4951\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23355\
        );

    \I__4950\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23355\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__23355\,
            I => \N__23352\
        );

    \I__4948\ : Odrv12
    port map (
            O => \N__23352\,
            I => \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0Z0Z_0\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__23349\,
            I => \N_87_0_cascade_\
        );

    \I__4946\ : CascadeMux
    port map (
            O => \N__23346\,
            I => \N__23339\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \N__23336\
        );

    \I__4944\ : CascadeMux
    port map (
            O => \N__23344\,
            I => \N__23333\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__23343\,
            I => \N__23330\
        );

    \I__4942\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23327\
        );

    \I__4941\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23324\
        );

    \I__4940\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23321\
        );

    \I__4939\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23316\
        );

    \I__4938\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23316\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23312\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__23324\,
            I => \N__23309\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23304\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__23316\,
            I => \N__23304\
        );

    \I__4933\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23301\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__23312\,
            I => \N__23294\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__23309\,
            I => \N__23294\
        );

    \I__4930\ : Span4Mux_v
    port map (
            O => \N__23304\,
            I => \N__23294\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__23301\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__23294\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__23289\,
            I => \N__23286\
        );

    \I__4926\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23274\
        );

    \I__4925\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23274\
        );

    \I__4924\ : InMux
    port map (
            O => \N__23284\,
            I => \N__23274\
        );

    \I__4923\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23274\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__4921\ : Span4Mux_v
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__4920\ : Span4Mux_h
    port map (
            O => \N__23268\,
            I => \N__23265\
        );

    \I__4919\ : Span4Mux_h
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__4918\ : Sp12to4
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__4917\ : Span12Mux_h
    port map (
            O => \N__23259\,
            I => \N__23256\
        );

    \I__4916\ : Odrv12
    port map (
            O => \N__23256\,
            I => port_enb_c
        );

    \I__4915\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23247\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__23247\,
            I => \N__23241\
        );

    \I__4912\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23234\
        );

    \I__4911\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23234\
        );

    \I__4910\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23234\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__23241\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__23234\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__4907\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23226\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__23226\,
            I => \this_reset_cond.M_stage_qZ0Z_4\
        );

    \I__4905\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23218\
        );

    \I__4904\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23214\
        );

    \I__4903\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23211\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__23218\,
            I => \N__23207\
        );

    \I__4901\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23204\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23197\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__23211\,
            I => \N__23197\
        );

    \I__4898\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23194\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__23207\,
            I => \N__23189\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__23204\,
            I => \N__23189\
        );

    \I__4895\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23186\
        );

    \I__4894\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23183\
        );

    \I__4893\ : Span4Mux_h
    port map (
            O => \N__23197\,
            I => \N__23180\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__23194\,
            I => \N__23175\
        );

    \I__4891\ : Span4Mux_h
    port map (
            O => \N__23189\,
            I => \N__23175\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__23186\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__23183\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__4888\ : Odrv4
    port map (
            O => \N__23180\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__23175\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__4886\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23163\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23160\
        );

    \I__4884\ : Odrv12
    port map (
            O => \N__23160\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__23157\,
            I => \N__23154\
        );

    \I__4882\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23151\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__23151\,
            I => \N_126\
        );

    \I__4880\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23145\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__23145\,
            I => \N__23141\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23134\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__23141\,
            I => \N__23131\
        );

    \I__4876\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23124\
        );

    \I__4875\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23124\
        );

    \I__4874\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23124\
        );

    \I__4873\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23121\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__23134\,
            I => \N__23118\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__23131\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__23124\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__23121\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4868\ : Odrv12
    port map (
            O => \N__23118\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__23109\,
            I => \port_dmab_ac0_1_3_cascade_\
        );

    \I__4866\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23103\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__23103\,
            I => port_dmab_ac0_1_4
        );

    \I__4864\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23096\
        );

    \I__4863\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23092\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__23096\,
            I => \N__23087\
        );

    \I__4861\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23084\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__23081\
        );

    \I__4859\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23078\
        );

    \I__4858\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23074\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__23087\,
            I => \N__23069\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23066\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__23081\,
            I => \N__23061\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__23078\,
            I => \N__23061\
        );

    \I__4853\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23058\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__23074\,
            I => \N__23055\
        );

    \I__4851\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23052\
        );

    \I__4850\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23049\
        );

    \I__4849\ : Span4Mux_v
    port map (
            O => \N__23069\,
            I => \N__23044\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__23066\,
            I => \N__23044\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__23061\,
            I => \N__23039\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23039\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__23055\,
            I => \N__23036\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23033\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__23049\,
            I => \N__23030\
        );

    \I__4842\ : Span4Mux_v
    port map (
            O => \N__23044\,
            I => \N__23027\
        );

    \I__4841\ : Sp12to4
    port map (
            O => \N__23039\,
            I => \N__23024\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__23036\,
            I => \N__23019\
        );

    \I__4839\ : Span4Mux_h
    port map (
            O => \N__23033\,
            I => \N__23019\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__23030\,
            I => \N__23016\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__23027\,
            I => \N__23013\
        );

    \I__4836\ : Span12Mux_v
    port map (
            O => \N__23024\,
            I => \N__23010\
        );

    \I__4835\ : Span4Mux_h
    port map (
            O => \N__23019\,
            I => \N__23005\
        );

    \I__4834\ : Span4Mux_h
    port map (
            O => \N__23016\,
            I => \N__23005\
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__23013\,
            I => \N_15\
        );

    \I__4832\ : Odrv12
    port map (
            O => \N__23010\,
            I => \N_15\
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__23005\,
            I => \N_15\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__22998\,
            I => \N_809_cascade_\
        );

    \I__4829\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22988\
        );

    \I__4828\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22985\
        );

    \I__4827\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22982\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__22992\,
            I => \N__22978\
        );

    \I__4825\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22975\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22972\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__22985\,
            I => \N__22969\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__22982\,
            I => \N__22966\
        );

    \I__4821\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22963\
        );

    \I__4820\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22960\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__22975\,
            I => \N__22957\
        );

    \I__4818\ : Span12Mux_h
    port map (
            O => \N__22972\,
            I => \N__22954\
        );

    \I__4817\ : Span4Mux_h
    port map (
            O => \N__22969\,
            I => \N__22949\
        );

    \I__4816\ : Span4Mux_h
    port map (
            O => \N__22966\,
            I => \N__22949\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__22963\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__22960\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__22957\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__4812\ : Odrv12
    port map (
            O => \N__22954\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__22949\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__4810\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22934\
        );

    \I__4809\ : InMux
    port map (
            O => \N__22937\,
            I => \N__22931\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22925\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__22931\,
            I => \N__22922\
        );

    \I__4806\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22919\
        );

    \I__4805\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22916\
        );

    \I__4804\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22913\
        );

    \I__4803\ : Span4Mux_h
    port map (
            O => \N__22925\,
            I => \N__22910\
        );

    \I__4802\ : Span4Mux_h
    port map (
            O => \N__22922\,
            I => \N__22907\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__22919\,
            I => \N__22902\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22902\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__22913\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__22910\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__22907\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4796\ : Odrv12
    port map (
            O => \N__22902\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__4795\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22889\
        );

    \I__4794\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22886\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__22889\,
            I => \N__22883\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__22886\,
            I => \N__22878\
        );

    \I__4791\ : Span4Mux_h
    port map (
            O => \N__22883\,
            I => \N__22875\
        );

    \I__4790\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22870\
        );

    \I__4789\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22870\
        );

    \I__4788\ : Odrv12
    port map (
            O => \N__22878\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__22875\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__22870\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__22863\,
            I => \N__22860\
        );

    \I__4784\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22857\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N_792\
        );

    \I__4782\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__22851\,
            I => \M_this_sprites_address_qc_0_0_0\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__4779\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__22842\,
            I => \N_795\
        );

    \I__4777\ : CascadeMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__4776\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__22830\,
            I => \N_773_0\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__22827\,
            I => \N_773_0_cascade_\
        );

    \I__4772\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22821\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__22821\,
            I => \this_vga_signals.N_485\
        );

    \I__4770\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22814\
        );

    \I__4769\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22808\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__22814\,
            I => \N__22804\
        );

    \I__4767\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22801\
        );

    \I__4766\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22797\
        );

    \I__4765\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22794\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__22808\,
            I => \N__22790\
        );

    \I__4763\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22787\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__22804\,
            I => \N__22782\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__22801\,
            I => \N__22782\
        );

    \I__4760\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22779\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__22797\,
            I => \N__22776\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22773\
        );

    \I__4757\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22770\
        );

    \I__4756\ : Sp12to4
    port map (
            O => \N__22790\,
            I => \N__22765\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__22787\,
            I => \N__22765\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__22782\,
            I => \N__22760\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__22779\,
            I => \N__22760\
        );

    \I__4752\ : Span4Mux_h
    port map (
            O => \N__22776\,
            I => \N__22757\
        );

    \I__4751\ : Span4Mux_h
    port map (
            O => \N__22773\,
            I => \N__22754\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__22770\,
            I => \N__22751\
        );

    \I__4749\ : Span12Mux_v
    port map (
            O => \N__22765\,
            I => \N__22748\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__22760\,
            I => \N__22745\
        );

    \I__4747\ : Span4Mux_v
    port map (
            O => \N__22757\,
            I => \N__22738\
        );

    \I__4746\ : Span4Mux_v
    port map (
            O => \N__22754\,
            I => \N__22738\
        );

    \I__4745\ : Span4Mux_h
    port map (
            O => \N__22751\,
            I => \N__22738\
        );

    \I__4744\ : Span12Mux_h
    port map (
            O => \N__22748\,
            I => \N__22735\
        );

    \I__4743\ : Span4Mux_h
    port map (
            O => \N__22745\,
            I => \N__22732\
        );

    \I__4742\ : Span4Mux_h
    port map (
            O => \N__22738\,
            I => \N__22729\
        );

    \I__4741\ : Odrv12
    port map (
            O => \N__22735\,
            I => \N_17\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__22732\,
            I => \N_17\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__22729\,
            I => \N_17\
        );

    \I__4738\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22719\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__22719\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__22716\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\
        );

    \I__4735\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__22710\,
            I => \N__22707\
        );

    \I__4733\ : Span12Mux_s9_v
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__4732\ : Span12Mux_h
    port map (
            O => \N__22704\,
            I => \N__22700\
        );

    \I__4731\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22697\
        );

    \I__4730\ : Odrv12
    port map (
            O => \N__22700\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__22697\,
            I => \M_this_ppu_vram_data_1\
        );

    \I__4728\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22689\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__22689\,
            I => \N__22686\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__22686\,
            I => \N__22683\
        );

    \I__4725\ : Span4Mux_v
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__4724\ : Span4Mux_h
    port map (
            O => \N__22680\,
            I => \N__22677\
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__22677\,
            I => \this_sprites_ram.mem_out_bus7_2\
        );

    \I__4722\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22671\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__22671\,
            I => \N__22668\
        );

    \I__4720\ : Span4Mux_v
    port map (
            O => \N__22668\,
            I => \N__22665\
        );

    \I__4719\ : Sp12to4
    port map (
            O => \N__22665\,
            I => \N__22662\
        );

    \I__4718\ : Odrv12
    port map (
            O => \N__22662\,
            I => \this_sprites_ram.mem_out_bus3_2\
        );

    \I__4717\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__4715\ : Span12Mux_v
    port map (
            O => \N__22653\,
            I => \N__22650\
        );

    \I__4714\ : Odrv12
    port map (
            O => \N__22650\,
            I => \this_sprites_ram.mem_out_bus4_2\
        );

    \I__4713\ : InMux
    port map (
            O => \N__22647\,
            I => \N__22644\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__22644\,
            I => \N__22641\
        );

    \I__4711\ : Span4Mux_v
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__22638\,
            I => \N__22635\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__22635\,
            I => \this_sprites_ram.mem_out_bus0_2\
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__22632\,
            I => \N__22629\
        );

    \I__4707\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22625\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__22628\,
            I => \N__22621\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__22625\,
            I => \N__22617\
        );

    \I__4704\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22614\
        );

    \I__4703\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22611\
        );

    \I__4702\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22608\
        );

    \I__4701\ : Span4Mux_v
    port map (
            O => \N__22617\,
            I => \N__22605\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__22614\,
            I => \N__22602\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__22611\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__22608\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__22605\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__22602\,
            I => \this_sprites_ram.mem_radregZ0Z_12\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__22593\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\
        );

    \I__4694\ : InMux
    port map (
            O => \N__22590\,
            I => \N__22587\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__22587\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__22584\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\
        );

    \I__4691\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__22578\,
            I => \N__22575\
        );

    \I__4689\ : Span12Mux_s9_v
    port map (
            O => \N__22575\,
            I => \N__22572\
        );

    \I__4688\ : Span12Mux_h
    port map (
            O => \N__22572\,
            I => \N__22568\
        );

    \I__4687\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22565\
        );

    \I__4686\ : Odrv12
    port map (
            O => \N__22568\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__22565\,
            I => \M_this_ppu_vram_data_2\
        );

    \I__4684\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22557\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__22557\,
            I => \N__22554\
        );

    \I__4682\ : Span4Mux_v
    port map (
            O => \N__22554\,
            I => \N__22551\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__22551\,
            I => \N__22548\
        );

    \I__4680\ : Sp12to4
    port map (
            O => \N__22548\,
            I => \N__22545\
        );

    \I__4679\ : Span12Mux_v
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__4678\ : Span12Mux_h
    port map (
            O => \N__22542\,
            I => \N__22539\
        );

    \I__4677\ : Odrv12
    port map (
            O => \N__22539\,
            I => \M_this_map_ram_read_data_0\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__22536\,
            I => \N__22532\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__22535\,
            I => \N__22521\
        );

    \I__4674\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22518\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__22531\,
            I => \N__22515\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__22530\,
            I => \N__22512\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__22529\,
            I => \N__22508\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__22528\,
            I => \N__22503\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__22527\,
            I => \N__22500\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__22526\,
            I => \N__22497\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__22525\,
            I => \N__22494\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__22524\,
            I => \N__22491\
        );

    \I__4665\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22488\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__22518\,
            I => \N__22484\
        );

    \I__4663\ : InMux
    port map (
            O => \N__22515\,
            I => \N__22481\
        );

    \I__4662\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22477\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__22511\,
            I => \N__22474\
        );

    \I__4660\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22471\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__22507\,
            I => \N__22468\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__22506\,
            I => \N__22465\
        );

    \I__4657\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22461\
        );

    \I__4656\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22458\
        );

    \I__4655\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22455\
        );

    \I__4654\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22452\
        );

    \I__4653\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22449\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__22488\,
            I => \N__22446\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__22487\,
            I => \N__22443\
        );

    \I__4650\ : Span4Mux_v
    port map (
            O => \N__22484\,
            I => \N__22438\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__22481\,
            I => \N__22438\
        );

    \I__4648\ : CascadeMux
    port map (
            O => \N__22480\,
            I => \N__22435\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__22477\,
            I => \N__22432\
        );

    \I__4646\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22429\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__22471\,
            I => \N__22426\
        );

    \I__4644\ : InMux
    port map (
            O => \N__22468\,
            I => \N__22423\
        );

    \I__4643\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22420\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__22464\,
            I => \N__22417\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__22461\,
            I => \N__22414\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22405\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__22455\,
            I => \N__22405\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__22452\,
            I => \N__22405\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__22449\,
            I => \N__22405\
        );

    \I__4636\ : Span4Mux_s2_v
    port map (
            O => \N__22446\,
            I => \N__22402\
        );

    \I__4635\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22399\
        );

    \I__4634\ : Span4Mux_v
    port map (
            O => \N__22438\,
            I => \N__22396\
        );

    \I__4633\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22393\
        );

    \I__4632\ : Span4Mux_h
    port map (
            O => \N__22432\,
            I => \N__22390\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__22429\,
            I => \N__22387\
        );

    \I__4630\ : Span4Mux_h
    port map (
            O => \N__22426\,
            I => \N__22384\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__22423\,
            I => \N__22381\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22378\
        );

    \I__4627\ : InMux
    port map (
            O => \N__22417\,
            I => \N__22375\
        );

    \I__4626\ : Span4Mux_h
    port map (
            O => \N__22414\,
            I => \N__22372\
        );

    \I__4625\ : Span12Mux_v
    port map (
            O => \N__22405\,
            I => \N__22369\
        );

    \I__4624\ : Sp12to4
    port map (
            O => \N__22402\,
            I => \N__22364\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__22399\,
            I => \N__22364\
        );

    \I__4622\ : Sp12to4
    port map (
            O => \N__22396\,
            I => \N__22359\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22359\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__22390\,
            I => \N__22354\
        );

    \I__4619\ : Span4Mux_h
    port map (
            O => \N__22387\,
            I => \N__22354\
        );

    \I__4618\ : Span4Mux_v
    port map (
            O => \N__22384\,
            I => \N__22349\
        );

    \I__4617\ : Span4Mux_h
    port map (
            O => \N__22381\,
            I => \N__22349\
        );

    \I__4616\ : Span4Mux_h
    port map (
            O => \N__22378\,
            I => \N__22346\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__22375\,
            I => \N__22343\
        );

    \I__4614\ : Sp12to4
    port map (
            O => \N__22372\,
            I => \N__22340\
        );

    \I__4613\ : Span12Mux_h
    port map (
            O => \N__22369\,
            I => \N__22333\
        );

    \I__4612\ : Span12Mux_h
    port map (
            O => \N__22364\,
            I => \N__22333\
        );

    \I__4611\ : Span12Mux_h
    port map (
            O => \N__22359\,
            I => \N__22333\
        );

    \I__4610\ : Span4Mux_h
    port map (
            O => \N__22354\,
            I => \N__22328\
        );

    \I__4609\ : Span4Mux_h
    port map (
            O => \N__22349\,
            I => \N__22328\
        );

    \I__4608\ : Span4Mux_v
    port map (
            O => \N__22346\,
            I => \N__22323\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__22343\,
            I => \N__22323\
        );

    \I__4606\ : Odrv12
    port map (
            O => \N__22340\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__4605\ : Odrv12
    port map (
            O => \N__22333\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__22328\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__4603\ : Odrv4
    port map (
            O => \N__22323\,
            I => \M_this_ppu_sprites_addr_6\
        );

    \I__4602\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22308\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__22302\,
            I => \this_sprites_ram.mem_out_bus6_2\
        );

    \I__4597\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22296\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__4595\ : Span12Mux_v
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__4594\ : Odrv12
    port map (
            O => \N__22290\,
            I => \this_sprites_ram.mem_out_bus2_2\
        );

    \I__4593\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__22284\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\
        );

    \I__4591\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22277\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22274\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__22277\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__22274\,
            I => \this_ppu.M_this_ppu_map_addr_i_3\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__22269\,
            I => \N__22266\
        );

    \I__4586\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22262\
        );

    \I__4585\ : InMux
    port map (
            O => \N__22265\,
            I => \N__22259\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__22262\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__22259\,
            I => \this_ppu.M_this_ppu_map_addr_i_4\
        );

    \I__4582\ : InMux
    port map (
            O => \N__22254\,
            I => \bfn_19_20_0_\
        );

    \I__4581\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22248\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__22248\,
            I => \this_ppu.vscroll8_1\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__4578\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__4576\ : Span4Mux_v
    port map (
            O => \N__22236\,
            I => \N__22233\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__22233\,
            I => \N__22230\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__22230\,
            I => \this_ppu.un1_M_vaddress_q_3_4\
        );

    \I__4573\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22224\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__22224\,
            I => \N__22221\
        );

    \I__4571\ : Span12Mux_v
    port map (
            O => \N__22221\,
            I => \N__22218\
        );

    \I__4570\ : Span12Mux_h
    port map (
            O => \N__22218\,
            I => \N__22215\
        );

    \I__4569\ : Odrv12
    port map (
            O => \N__22215\,
            I => \this_sprites_ram.mem_out_bus4_1\
        );

    \I__4568\ : InMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__22209\,
            I => \N__22206\
        );

    \I__4566\ : Span4Mux_v
    port map (
            O => \N__22206\,
            I => \N__22203\
        );

    \I__4565\ : Span4Mux_h
    port map (
            O => \N__22203\,
            I => \N__22200\
        );

    \I__4564\ : Span4Mux_v
    port map (
            O => \N__22200\,
            I => \N__22197\
        );

    \I__4563\ : Odrv4
    port map (
            O => \N__22197\,
            I => \this_sprites_ram.mem_out_bus0_1\
        );

    \I__4562\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22191\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__22191\,
            I => \N__22188\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__22188\,
            I => \N__22185\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__22185\,
            I => \N__22182\
        );

    \I__4558\ : Span4Mux_h
    port map (
            O => \N__22182\,
            I => \N__22179\
        );

    \I__4557\ : Odrv4
    port map (
            O => \N__22179\,
            I => \this_sprites_ram.mem_out_bus7_1\
        );

    \I__4556\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22173\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__22173\,
            I => \N__22170\
        );

    \I__4554\ : Sp12to4
    port map (
            O => \N__22170\,
            I => \N__22167\
        );

    \I__4553\ : Odrv12
    port map (
            O => \N__22167\,
            I => \this_sprites_ram.mem_out_bus3_1\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__22164\,
            I => \N__22161\
        );

    \I__4551\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22158\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__22158\,
            I => \N__22155\
        );

    \I__4549\ : Span12Mux_v
    port map (
            O => \N__22155\,
            I => \N__22152\
        );

    \I__4548\ : Span12Mux_h
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__4547\ : Odrv12
    port map (
            O => \N__22149\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__4546\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22143\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__22143\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__4543\ : CascadeBuf
    port map (
            O => \N__22137\,
            I => \N__22134\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__22134\,
            I => \N__22131\
        );

    \I__4541\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22128\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__4539\ : Sp12to4
    port map (
            O => \N__22125\,
            I => \N__22120\
        );

    \I__4538\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22117\
        );

    \I__4537\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22114\
        );

    \I__4536\ : Span12Mux_v
    port map (
            O => \N__22120\,
            I => \N__22111\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__22117\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__22114\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__4533\ : Odrv12
    port map (
            O => \N__22111\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__4532\ : InMux
    port map (
            O => \N__22104\,
            I => \bfn_19_18_0_\
        );

    \I__4531\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22098\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__22095\,
            I => \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\
        );

    \I__4528\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__22086\,
            I => \N__22083\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__22083\,
            I => \this_reset_cond.M_stage_qZ0Z_3\
        );

    \I__4524\ : InMux
    port map (
            O => \N__22080\,
            I => \N__22076\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22073\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__22076\,
            I => \this_ppu.M_this_ppu_vram_addr_i_0\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__22073\,
            I => \this_ppu.M_this_ppu_vram_addr_i_0\
        );

    \I__4520\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22064\
        );

    \I__4519\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22061\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__22064\,
            I => \this_ppu.M_this_ppu_vram_addr_i_1\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__22061\,
            I => \this_ppu.M_this_ppu_vram_addr_i_1\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__22056\,
            I => \N__22053\
        );

    \I__4515\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22050\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__22050\,
            I => \N__22046\
        );

    \I__4513\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22043\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__22046\,
            I => \this_ppu.M_this_ppu_vram_addr_i_2\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__22043\,
            I => \this_ppu.M_this_ppu_vram_addr_i_2\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__22038\,
            I => \N__22034\
        );

    \I__4509\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22031\
        );

    \I__4508\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22028\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__22031\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__22028\,
            I => \this_ppu.M_this_ppu_map_addr_i_0\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__22023\,
            I => \N__22019\
        );

    \I__4504\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22016\
        );

    \I__4503\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22013\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__22016\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__22013\,
            I => \this_ppu.M_this_ppu_map_addr_i_1\
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__22008\,
            I => \N__22004\
        );

    \I__4499\ : InMux
    port map (
            O => \N__22007\,
            I => \N__22001\
        );

    \I__4498\ : InMux
    port map (
            O => \N__22004\,
            I => \N__21998\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__22001\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__21998\,
            I => \this_ppu.M_this_ppu_map_addr_i_2\
        );

    \I__4495\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21987\
        );

    \I__4494\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21987\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21984\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__21984\,
            I => \this_ppu.un1_M_vaddress_q_2_c2\
        );

    \I__4491\ : SRMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__4489\ : Span4Mux_v
    port map (
            O => \N__21975\,
            I => \N__21971\
        );

    \I__4488\ : SRMux
    port map (
            O => \N__21974\,
            I => \N__21968\
        );

    \I__4487\ : Span4Mux_h
    port map (
            O => \N__21971\,
            I => \N__21963\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21963\
        );

    \I__4485\ : Span4Mux_h
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__21960\,
            I => \this_ppu.M_state_q_RNILG0GDZ0Z_0\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__21957\,
            I => \N__21954\
        );

    \I__4482\ : CascadeBuf
    port map (
            O => \N__21954\,
            I => \N__21951\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__4480\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21945\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__21945\,
            I => \N__21942\
        );

    \I__4478\ : Sp12to4
    port map (
            O => \N__21942\,
            I => \N__21938\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__21941\,
            I => \N__21935\
        );

    \I__4476\ : Span12Mux_s4_v
    port map (
            O => \N__21938\,
            I => \N__21929\
        );

    \I__4475\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21924\
        );

    \I__4474\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21924\
        );

    \I__4473\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21921\
        );

    \I__4472\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21918\
        );

    \I__4471\ : Span12Mux_v
    port map (
            O => \N__21929\,
            I => \N__21915\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__21924\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__21921\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__21918\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__4467\ : Odrv12
    port map (
            O => \N__21915\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__4465\ : CascadeBuf
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__21900\,
            I => \N__21897\
        );

    \I__4463\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__21894\,
            I => \N__21888\
        );

    \I__4461\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21885\
        );

    \I__4460\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21882\
        );

    \I__4459\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21879\
        );

    \I__4458\ : Span12Mux_v
    port map (
            O => \N__21888\,
            I => \N__21876\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__21885\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__21882\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__21879\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__4454\ : Odrv12
    port map (
            O => \N__21876\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__21867\,
            I => \N__21864\
        );

    \I__4452\ : CascadeBuf
    port map (
            O => \N__21864\,
            I => \N__21861\
        );

    \I__4451\ : CascadeMux
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__4450\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21855\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__21855\,
            I => \N__21852\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__4447\ : Span4Mux_v
    port map (
            O => \N__21849\,
            I => \N__21846\
        );

    \I__4446\ : Span4Mux_v
    port map (
            O => \N__21846\,
            I => \N__21839\
        );

    \I__4445\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21832\
        );

    \I__4444\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21832\
        );

    \I__4443\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21832\
        );

    \I__4442\ : InMux
    port map (
            O => \N__21842\,
            I => \N__21829\
        );

    \I__4441\ : Sp12to4
    port map (
            O => \N__21839\,
            I => \N__21826\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__21832\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__21829\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4438\ : Odrv12
    port map (
            O => \N__21826\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__21819\,
            I => \N__21816\
        );

    \I__4436\ : CascadeBuf
    port map (
            O => \N__21816\,
            I => \N__21813\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__21813\,
            I => \N__21810\
        );

    \I__4434\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21806\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__21809\,
            I => \N__21803\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__21806\,
            I => \N__21798\
        );

    \I__4431\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21793\
        );

    \I__4430\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21793\
        );

    \I__4429\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21790\
        );

    \I__4428\ : Span12Mux_v
    port map (
            O => \N__21798\,
            I => \N__21787\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__21793\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__21790\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__4425\ : Odrv12
    port map (
            O => \N__21787\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__21780\,
            I => \this_vga_signals.M_this_state_q_srsts_i_a3_0_7_cascade_\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__21777\,
            I => \this_vga_signals.M_this_state_q_srsts_i_0Z0Z_7_cascade_\
        );

    \I__4422\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21771\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__21771\,
            I => \N__21768\
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__21768\,
            I => \M_this_state_q_RNI6Q0SZ0Z_5\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__21765\,
            I => \N__21762\
        );

    \I__4418\ : InMux
    port map (
            O => \N__21762\,
            I => \N__21759\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__21759\,
            I => \N__21753\
        );

    \I__4416\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21750\
        );

    \I__4415\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21747\
        );

    \I__4414\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21744\
        );

    \I__4413\ : Span4Mux_v
    port map (
            O => \N__21753\,
            I => \N__21741\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__21750\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__21747\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__21744\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__21741\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__4408\ : InMux
    port map (
            O => \N__21732\,
            I => \N__21723\
        );

    \I__4407\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21723\
        );

    \I__4406\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21717\
        );

    \I__4405\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21714\
        );

    \I__4404\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21711\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__21723\,
            I => \N__21708\
        );

    \I__4402\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21703\
        );

    \I__4401\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21703\
        );

    \I__4400\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21700\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__21717\,
            I => \N_848\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__21714\,
            I => \N_848\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__21711\,
            I => \N_848\
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__21708\,
            I => \N_848\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__21703\,
            I => \N_848\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__21700\,
            I => \N_848\
        );

    \I__4393\ : InMux
    port map (
            O => \N__21687\,
            I => \N__21681\
        );

    \I__4392\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21681\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__21681\,
            I => \this_vga_signals.N_93_0\
        );

    \I__4390\ : InMux
    port map (
            O => \N__21678\,
            I => \N__21675\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__21675\,
            I => \N__21670\
        );

    \I__4388\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21667\
        );

    \I__4387\ : CascadeMux
    port map (
            O => \N__21673\,
            I => \N__21664\
        );

    \I__4386\ : Span4Mux_v
    port map (
            O => \N__21670\,
            I => \N__21658\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21655\
        );

    \I__4384\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21648\
        );

    \I__4383\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21648\
        );

    \I__4382\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21648\
        );

    \I__4381\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21645\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__21658\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__21655\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__21648\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__21645\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__4376\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21633\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__4374\ : Span4Mux_v
    port map (
            O => \N__21630\,
            I => \N__21624\
        );

    \I__4373\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21617\
        );

    \I__4372\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21617\
        );

    \I__4371\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21617\
        );

    \I__4370\ : Span4Mux_h
    port map (
            O => \N__21624\,
            I => \N__21611\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__21617\,
            I => \N__21611\
        );

    \I__4368\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21608\
        );

    \I__4367\ : Odrv4
    port map (
            O => \N__21611\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__21608\,
            I => \M_this_vga_signals_line_clk_0\
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__21603\,
            I => \N__21599\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__21602\,
            I => \N__21596\
        );

    \I__4363\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21593\
        );

    \I__4362\ : InMux
    port map (
            O => \N__21596\,
            I => \N__21588\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__21593\,
            I => \N__21585\
        );

    \I__4360\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21580\
        );

    \I__4359\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21580\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__21588\,
            I => \N__21577\
        );

    \I__4357\ : Span12Mux_v
    port map (
            O => \N__21585\,
            I => \N__21572\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__21580\,
            I => \N__21567\
        );

    \I__4355\ : Span4Mux_h
    port map (
            O => \N__21577\,
            I => \N__21567\
        );

    \I__4354\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21564\
        );

    \I__4353\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21561\
        );

    \I__4352\ : Odrv12
    port map (
            O => \N__21572\,
            I => \this_ppu.M_last_q\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__21567\,
            I => \this_ppu.M_last_q\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__21564\,
            I => \this_ppu.M_last_q\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__21561\,
            I => \this_ppu.M_last_q\
        );

    \I__4348\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21543\
        );

    \I__4347\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21543\
        );

    \I__4346\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21538\
        );

    \I__4345\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21538\
        );

    \I__4344\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21535\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__21543\,
            I => \N__21528\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__21538\,
            I => \N__21528\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__21535\,
            I => \N__21524\
        );

    \I__4340\ : InMux
    port map (
            O => \N__21534\,
            I => \N__21521\
        );

    \I__4339\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21518\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__21528\,
            I => \N__21515\
        );

    \I__4337\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21512\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__21524\,
            I => \N__21509\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__21521\,
            I => \N__21502\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21502\
        );

    \I__4333\ : Span4Mux_h
    port map (
            O => \N__21515\,
            I => \N__21502\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__21512\,
            I => \this_ppu.N_132_0\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__21509\,
            I => \this_ppu.N_132_0\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__21502\,
            I => \this_ppu.N_132_0\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__21495\,
            I => \M_this_state_q_RNIH92SZ0Z_10_cascade_\
        );

    \I__4328\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21488\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__21491\,
            I => \N__21485\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__21488\,
            I => \N__21480\
        );

    \I__4325\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21477\
        );

    \I__4324\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21471\
        );

    \I__4323\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21471\
        );

    \I__4322\ : Span4Mux_v
    port map (
            O => \N__21480\,
            I => \N__21464\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__21477\,
            I => \N__21464\
        );

    \I__4320\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21461\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__21471\,
            I => \N__21458\
        );

    \I__4318\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21453\
        );

    \I__4317\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21453\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__21464\,
            I => \this_vga_signals.N_83\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__21461\,
            I => \this_vga_signals.N_83\
        );

    \I__4314\ : Odrv12
    port map (
            O => \N__21458\,
            I => \this_vga_signals.N_83\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__21453\,
            I => \this_vga_signals.N_83\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__21444\,
            I => \N__21441\
        );

    \I__4311\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21438\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__21438\,
            I => \N__21435\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__21435\,
            I => \N__21432\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__21432\,
            I => \this_vga_signals.N_94_0\
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__21429\,
            I => \this_vga_signals.N_94_0_cascade_\
        );

    \I__4306\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__21423\,
            I => \this_vga_signals.M_this_state_q_srsts_i_i_0Z0Z_12\
        );

    \I__4304\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21414\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__21414\,
            I => \M_this_state_q_RNI373A1Z0Z_8\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__21411\,
            I => \this_vga_signals_un21_i_a3_1_1_cascade_\
        );

    \I__4300\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21405\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__21405\,
            I => \N__21401\
        );

    \I__4298\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21397\
        );

    \I__4297\ : Span4Mux_h
    port map (
            O => \N__21401\,
            I => \N__21394\
        );

    \I__4296\ : IoInMux
    port map (
            O => \N__21400\,
            I => \N__21391\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21388\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__21394\,
            I => \N__21385\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__21391\,
            I => \N__21381\
        );

    \I__4292\ : Sp12to4
    port map (
            O => \N__21388\,
            I => \N__21378\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__21385\,
            I => \N__21375\
        );

    \I__4290\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21372\
        );

    \I__4289\ : Span12Mux_s6_h
    port map (
            O => \N__21381\,
            I => \N__21368\
        );

    \I__4288\ : Span12Mux_v
    port map (
            O => \N__21378\,
            I => \N__21365\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__21375\,
            I => \N__21362\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__21372\,
            I => \N__21359\
        );

    \I__4285\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21356\
        );

    \I__4284\ : Span12Mux_h
    port map (
            O => \N__21368\,
            I => \N__21353\
        );

    \I__4283\ : Span12Mux_h
    port map (
            O => \N__21365\,
            I => \N__21350\
        );

    \I__4282\ : Span4Mux_h
    port map (
            O => \N__21362\,
            I => \N__21345\
        );

    \I__4281\ : Span4Mux_v
    port map (
            O => \N__21359\,
            I => \N__21345\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21342\
        );

    \I__4279\ : Odrv12
    port map (
            O => \N__21353\,
            I => port_dmab_c
        );

    \I__4278\ : Odrv12
    port map (
            O => \N__21350\,
            I => port_dmab_c
        );

    \I__4277\ : Odrv4
    port map (
            O => \N__21345\,
            I => port_dmab_c
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__21342\,
            I => port_dmab_c
        );

    \I__4275\ : InMux
    port map (
            O => \N__21333\,
            I => \N__21329\
        );

    \I__4274\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21325\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N__21322\
        );

    \I__4272\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21319\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__21325\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__21322\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__21319\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__4268\ : CascadeMux
    port map (
            O => \N__21312\,
            I => \N__21309\
        );

    \I__4267\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21305\
        );

    \I__4266\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21302\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21296\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__21302\,
            I => \N__21296\
        );

    \I__4263\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21293\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__21296\,
            I => \N__21290\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__21293\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__21290\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__21285\,
            I => \N__21282\
        );

    \I__4258\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21277\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__21281\,
            I => \N__21274\
        );

    \I__4256\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21271\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__21277\,
            I => \N__21268\
        );

    \I__4254\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21265\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__21271\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4252\ : Odrv4
    port map (
            O => \N__21268\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__21265\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__4250\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21253\
        );

    \I__4249\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21250\
        );

    \I__4248\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21247\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__21253\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__21250\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__21247\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__4244\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__4242\ : Odrv4
    port map (
            O => \N__21234\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_8\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__21231\,
            I => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_\
        );

    \I__4240\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21225\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__21225\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__21222\,
            I => \N__21219\
        );

    \I__4237\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21216\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__21216\,
            I => \N__21213\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__21213\,
            I => \N__21210\
        );

    \I__4234\ : Sp12to4
    port map (
            O => \N__21210\,
            I => \N__21207\
        );

    \I__4233\ : Span12Mux_v
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__4232\ : Span12Mux_h
    port map (
            O => \N__21204\,
            I => \N__21201\
        );

    \I__4231\ : Odrv12
    port map (
            O => \N__21201\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__4230\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21195\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__21195\,
            I => \N__21192\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21186\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__21186\,
            I => \N__21183\
        );

    \I__4225\ : Span4Mux_h
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__21180\,
            I => \this_sprites_ram.mem_out_bus7_3\
        );

    \I__4223\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21174\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21171\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__21171\,
            I => \N__21168\
        );

    \I__4220\ : Span4Mux_h
    port map (
            O => \N__21168\,
            I => \N__21165\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__21165\,
            I => \N__21162\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__21162\,
            I => \this_sprites_ram.mem_out_bus3_3\
        );

    \I__4217\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__21156\,
            I => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\
        );

    \I__4215\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__21150\,
            I => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\
        );

    \I__4213\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__21144\,
            I => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__21141\,
            I => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\
        );

    \I__4210\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__4208\ : Span4Mux_v
    port map (
            O => \N__21132\,
            I => \N__21129\
        );

    \I__4207\ : Sp12to4
    port map (
            O => \N__21129\,
            I => \N__21126\
        );

    \I__4206\ : Span12Mux_h
    port map (
            O => \N__21126\,
            I => \N__21122\
        );

    \I__4205\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21119\
        );

    \I__4204\ : Odrv12
    port map (
            O => \N__21122\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__21119\,
            I => \M_this_ppu_vram_data_3\
        );

    \I__4202\ : InMux
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__21111\,
            I => \N__21106\
        );

    \I__4200\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21103\
        );

    \I__4199\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21100\
        );

    \I__4198\ : Odrv12
    port map (
            O => \N__21106\,
            I => \this_ppu.N_156\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__21103\,
            I => \this_ppu.N_156\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__21100\,
            I => \this_ppu.N_156\
        );

    \I__4195\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__21090\,
            I => \this_ppu.N_150\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__21087\,
            I => \N__21083\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__21086\,
            I => \N__21080\
        );

    \I__4191\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21074\
        );

    \I__4190\ : InMux
    port map (
            O => \N__21080\,
            I => \N__21069\
        );

    \I__4189\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21069\
        );

    \I__4188\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21066\
        );

    \I__4187\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21063\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__21074\,
            I => \N__21060\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__21069\,
            I => \N__21057\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21054\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__21063\,
            I => \N__21051\
        );

    \I__4182\ : Span4Mux_h
    port map (
            O => \N__21060\,
            I => \N__21048\
        );

    \I__4181\ : Span4Mux_v
    port map (
            O => \N__21057\,
            I => \N__21045\
        );

    \I__4180\ : Span4Mux_h
    port map (
            O => \N__21054\,
            I => \N__21040\
        );

    \I__4179\ : Span4Mux_h
    port map (
            O => \N__21051\,
            I => \N__21040\
        );

    \I__4178\ : Span4Mux_v
    port map (
            O => \N__21048\,
            I => \N__21037\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__21045\,
            I => \N__21034\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__21040\,
            I => \N__21031\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__21037\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__21034\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__21031\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__4171\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21017\
        );

    \I__4170\ : CascadeMux
    port map (
            O => \N__21020\,
            I => \N__21013\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__21008\
        );

    \I__4168\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21005\
        );

    \I__4167\ : InMux
    port map (
            O => \N__21013\,
            I => \N__21002\
        );

    \I__4166\ : InMux
    port map (
            O => \N__21012\,
            I => \N__20999\
        );

    \I__4165\ : InMux
    port map (
            O => \N__21011\,
            I => \N__20996\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__21008\,
            I => \N__20990\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__20990\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__21002\,
            I => \N__20985\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20985\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__20996\,
            I => \N__20982\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__20995\,
            I => \N__20979\
        );

    \I__4158\ : Span4Mux_v
    port map (
            O => \N__20990\,
            I => \N__20974\
        );

    \I__4157\ : Span4Mux_v
    port map (
            O => \N__20985\,
            I => \N__20971\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__20982\,
            I => \N__20968\
        );

    \I__4155\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20965\
        );

    \I__4154\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20960\
        );

    \I__4153\ : InMux
    port map (
            O => \N__20977\,
            I => \N__20960\
        );

    \I__4152\ : Span4Mux_v
    port map (
            O => \N__20974\,
            I => \N__20957\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__20971\,
            I => \N__20952\
        );

    \I__4150\ : Span4Mux_v
    port map (
            O => \N__20968\,
            I => \N__20952\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__20965\,
            I => \N__20947\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__20960\,
            I => \N__20947\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__20957\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__20952\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__4145\ : Odrv12
    port map (
            O => \N__20947\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__4144\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20937\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__20937\,
            I => \N__20934\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__20934\,
            I => \N__20931\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__20931\,
            I => \N__20928\
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__20928\,
            I => \this_sprites_ram.mem_out_bus5_3\
        );

    \I__4139\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20922\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__20922\,
            I => \N__20919\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__20919\,
            I => \N__20916\
        );

    \I__4136\ : Span4Mux_h
    port map (
            O => \N__20916\,
            I => \N__20913\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__20913\,
            I => \N__20910\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__20910\,
            I => \this_sprites_ram.mem_out_bus1_3\
        );

    \I__4133\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__20904\,
            I => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\
        );

    \I__4131\ : InMux
    port map (
            O => \N__20901\,
            I => \N__20895\
        );

    \I__4130\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20892\
        );

    \I__4129\ : InMux
    port map (
            O => \N__20899\,
            I => \N__20889\
        );

    \I__4128\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20886\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__20895\,
            I => \N__20883\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__20892\,
            I => \N__20880\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20875\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__20886\,
            I => \N__20875\
        );

    \I__4123\ : Odrv12
    port map (
            O => \N__20883\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__20880\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__4121\ : Odrv4
    port map (
            O => \N__20875\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__4120\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20865\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__20865\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__20862\,
            I => \N__20859\
        );

    \I__4117\ : CascadeBuf
    port map (
            O => \N__20859\,
            I => \N__20856\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__20856\,
            I => \N__20853\
        );

    \I__4115\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__20847\,
            I => \N__20843\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__20846\,
            I => \N__20839\
        );

    \I__4111\ : Span4Mux_h
    port map (
            O => \N__20843\,
            I => \N__20834\
        );

    \I__4110\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20831\
        );

    \I__4109\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20826\
        );

    \I__4108\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20826\
        );

    \I__4107\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20823\
        );

    \I__4106\ : Span4Mux_h
    port map (
            O => \N__20834\,
            I => \N__20820\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__20831\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__20826\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__20823\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__20820\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__4101\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20807\
        );

    \I__4100\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20804\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__20807\,
            I => \this_ppu.N_144_4\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__20804\,
            I => \this_ppu.N_144_4\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__20799\,
            I => \N__20795\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__20798\,
            I => \N__20792\
        );

    \I__4095\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20789\
        );

    \I__4094\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20786\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__20789\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__20786\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__4091\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20775\
        );

    \I__4089\ : Sp12to4
    port map (
            O => \N__20775\,
            I => \N__20772\
        );

    \I__4088\ : Odrv12
    port map (
            O => \N__20772\,
            I => \this_ppu.N_144\
        );

    \I__4087\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__20766\,
            I => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\
        );

    \I__4085\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20760\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__4083\ : Span4Mux_v
    port map (
            O => \N__20757\,
            I => \N__20754\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__20754\,
            I => \N__20751\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__20751\,
            I => \N__20748\
        );

    \I__4080\ : Span4Mux_h
    port map (
            O => \N__20748\,
            I => \N__20745\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__20745\,
            I => \M_this_ppu_vram_data_0\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__20742\,
            I => \M_this_ppu_vram_data_0_cascade_\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__20739\,
            I => \this_ppu.N_156_cascade_\
        );

    \I__4076\ : CEMux
    port map (
            O => \N__20736\,
            I => \N__20733\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__20733\,
            I => \N__20730\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__4073\ : Span4Mux_v
    port map (
            O => \N__20727\,
            I => \N__20724\
        );

    \I__4072\ : Span4Mux_h
    port map (
            O => \N__20724\,
            I => \N__20719\
        );

    \I__4071\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20716\
        );

    \I__4070\ : InMux
    port map (
            O => \N__20722\,
            I => \N__20712\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__20719\,
            I => \N__20707\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20707\
        );

    \I__4067\ : InMux
    port map (
            O => \N__20715\,
            I => \N__20704\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__20712\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__20707\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__20704\,
            I => \M_this_ppu_vram_en_0\
        );

    \I__4063\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20694\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__4061\ : Span4Mux_h
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__4060\ : Span4Mux_v
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__20685\,
            I => \N__20682\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__20682\,
            I => \this_sprites_ram.mem_out_bus6_3\
        );

    \I__4057\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__20676\,
            I => \N__20673\
        );

    \I__4055\ : Span12Mux_h
    port map (
            O => \N__20673\,
            I => \N__20670\
        );

    \I__4054\ : Odrv12
    port map (
            O => \N__20670\,
            I => \this_sprites_ram.mem_out_bus2_3\
        );

    \I__4053\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20664\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__4051\ : Span4Mux_v
    port map (
            O => \N__20661\,
            I => \N__20658\
        );

    \I__4050\ : Sp12to4
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__4049\ : Odrv12
    port map (
            O => \N__20655\,
            I => \this_sprites_ram.mem_out_bus4_0\
        );

    \I__4048\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20649\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__20649\,
            I => \N__20646\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__4045\ : Span4Mux_h
    port map (
            O => \N__20643\,
            I => \N__20640\
        );

    \I__4044\ : Span4Mux_v
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__4043\ : Span4Mux_v
    port map (
            O => \N__20637\,
            I => \N__20634\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__20634\,
            I => \this_sprites_ram.mem_out_bus0_0\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__20631\,
            I => \N__20628\
        );

    \I__4040\ : CascadeBuf
    port map (
            O => \N__20628\,
            I => \N__20625\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__20625\,
            I => \N__20622\
        );

    \I__4038\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__20619\,
            I => \N__20615\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__20618\,
            I => \N__20611\
        );

    \I__4035\ : Span4Mux_h
    port map (
            O => \N__20615\,
            I => \N__20608\
        );

    \I__4034\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20605\
        );

    \I__4033\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20602\
        );

    \I__4032\ : Sp12to4
    port map (
            O => \N__20608\,
            I => \N__20599\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__20605\,
            I => \N__20594\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__20602\,
            I => \N__20591\
        );

    \I__4029\ : Span12Mux_v
    port map (
            O => \N__20599\,
            I => \N__20588\
        );

    \I__4028\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20585\
        );

    \I__4027\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20582\
        );

    \I__4026\ : Span12Mux_v
    port map (
            O => \N__20594\,
            I => \N__20575\
        );

    \I__4025\ : Span12Mux_h
    port map (
            O => \N__20591\,
            I => \N__20575\
        );

    \I__4024\ : Span12Mux_h
    port map (
            O => \N__20588\,
            I => \N__20575\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__20585\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__20582\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4021\ : Odrv12
    port map (
            O => \N__20575\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__20568\,
            I => \N__20565\
        );

    \I__4019\ : CascadeBuf
    port map (
            O => \N__20565\,
            I => \N__20562\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__20562\,
            I => \N__20558\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__20561\,
            I => \N__20555\
        );

    \I__4016\ : InMux
    port map (
            O => \N__20558\,
            I => \N__20552\
        );

    \I__4015\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20549\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__20552\,
            I => \N__20546\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__20549\,
            I => \N__20542\
        );

    \I__4012\ : Span4Mux_h
    port map (
            O => \N__20546\,
            I => \N__20539\
        );

    \I__4011\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20536\
        );

    \I__4010\ : Span4Mux_h
    port map (
            O => \N__20542\,
            I => \N__20533\
        );

    \I__4009\ : Span4Mux_v
    port map (
            O => \N__20539\,
            I => \N__20530\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20524\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__20533\,
            I => \N__20521\
        );

    \I__4006\ : Sp12to4
    port map (
            O => \N__20530\,
            I => \N__20518\
        );

    \I__4005\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20515\
        );

    \I__4004\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20512\
        );

    \I__4003\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20509\
        );

    \I__4002\ : Span12Mux_h
    port map (
            O => \N__20524\,
            I => \N__20506\
        );

    \I__4001\ : Sp12to4
    port map (
            O => \N__20521\,
            I => \N__20501\
        );

    \I__4000\ : Span12Mux_v
    port map (
            O => \N__20518\,
            I => \N__20501\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__20515\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__20512\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__20509\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__3996\ : Odrv12
    port map (
            O => \N__20506\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__3995\ : Odrv12
    port map (
            O => \N__20501\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__20490\,
            I => \N__20487\
        );

    \I__3993\ : CascadeBuf
    port map (
            O => \N__20487\,
            I => \N__20484\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__20484\,
            I => \N__20481\
        );

    \I__3991\ : InMux
    port map (
            O => \N__20481\,
            I => \N__20477\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__20480\,
            I => \N__20474\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__20477\,
            I => \N__20471\
        );

    \I__3988\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20468\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__20471\,
            I => \N__20464\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20461\
        );

    \I__3985\ : InMux
    port map (
            O => \N__20467\,
            I => \N__20458\
        );

    \I__3984\ : Sp12to4
    port map (
            O => \N__20464\,
            I => \N__20455\
        );

    \I__3983\ : Span4Mux_v
    port map (
            O => \N__20461\,
            I => \N__20450\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__20458\,
            I => \N__20445\
        );

    \I__3981\ : Span12Mux_h
    port map (
            O => \N__20455\,
            I => \N__20445\
        );

    \I__3980\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20442\
        );

    \I__3979\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20439\
        );

    \I__3978\ : Sp12to4
    port map (
            O => \N__20450\,
            I => \N__20436\
        );

    \I__3977\ : Span12Mux_v
    port map (
            O => \N__20445\,
            I => \N__20433\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__20442\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__20439\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3974\ : Odrv12
    port map (
            O => \N__20436\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3973\ : Odrv12
    port map (
            O => \N__20433\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__20424\,
            I => \N__20421\
        );

    \I__3971\ : CascadeBuf
    port map (
            O => \N__20421\,
            I => \N__20418\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__20418\,
            I => \N__20415\
        );

    \I__3969\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20412\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__20412\,
            I => \N__20408\
        );

    \I__3967\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20405\
        );

    \I__3966\ : Span4Mux_h
    port map (
            O => \N__20408\,
            I => \N__20402\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__20405\,
            I => \N__20398\
        );

    \I__3964\ : Sp12to4
    port map (
            O => \N__20402\,
            I => \N__20395\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__20401\,
            I => \N__20392\
        );

    \I__3962\ : Span4Mux_v
    port map (
            O => \N__20398\,
            I => \N__20389\
        );

    \I__3961\ : Span12Mux_v
    port map (
            O => \N__20395\,
            I => \N__20386\
        );

    \I__3960\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20383\
        );

    \I__3959\ : Span4Mux_v
    port map (
            O => \N__20389\,
            I => \N__20380\
        );

    \I__3958\ : Span12Mux_h
    port map (
            O => \N__20386\,
            I => \N__20377\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__20383\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__20380\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__3955\ : Odrv12
    port map (
            O => \N__20377\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__3954\ : InMux
    port map (
            O => \N__20370\,
            I => \bfn_18_20_0_\
        );

    \I__3953\ : InMux
    port map (
            O => \N__20367\,
            I => \N__20363\
        );

    \I__3952\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20358\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20355\
        );

    \I__3950\ : InMux
    port map (
            O => \N__20362\,
            I => \N__20350\
        );

    \I__3949\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20350\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__20358\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__20355\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__20350\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__20343\,
            I => \N__20340\
        );

    \I__3944\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20337\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__20337\,
            I => \N__20334\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__20334\,
            I => \this_ppu.un1_M_haddress_q_2_4\
        );

    \I__3941\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20328\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__20328\,
            I => \this_ppu.N_148\
        );

    \I__3939\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20320\
        );

    \I__3938\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20316\
        );

    \I__3937\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20313\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__20320\,
            I => \N__20310\
        );

    \I__3935\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20307\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__20316\,
            I => \this_ppu.vscroll8\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__20313\,
            I => \this_ppu.vscroll8\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__20310\,
            I => \this_ppu.vscroll8\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__20307\,
            I => \this_ppu.vscroll8\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__3929\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20292\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__20289\,
            I => \this_ppu.un1_M_haddress_q_2_5\
        );

    \I__3926\ : CascadeMux
    port map (
            O => \N__20286\,
            I => \this_ppu.un1_M_vaddress_q_2_c2_cascade_\
        );

    \I__3925\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20274\
        );

    \I__3924\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20274\
        );

    \I__3923\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20274\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__20274\,
            I => \this_ppu.un1_M_vaddress_q_2_c5\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__20271\,
            I => \N__20268\
        );

    \I__3920\ : CascadeBuf
    port map (
            O => \N__20268\,
            I => \N__20265\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__20265\,
            I => \N__20261\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__20264\,
            I => \N__20258\
        );

    \I__3917\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20255\
        );

    \I__3916\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20252\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__20255\,
            I => \N__20249\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__20252\,
            I => \N__20245\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__20249\,
            I => \N__20242\
        );

    \I__3912\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20239\
        );

    \I__3911\ : Span4Mux_v
    port map (
            O => \N__20245\,
            I => \N__20236\
        );

    \I__3910\ : Sp12to4
    port map (
            O => \N__20242\,
            I => \N__20233\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__20239\,
            I => \N__20227\
        );

    \I__3908\ : Sp12to4
    port map (
            O => \N__20236\,
            I => \N__20224\
        );

    \I__3907\ : Span12Mux_v
    port map (
            O => \N__20233\,
            I => \N__20221\
        );

    \I__3906\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20216\
        );

    \I__3905\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20216\
        );

    \I__3904\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20213\
        );

    \I__3903\ : Span12Mux_v
    port map (
            O => \N__20227\,
            I => \N__20206\
        );

    \I__3902\ : Span12Mux_h
    port map (
            O => \N__20224\,
            I => \N__20206\
        );

    \I__3901\ : Span12Mux_h
    port map (
            O => \N__20221\,
            I => \N__20206\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__20216\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__20213\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__3898\ : Odrv12
    port map (
            O => \N__20206\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__3897\ : InMux
    port map (
            O => \N__20199\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__3896\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__20190\,
            I => \M_this_data_count_q_cry_7_THRU_CO\
        );

    \I__3893\ : InMux
    port map (
            O => \N__20187\,
            I => \bfn_18_16_0_\
        );

    \I__3892\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__20178\,
            I => \M_this_data_count_q_cry_8_THRU_CO\
        );

    \I__3889\ : InMux
    port map (
            O => \N__20175\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__3888\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20168\
        );

    \I__3887\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20165\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__20168\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__20165\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__3884\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20157\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__20157\,
            I => \M_this_data_count_q_s_10\
        );

    \I__3882\ : InMux
    port map (
            O => \N__20154\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__3880\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20144\
        );

    \I__3879\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20140\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20137\
        );

    \I__3877\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20134\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__20140\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3875\ : Odrv12
    port map (
            O => \N__20137\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__20134\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__3873\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20124\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__20121\,
            I => \M_this_data_count_q_cry_10_THRU_CO\
        );

    \I__3870\ : InMux
    port map (
            O => \N__20118\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__3869\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20110\
        );

    \I__3868\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20105\
        );

    \I__3867\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20105\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__20110\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__20105\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__3864\ : SRMux
    port map (
            O => \N__20100\,
            I => \N__20093\
        );

    \I__3863\ : SRMux
    port map (
            O => \N__20099\,
            I => \N__20088\
        );

    \I__3862\ : SRMux
    port map (
            O => \N__20098\,
            I => \N__20077\
        );

    \I__3861\ : SRMux
    port map (
            O => \N__20097\,
            I => \N__20072\
        );

    \I__3860\ : SRMux
    port map (
            O => \N__20096\,
            I => \N__20069\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__20093\,
            I => \N__20064\
        );

    \I__3858\ : SRMux
    port map (
            O => \N__20092\,
            I => \N__20061\
        );

    \I__3857\ : SRMux
    port map (
            O => \N__20091\,
            I => \N__20058\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__20088\,
            I => \N__20053\
        );

    \I__3855\ : SRMux
    port map (
            O => \N__20087\,
            I => \N__20050\
        );

    \I__3854\ : SRMux
    port map (
            O => \N__20086\,
            I => \N__20047\
        );

    \I__3853\ : SRMux
    port map (
            O => \N__20085\,
            I => \N__20043\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__20084\,
            I => \N__20038\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__20083\,
            I => \N__20035\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__20082\,
            I => \N__20031\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__20081\,
            I => \N__20027\
        );

    \I__3848\ : SRMux
    port map (
            O => \N__20080\,
            I => \N__20024\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__20077\,
            I => \N__20020\
        );

    \I__3846\ : SRMux
    port map (
            O => \N__20076\,
            I => \N__20017\
        );

    \I__3845\ : SRMux
    port map (
            O => \N__20075\,
            I => \N__20014\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__20072\,
            I => \N__20007\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__20069\,
            I => \N__20007\
        );

    \I__3842\ : SRMux
    port map (
            O => \N__20068\,
            I => \N__20004\
        );

    \I__3841\ : SRMux
    port map (
            O => \N__20067\,
            I => \N__20001\
        );

    \I__3840\ : Span4Mux_s2_v
    port map (
            O => \N__20064\,
            I => \N__19994\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__20061\,
            I => \N__19994\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__20058\,
            I => \N__19994\
        );

    \I__3837\ : SRMux
    port map (
            O => \N__20057\,
            I => \N__19991\
        );

    \I__3836\ : SRMux
    port map (
            O => \N__20056\,
            I => \N__19988\
        );

    \I__3835\ : Span4Mux_v
    port map (
            O => \N__20053\,
            I => \N__19979\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__20050\,
            I => \N__19979\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__20047\,
            I => \N__19979\
        );

    \I__3832\ : SRMux
    port map (
            O => \N__20046\,
            I => \N__19976\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__19972\
        );

    \I__3830\ : SRMux
    port map (
            O => \N__20042\,
            I => \N__19969\
        );

    \I__3829\ : IoInMux
    port map (
            O => \N__20041\,
            I => \N__19965\
        );

    \I__3828\ : InMux
    port map (
            O => \N__20038\,
            I => \N__19957\
        );

    \I__3827\ : InMux
    port map (
            O => \N__20035\,
            I => \N__19957\
        );

    \I__3826\ : InMux
    port map (
            O => \N__20034\,
            I => \N__19957\
        );

    \I__3825\ : InMux
    port map (
            O => \N__20031\,
            I => \N__19950\
        );

    \I__3824\ : InMux
    port map (
            O => \N__20030\,
            I => \N__19950\
        );

    \I__3823\ : InMux
    port map (
            O => \N__20027\,
            I => \N__19950\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__20024\,
            I => \N__19947\
        );

    \I__3821\ : SRMux
    port map (
            O => \N__20023\,
            I => \N__19944\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__20020\,
            I => \N__19937\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__20017\,
            I => \N__19937\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__19937\
        );

    \I__3817\ : SRMux
    port map (
            O => \N__20013\,
            I => \N__19934\
        );

    \I__3816\ : SRMux
    port map (
            O => \N__20012\,
            I => \N__19931\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__20007\,
            I => \N__19924\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__19924\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__20001\,
            I => \N__19924\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__19994\,
            I => \N__19917\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__19991\,
            I => \N__19917\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19917\
        );

    \I__3809\ : SRMux
    port map (
            O => \N__19987\,
            I => \N__19914\
        );

    \I__3808\ : SRMux
    port map (
            O => \N__19986\,
            I => \N__19907\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__19979\,
            I => \N__19902\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__19976\,
            I => \N__19902\
        );

    \I__3805\ : SRMux
    port map (
            O => \N__19975\,
            I => \N__19899\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__19972\,
            I => \N__19894\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__19969\,
            I => \N__19894\
        );

    \I__3802\ : SRMux
    port map (
            O => \N__19968\,
            I => \N__19891\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__19965\,
            I => \N__19888\
        );

    \I__3800\ : SRMux
    port map (
            O => \N__19964\,
            I => \N__19884\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__19957\,
            I => \N__19879\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__19950\,
            I => \N__19879\
        );

    \I__3797\ : Span4Mux_h
    port map (
            O => \N__19947\,
            I => \N__19874\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__19944\,
            I => \N__19871\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__19937\,
            I => \N__19866\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19866\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__19931\,
            I => \N__19862\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__19924\,
            I => \N__19859\
        );

    \I__3791\ : Span4Mux_v
    port map (
            O => \N__19917\,
            I => \N__19854\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__19914\,
            I => \N__19854\
        );

    \I__3789\ : SRMux
    port map (
            O => \N__19913\,
            I => \N__19851\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__19912\,
            I => \N__19846\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__19911\,
            I => \N__19842\
        );

    \I__3786\ : CascadeMux
    port map (
            O => \N__19910\,
            I => \N__19838\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19828\
        );

    \I__3784\ : Span4Mux_h
    port map (
            O => \N__19902\,
            I => \N__19828\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__19899\,
            I => \N__19828\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__19894\,
            I => \N__19823\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19823\
        );

    \I__3780\ : IoSpan4Mux
    port map (
            O => \N__19888\,
            I => \N__19819\
        );

    \I__3779\ : SRMux
    port map (
            O => \N__19887\,
            I => \N__19816\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__19884\,
            I => \N__19813\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__19879\,
            I => \N__19810\
        );

    \I__3776\ : SRMux
    port map (
            O => \N__19878\,
            I => \N__19806\
        );

    \I__3775\ : SRMux
    port map (
            O => \N__19877\,
            I => \N__19803\
        );

    \I__3774\ : Span4Mux_v
    port map (
            O => \N__19874\,
            I => \N__19797\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__19871\,
            I => \N__19797\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__19866\,
            I => \N__19794\
        );

    \I__3771\ : SRMux
    port map (
            O => \N__19865\,
            I => \N__19791\
        );

    \I__3770\ : Span4Mux_s2_v
    port map (
            O => \N__19862\,
            I => \N__19788\
        );

    \I__3769\ : Span4Mux_v
    port map (
            O => \N__19859\,
            I => \N__19781\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__19854\,
            I => \N__19781\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19781\
        );

    \I__3766\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19766\
        );

    \I__3765\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19766\
        );

    \I__3764\ : InMux
    port map (
            O => \N__19846\,
            I => \N__19766\
        );

    \I__3763\ : InMux
    port map (
            O => \N__19845\,
            I => \N__19766\
        );

    \I__3762\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19766\
        );

    \I__3761\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19766\
        );

    \I__3760\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19766\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__19837\,
            I => \N__19762\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__19836\,
            I => \N__19759\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__19835\,
            I => \N__19755\
        );

    \I__3756\ : Span4Mux_v
    port map (
            O => \N__19828\,
            I => \N__19750\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__19823\,
            I => \N__19750\
        );

    \I__3754\ : SRMux
    port map (
            O => \N__19822\,
            I => \N__19747\
        );

    \I__3753\ : Span4Mux_s2_h
    port map (
            O => \N__19819\,
            I => \N__19741\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__19816\,
            I => \N__19738\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__19813\,
            I => \N__19733\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__19810\,
            I => \N__19733\
        );

    \I__3749\ : SRMux
    port map (
            O => \N__19809\,
            I => \N__19730\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__19806\,
            I => \N__19724\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19724\
        );

    \I__3746\ : SRMux
    port map (
            O => \N__19802\,
            I => \N__19721\
        );

    \I__3745\ : Span4Mux_v
    port map (
            O => \N__19797\,
            I => \N__19714\
        );

    \I__3744\ : Span4Mux_v
    port map (
            O => \N__19794\,
            I => \N__19714\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__19791\,
            I => \N__19714\
        );

    \I__3742\ : Span4Mux_h
    port map (
            O => \N__19788\,
            I => \N__19711\
        );

    \I__3741\ : Span4Mux_h
    port map (
            O => \N__19781\,
            I => \N__19706\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__19766\,
            I => \N__19706\
        );

    \I__3739\ : InMux
    port map (
            O => \N__19765\,
            I => \N__19695\
        );

    \I__3738\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19695\
        );

    \I__3737\ : InMux
    port map (
            O => \N__19759\,
            I => \N__19695\
        );

    \I__3736\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19695\
        );

    \I__3735\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19695\
        );

    \I__3734\ : Span4Mux_v
    port map (
            O => \N__19750\,
            I => \N__19690\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__19747\,
            I => \N__19690\
        );

    \I__3732\ : SRMux
    port map (
            O => \N__19746\,
            I => \N__19687\
        );

    \I__3731\ : SRMux
    port map (
            O => \N__19745\,
            I => \N__19684\
        );

    \I__3730\ : SRMux
    port map (
            O => \N__19744\,
            I => \N__19681\
        );

    \I__3729\ : Sp12to4
    port map (
            O => \N__19741\,
            I => \N__19676\
        );

    \I__3728\ : Sp12to4
    port map (
            O => \N__19738\,
            I => \N__19676\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__19733\,
            I => \N__19671\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19671\
        );

    \I__3725\ : IoInMux
    port map (
            O => \N__19729\,
            I => \N__19668\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__19724\,
            I => \N__19662\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__19721\,
            I => \N__19662\
        );

    \I__3722\ : Span4Mux_h
    port map (
            O => \N__19714\,
            I => \N__19659\
        );

    \I__3721\ : Sp12to4
    port map (
            O => \N__19711\,
            I => \N__19655\
        );

    \I__3720\ : Span4Mux_h
    port map (
            O => \N__19706\,
            I => \N__19650\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__19695\,
            I => \N__19650\
        );

    \I__3718\ : Span4Mux_h
    port map (
            O => \N__19690\,
            I => \N__19647\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19642\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19642\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19639\
        );

    \I__3714\ : Span12Mux_h
    port map (
            O => \N__19676\,
            I => \N__19636\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__19671\,
            I => \N__19633\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__19668\,
            I => \N__19630\
        );

    \I__3711\ : SRMux
    port map (
            O => \N__19667\,
            I => \N__19627\
        );

    \I__3710\ : Span4Mux_v
    port map (
            O => \N__19662\,
            I => \N__19624\
        );

    \I__3709\ : Span4Mux_v
    port map (
            O => \N__19659\,
            I => \N__19621\
        );

    \I__3708\ : SRMux
    port map (
            O => \N__19658\,
            I => \N__19618\
        );

    \I__3707\ : Span12Mux_v
    port map (
            O => \N__19655\,
            I => \N__19614\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__19650\,
            I => \N__19611\
        );

    \I__3705\ : Span4Mux_v
    port map (
            O => \N__19647\,
            I => \N__19606\
        );

    \I__3704\ : Span4Mux_v
    port map (
            O => \N__19642\,
            I => \N__19606\
        );

    \I__3703\ : Span4Mux_v
    port map (
            O => \N__19639\,
            I => \N__19603\
        );

    \I__3702\ : Span12Mux_h
    port map (
            O => \N__19636\,
            I => \N__19598\
        );

    \I__3701\ : Sp12to4
    port map (
            O => \N__19633\,
            I => \N__19598\
        );

    \I__3700\ : IoSpan4Mux
    port map (
            O => \N__19630\,
            I => \N__19595\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__19627\,
            I => \N__19592\
        );

    \I__3698\ : Span4Mux_v
    port map (
            O => \N__19624\,
            I => \N__19585\
        );

    \I__3697\ : Span4Mux_v
    port map (
            O => \N__19621\,
            I => \N__19585\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__19618\,
            I => \N__19585\
        );

    \I__3695\ : SRMux
    port map (
            O => \N__19617\,
            I => \N__19582\
        );

    \I__3694\ : Span12Mux_h
    port map (
            O => \N__19614\,
            I => \N__19578\
        );

    \I__3693\ : Sp12to4
    port map (
            O => \N__19611\,
            I => \N__19575\
        );

    \I__3692\ : Sp12to4
    port map (
            O => \N__19606\,
            I => \N__19570\
        );

    \I__3691\ : Sp12to4
    port map (
            O => \N__19603\,
            I => \N__19570\
        );

    \I__3690\ : Span12Mux_v
    port map (
            O => \N__19598\,
            I => \N__19567\
        );

    \I__3689\ : IoSpan4Mux
    port map (
            O => \N__19595\,
            I => \N__19564\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__19592\,
            I => \N__19557\
        );

    \I__3687\ : Span4Mux_v
    port map (
            O => \N__19585\,
            I => \N__19557\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__19582\,
            I => \N__19557\
        );

    \I__3685\ : SRMux
    port map (
            O => \N__19581\,
            I => \N__19554\
        );

    \I__3684\ : Span12Mux_v
    port map (
            O => \N__19578\,
            I => \N__19551\
        );

    \I__3683\ : Span12Mux_h
    port map (
            O => \N__19575\,
            I => \N__19548\
        );

    \I__3682\ : Span12Mux_h
    port map (
            O => \N__19570\,
            I => \N__19543\
        );

    \I__3681\ : Span12Mux_v
    port map (
            O => \N__19567\,
            I => \N__19543\
        );

    \I__3680\ : Span4Mux_s2_h
    port map (
            O => \N__19564\,
            I => \N__19540\
        );

    \I__3679\ : Span4Mux_v
    port map (
            O => \N__19557\,
            I => \N__19535\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__19554\,
            I => \N__19535\
        );

    \I__3677\ : Odrv12
    port map (
            O => \N__19551\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3676\ : Odrv12
    port map (
            O => \N__19548\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3675\ : Odrv12
    port map (
            O => \N__19543\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__19540\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__19535\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3672\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19521\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__19521\,
            I => \M_this_data_count_q_cry_11_THRU_CO\
        );

    \I__3670\ : InMux
    port map (
            O => \N__19518\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__3669\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19511\
        );

    \I__3668\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \N__19508\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__19511\,
            I => \N__19505\
        );

    \I__3666\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19502\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__19505\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__19502\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__3663\ : InMux
    port map (
            O => \N__19497\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__3662\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19491\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19488\
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__19488\,
            I => \M_this_data_count_q_s_13\
        );

    \I__3659\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19482\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__19482\,
            I => \N_49\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__3656\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19473\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__19473\,
            I => \N__19470\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__19470\,
            I => \N__19467\
        );

    \I__3653\ : Span4Mux_h
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__19464\,
            I => this_vga_signals_vvisibility_1
        );

    \I__3651\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__19458\,
            I => \N__19443\
        );

    \I__3649\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19440\
        );

    \I__3648\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19437\
        );

    \I__3647\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19428\
        );

    \I__3646\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19428\
        );

    \I__3645\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19428\
        );

    \I__3644\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19428\
        );

    \I__3643\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19417\
        );

    \I__3642\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19417\
        );

    \I__3641\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19417\
        );

    \I__3640\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19417\
        );

    \I__3639\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19417\
        );

    \I__3638\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19414\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__19443\,
            I => \N_686_i\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__19440\,
            I => \N_686_i\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__19437\,
            I => \N_686_i\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__19428\,
            I => \N_686_i\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__19417\,
            I => \N_686_i\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__19414\,
            I => \N_686_i\
        );

    \I__3631\ : CEMux
    port map (
            O => \N__19401\,
            I => \N__19398\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__19398\,
            I => \N__19390\
        );

    \I__3629\ : CEMux
    port map (
            O => \N__19397\,
            I => \N__19387\
        );

    \I__3628\ : CEMux
    port map (
            O => \N__19396\,
            I => \N__19384\
        );

    \I__3627\ : CEMux
    port map (
            O => \N__19395\,
            I => \N__19381\
        );

    \I__3626\ : CEMux
    port map (
            O => \N__19394\,
            I => \N__19378\
        );

    \I__3625\ : CEMux
    port map (
            O => \N__19393\,
            I => \N__19375\
        );

    \I__3624\ : Odrv12
    port map (
            O => \N__19390\,
            I => \M_this_data_count_qlde_i_i\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__19387\,
            I => \M_this_data_count_qlde_i_i\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__19384\,
            I => \M_this_data_count_qlde_i_i\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__19381\,
            I => \M_this_data_count_qlde_i_i\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__19378\,
            I => \M_this_data_count_qlde_i_i\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__19375\,
            I => \M_this_data_count_qlde_i_i\
        );

    \I__3618\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19357\
        );

    \I__3617\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19352\
        );

    \I__3616\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19352\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__19357\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__19352\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__3612\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19339\
        );

    \I__3611\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19334\
        );

    \I__3610\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19334\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__19339\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__19334\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__3607\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__19326\,
            I => \M_this_data_count_q_cry_0_THRU_CO\
        );

    \I__3605\ : InMux
    port map (
            O => \N__19323\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__3604\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__19317\,
            I => \N__19312\
        );

    \I__3602\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19309\
        );

    \I__3601\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19306\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__19312\,
            I => \N__19303\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__19309\,
            I => \N__19300\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__19306\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__19303\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__19300\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__3595\ : InMux
    port map (
            O => \N__19293\,
            I => \N__19290\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__19290\,
            I => \N__19287\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__19287\,
            I => \N__19284\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__19284\,
            I => \M_this_data_count_q_cry_1_THRU_CO\
        );

    \I__3591\ : InMux
    port map (
            O => \N__19281\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__3589\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19272\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__19272\,
            I => \N__19267\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__19271\,
            I => \N__19264\
        );

    \I__3586\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19261\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__19267\,
            I => \N__19258\
        );

    \I__3584\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19255\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__19261\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__19258\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__19255\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__3580\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__19242\,
            I => \M_this_data_count_q_cry_2_THRU_CO\
        );

    \I__3577\ : InMux
    port map (
            O => \N__19239\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__3576\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__19233\,
            I => \M_this_data_count_q_cry_3_THRU_CO\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19230\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__3573\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__3571\ : Span4Mux_h
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__3570\ : Odrv4
    port map (
            O => \N__19218\,
            I => \M_this_data_count_q_cry_4_THRU_CO\
        );

    \I__3569\ : InMux
    port map (
            O => \N__19215\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__3568\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19208\
        );

    \I__3567\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19205\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__19208\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__19205\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__3564\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__19197\,
            I => \M_this_data_count_q_s_6\
        );

    \I__3562\ : InMux
    port map (
            O => \N__19194\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__19191\,
            I => \N__19188\
        );

    \I__3560\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__19185\,
            I => \N__19180\
        );

    \I__3558\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19175\
        );

    \I__3557\ : InMux
    port map (
            O => \N__19183\,
            I => \N__19175\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__19180\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__19175\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__3554\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19167\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__19167\,
            I => \M_this_data_count_q_cry_6_THRU_CO\
        );

    \I__3552\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19158\
        );

    \I__3551\ : InMux
    port map (
            O => \N__19163\,
            I => \N__19158\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__19158\,
            I => \this_ppu.un1_M_haddress_q_3_c2\
        );

    \I__3549\ : SRMux
    port map (
            O => \N__19155\,
            I => \N__19151\
        );

    \I__3548\ : SRMux
    port map (
            O => \N__19154\,
            I => \N__19148\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19145\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19142\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__19145\,
            I => \N__19134\
        );

    \I__3544\ : Span4Mux_v
    port map (
            O => \N__19142\,
            I => \N__19134\
        );

    \I__3543\ : SRMux
    port map (
            O => \N__19141\,
            I => \N__19131\
        );

    \I__3542\ : SRMux
    port map (
            O => \N__19140\,
            I => \N__19128\
        );

    \I__3541\ : SRMux
    port map (
            O => \N__19139\,
            I => \N__19125\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__19134\,
            I => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__19131\,
            I => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__19128\,
            I => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__19125\,
            I => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\
        );

    \I__3536\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19113\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__19113\,
            I => \N__19110\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__19110\,
            I => \N__19107\
        );

    \I__3533\ : Sp12to4
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__3532\ : Odrv12
    port map (
            O => \N__19104\,
            I => \this_sprites_ram.mem_out_bus4_3\
        );

    \I__3531\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19098\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__19098\,
            I => \N__19095\
        );

    \I__3529\ : Span4Mux_v
    port map (
            O => \N__19095\,
            I => \N__19092\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__19092\,
            I => \N__19089\
        );

    \I__3527\ : Span4Mux_h
    port map (
            O => \N__19089\,
            I => \N__19086\
        );

    \I__3526\ : Span4Mux_v
    port map (
            O => \N__19086\,
            I => \N__19083\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__19083\,
            I => \this_sprites_ram.mem_out_bus0_3\
        );

    \I__3524\ : CEMux
    port map (
            O => \N__19080\,
            I => \N__19077\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__19077\,
            I => \N__19073\
        );

    \I__3522\ : CEMux
    port map (
            O => \N__19076\,
            I => \N__19070\
        );

    \I__3521\ : Span4Mux_v
    port map (
            O => \N__19073\,
            I => \N__19065\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__19070\,
            I => \N__19065\
        );

    \I__3519\ : Span4Mux_h
    port map (
            O => \N__19065\,
            I => \N__19062\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__19062\,
            I => \N__19059\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__19059\,
            I => \this_sprites_ram.mem_WE_8\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__19056\,
            I => \N__19053\
        );

    \I__3515\ : CascadeBuf
    port map (
            O => \N__19053\,
            I => \N__19050\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__19050\,
            I => \N__19047\
        );

    \I__3513\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19042\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19039\
        );

    \I__3511\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19035\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__19042\,
            I => \N__19032\
        );

    \I__3509\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19029\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19026\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__19035\,
            I => \N__19023\
        );

    \I__3506\ : Span12Mux_v
    port map (
            O => \N__19032\,
            I => \N__19020\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__19029\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__19026\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__19023\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__3502\ : Odrv12
    port map (
            O => \N__19020\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__19011\,
            I => \N__19008\
        );

    \I__3500\ : CascadeBuf
    port map (
            O => \N__19008\,
            I => \N__19005\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__19005\,
            I => \N__19002\
        );

    \I__3498\ : InMux
    port map (
            O => \N__19002\,
            I => \N__18999\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__18999\,
            I => \N__18996\
        );

    \I__3496\ : Sp12to4
    port map (
            O => \N__18996\,
            I => \N__18989\
        );

    \I__3495\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18982\
        );

    \I__3494\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18982\
        );

    \I__3493\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18982\
        );

    \I__3492\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18979\
        );

    \I__3491\ : Span12Mux_v
    port map (
            O => \N__18989\,
            I => \N__18976\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__18982\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__18979\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__3488\ : Odrv12
    port map (
            O => \N__18976\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__18969\,
            I => \N__18965\
        );

    \I__3486\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18962\
        );

    \I__3485\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18959\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__18962\,
            I => \this_ppu.M_oam_idx_qZ0Z_4\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__18959\,
            I => \this_ppu.M_oam_idx_qZ0Z_4\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__18954\,
            I => \N__18951\
        );

    \I__3481\ : CascadeBuf
    port map (
            O => \N__18951\,
            I => \N__18948\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__3479\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18942\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__18942\,
            I => \N__18938\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \N__18934\
        );

    \I__3476\ : Span4Mux_v
    port map (
            O => \N__18938\,
            I => \N__18930\
        );

    \I__3475\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18927\
        );

    \I__3474\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18922\
        );

    \I__3473\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18922\
        );

    \I__3472\ : Span4Mux_h
    port map (
            O => \N__18930\,
            I => \N__18919\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__18927\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__18922\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__18919\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__18912\,
            I => \this_ppu.un1_M_haddress_q_3_c2_cascade_\
        );

    \I__3467\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18904\
        );

    \I__3466\ : InMux
    port map (
            O => \N__18908\,
            I => \N__18901\
        );

    \I__3465\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18898\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__18904\,
            I => \this_ppu.un1_M_haddress_q_3_c5\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__18901\,
            I => \this_ppu.un1_M_haddress_q_3_c5\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__18898\,
            I => \this_ppu.un1_M_haddress_q_3_c5\
        );

    \I__3461\ : InMux
    port map (
            O => \N__18891\,
            I => \N__18888\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__18888\,
            I => \N__18885\
        );

    \I__3459\ : Span4Mux_h
    port map (
            O => \N__18885\,
            I => \N__18882\
        );

    \I__3458\ : Span4Mux_h
    port map (
            O => \N__18882\,
            I => \N__18879\
        );

    \I__3457\ : Sp12to4
    port map (
            O => \N__18879\,
            I => \N__18876\
        );

    \I__3456\ : Odrv12
    port map (
            O => \N__18876\,
            I => \this_sprites_ram.mem_out_bus7_0\
        );

    \I__3455\ : InMux
    port map (
            O => \N__18873\,
            I => \N__18870\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__18870\,
            I => \N__18867\
        );

    \I__3453\ : Span12Mux_h
    port map (
            O => \N__18867\,
            I => \N__18864\
        );

    \I__3452\ : Odrv12
    port map (
            O => \N__18864\,
            I => \this_sprites_ram.mem_out_bus3_0\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__18861\,
            I => \this_ppu.un2_hscroll_axb_0_cascade_\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__18858\,
            I => \N__18855\
        );

    \I__3449\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18848\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__18854\,
            I => \N__18845\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__18853\,
            I => \N__18840\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__18852\,
            I => \N__18837\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__18851\,
            I => \N__18834\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__18848\,
            I => \N__18826\
        );

    \I__3443\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18823\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__18844\,
            I => \N__18820\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__18843\,
            I => \N__18817\
        );

    \I__3440\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18813\
        );

    \I__3439\ : InMux
    port map (
            O => \N__18837\,
            I => \N__18810\
        );

    \I__3438\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18807\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__18833\,
            I => \N__18804\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__18832\,
            I => \N__18800\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__18831\,
            I => \N__18797\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__18830\,
            I => \N__18794\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__18829\,
            I => \N__18791\
        );

    \I__3432\ : Span4Mux_s0_v
    port map (
            O => \N__18826\,
            I => \N__18784\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18784\
        );

    \I__3430\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18781\
        );

    \I__3429\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18778\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__18816\,
            I => \N__18775\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__18813\,
            I => \N__18770\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__18810\,
            I => \N__18770\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__18807\,
            I => \N__18767\
        );

    \I__3424\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18764\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__18803\,
            I => \N__18761\
        );

    \I__3422\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18758\
        );

    \I__3421\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18755\
        );

    \I__3420\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18752\
        );

    \I__3419\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18749\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__18790\,
            I => \N__18746\
        );

    \I__3417\ : CascadeMux
    port map (
            O => \N__18789\,
            I => \N__18743\
        );

    \I__3416\ : Span4Mux_v
    port map (
            O => \N__18784\,
            I => \N__18738\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__18781\,
            I => \N__18738\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__18778\,
            I => \N__18735\
        );

    \I__3413\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18732\
        );

    \I__3412\ : Span4Mux_v
    port map (
            O => \N__18770\,
            I => \N__18725\
        );

    \I__3411\ : Span4Mux_h
    port map (
            O => \N__18767\,
            I => \N__18725\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__18764\,
            I => \N__18725\
        );

    \I__3409\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18722\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__18758\,
            I => \N__18719\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__18755\,
            I => \N__18716\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18711\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__18749\,
            I => \N__18711\
        );

    \I__3404\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18708\
        );

    \I__3403\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18705\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__18738\,
            I => \N__18702\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__18735\,
            I => \N__18697\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__18732\,
            I => \N__18697\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__18725\,
            I => \N__18692\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__18722\,
            I => \N__18692\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__18719\,
            I => \N__18689\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__18716\,
            I => \N__18682\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__18711\,
            I => \N__18682\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__18708\,
            I => \N__18682\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__18705\,
            I => \N__18679\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__18702\,
            I => \N__18674\
        );

    \I__3391\ : Span4Mux_h
    port map (
            O => \N__18697\,
            I => \N__18674\
        );

    \I__3390\ : Span4Mux_h
    port map (
            O => \N__18692\,
            I => \N__18671\
        );

    \I__3389\ : Span4Mux_v
    port map (
            O => \N__18689\,
            I => \N__18666\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__18682\,
            I => \N__18666\
        );

    \I__3387\ : Span4Mux_h
    port map (
            O => \N__18679\,
            I => \N__18663\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__18674\,
            I => \N__18658\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__18671\,
            I => \N__18658\
        );

    \I__3384\ : Span4Mux_h
    port map (
            O => \N__18666\,
            I => \N__18653\
        );

    \I__3383\ : Span4Mux_h
    port map (
            O => \N__18663\,
            I => \N__18653\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__18658\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__18653\,
            I => \M_this_ppu_sprites_addr_0\
        );

    \I__3380\ : IoInMux
    port map (
            O => \N__18648\,
            I => \N__18644\
        );

    \I__3379\ : IoInMux
    port map (
            O => \N__18647\,
            I => \N__18637\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__18644\,
            I => \N__18633\
        );

    \I__3377\ : IoInMux
    port map (
            O => \N__18643\,
            I => \N__18630\
        );

    \I__3376\ : IoInMux
    port map (
            O => \N__18642\,
            I => \N__18627\
        );

    \I__3375\ : IoInMux
    port map (
            O => \N__18641\,
            I => \N__18623\
        );

    \I__3374\ : IoInMux
    port map (
            O => \N__18640\,
            I => \N__18620\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18617\
        );

    \I__3372\ : IoInMux
    port map (
            O => \N__18636\,
            I => \N__18614\
        );

    \I__3371\ : IoSpan4Mux
    port map (
            O => \N__18633\,
            I => \N__18604\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__18630\,
            I => \N__18604\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__18627\,
            I => \N__18601\
        );

    \I__3368\ : IoInMux
    port map (
            O => \N__18626\,
            I => \N__18598\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__18623\,
            I => \N__18591\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__18620\,
            I => \N__18591\
        );

    \I__3365\ : IoSpan4Mux
    port map (
            O => \N__18617\,
            I => \N__18585\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__18614\,
            I => \N__18585\
        );

    \I__3363\ : IoInMux
    port map (
            O => \N__18613\,
            I => \N__18582\
        );

    \I__3362\ : IoInMux
    port map (
            O => \N__18612\,
            I => \N__18579\
        );

    \I__3361\ : IoInMux
    port map (
            O => \N__18611\,
            I => \N__18576\
        );

    \I__3360\ : IoInMux
    port map (
            O => \N__18610\,
            I => \N__18573\
        );

    \I__3359\ : IoInMux
    port map (
            O => \N__18609\,
            I => \N__18570\
        );

    \I__3358\ : IoSpan4Mux
    port map (
            O => \N__18604\,
            I => \N__18563\
        );

    \I__3357\ : IoSpan4Mux
    port map (
            O => \N__18601\,
            I => \N__18563\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__18598\,
            I => \N__18563\
        );

    \I__3355\ : IoInMux
    port map (
            O => \N__18597\,
            I => \N__18560\
        );

    \I__3354\ : IoInMux
    port map (
            O => \N__18596\,
            I => \N__18557\
        );

    \I__3353\ : IoSpan4Mux
    port map (
            O => \N__18591\,
            I => \N__18553\
        );

    \I__3352\ : IoInMux
    port map (
            O => \N__18590\,
            I => \N__18550\
        );

    \I__3351\ : IoSpan4Mux
    port map (
            O => \N__18585\,
            I => \N__18541\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__18582\,
            I => \N__18541\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__18579\,
            I => \N__18541\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__18576\,
            I => \N__18541\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18536\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__18570\,
            I => \N__18536\
        );

    \I__3345\ : IoSpan4Mux
    port map (
            O => \N__18563\,
            I => \N__18531\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__18560\,
            I => \N__18531\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__18557\,
            I => \N__18528\
        );

    \I__3342\ : IoInMux
    port map (
            O => \N__18556\,
            I => \N__18525\
        );

    \I__3341\ : Sp12to4
    port map (
            O => \N__18553\,
            I => \N__18522\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18519\
        );

    \I__3339\ : IoSpan4Mux
    port map (
            O => \N__18541\,
            I => \N__18514\
        );

    \I__3338\ : IoSpan4Mux
    port map (
            O => \N__18536\,
            I => \N__18514\
        );

    \I__3337\ : IoSpan4Mux
    port map (
            O => \N__18531\,
            I => \N__18509\
        );

    \I__3336\ : IoSpan4Mux
    port map (
            O => \N__18528\,
            I => \N__18509\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__18525\,
            I => \N__18506\
        );

    \I__3334\ : Span12Mux_s1_h
    port map (
            O => \N__18522\,
            I => \N__18503\
        );

    \I__3333\ : IoSpan4Mux
    port map (
            O => \N__18519\,
            I => \N__18500\
        );

    \I__3332\ : Span4Mux_s0_h
    port map (
            O => \N__18514\,
            I => \N__18497\
        );

    \I__3331\ : Span4Mux_s2_v
    port map (
            O => \N__18509\,
            I => \N__18492\
        );

    \I__3330\ : Span4Mux_s2_v
    port map (
            O => \N__18506\,
            I => \N__18492\
        );

    \I__3329\ : Span12Mux_h
    port map (
            O => \N__18503\,
            I => \N__18489\
        );

    \I__3328\ : Sp12to4
    port map (
            O => \N__18500\,
            I => \N__18486\
        );

    \I__3327\ : Span4Mux_h
    port map (
            O => \N__18497\,
            I => \N__18483\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__18492\,
            I => \N__18480\
        );

    \I__3325\ : Span12Mux_v
    port map (
            O => \N__18489\,
            I => \N__18475\
        );

    \I__3324\ : Span12Mux_s6_h
    port map (
            O => \N__18486\,
            I => \N__18475\
        );

    \I__3323\ : Sp12to4
    port map (
            O => \N__18483\,
            I => \N__18472\
        );

    \I__3322\ : Span4Mux_v
    port map (
            O => \N__18480\,
            I => \N__18469\
        );

    \I__3321\ : Odrv12
    port map (
            O => \N__18475\,
            I => port_dmab_c_i
        );

    \I__3320\ : Odrv12
    port map (
            O => \N__18472\,
            I => port_dmab_c_i
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__18469\,
            I => port_dmab_c_i
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__18462\,
            I => \this_ppu.un1_M_oam_idx_q_1_c1_cascade_\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__18459\,
            I => \this_ppu.un1_M_oam_idx_q_1_c3_cascade_\
        );

    \I__3316\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18452\
        );

    \I__3315\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18449\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__18452\,
            I => \N__18443\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__18449\,
            I => \N__18443\
        );

    \I__3312\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18439\
        );

    \I__3311\ : Span12Mux_v
    port map (
            O => \N__18443\,
            I => \N__18436\
        );

    \I__3310\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18433\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__18439\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_7\
        );

    \I__3308\ : Odrv12
    port map (
            O => \N__18436\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_7\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__18433\,
            I => \this_ppu.M_count_d_0_sqmuxa_1_7\
        );

    \I__3306\ : InMux
    port map (
            O => \N__18426\,
            I => \N__18423\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__18423\,
            I => \this_ppu.un1_M_oam_idx_q_1_c3\
        );

    \I__3304\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18414\
        );

    \I__3303\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18414\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__18414\,
            I => \this_ppu.un1_M_oam_idx_q_1_c1\
        );

    \I__3301\ : InMux
    port map (
            O => \N__18411\,
            I => \N__18407\
        );

    \I__3300\ : InMux
    port map (
            O => \N__18410\,
            I => \N__18401\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__18407\,
            I => \N__18398\
        );

    \I__3298\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18391\
        );

    \I__3297\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18391\
        );

    \I__3296\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18391\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__18401\,
            I => \this_ppu.N_1156_0\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__18398\,
            I => \this_ppu.N_1156_0\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__18391\,
            I => \this_ppu.N_1156_0\
        );

    \I__3292\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__18381\,
            I => \N__18378\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__18378\,
            I => \N__18374\
        );

    \I__3289\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18371\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__18374\,
            I => \this_vga_signals.N_97\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__18371\,
            I => \this_vga_signals.N_97\
        );

    \I__3286\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__18363\,
            I => \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_2_0\
        );

    \I__3284\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18357\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__18357\,
            I => \this_vga_signals.N_154\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__18354\,
            I => \this_vga_signals.N_62_cascade_\
        );

    \I__3281\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18348\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__18348\,
            I => \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0\
        );

    \I__3279\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18339\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__18339\,
            I => \N__18336\
        );

    \I__3276\ : Sp12to4
    port map (
            O => \N__18336\,
            I => \N__18333\
        );

    \I__3275\ : Span12Mux_h
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__3274\ : Odrv12
    port map (
            O => \N__18330\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__18327\,
            I => \N__18322\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__18326\,
            I => \N__18318\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__18325\,
            I => \N__18314\
        );

    \I__3270\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18310\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__18321\,
            I => \N__18307\
        );

    \I__3268\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18303\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__18317\,
            I => \N__18300\
        );

    \I__3266\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18296\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__18313\,
            I => \N__18293\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__18310\,
            I => \N__18289\
        );

    \I__3263\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18286\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__18306\,
            I => \N__18283\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__18303\,
            I => \N__18279\
        );

    \I__3260\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18276\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__18299\,
            I => \N__18273\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18269\
        );

    \I__3257\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18266\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__18292\,
            I => \N__18263\
        );

    \I__3255\ : Span4Mux_v
    port map (
            O => \N__18289\,
            I => \N__18256\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__18286\,
            I => \N__18256\
        );

    \I__3253\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18253\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__18282\,
            I => \N__18250\
        );

    \I__3251\ : Span4Mux_v
    port map (
            O => \N__18279\,
            I => \N__18243\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__18276\,
            I => \N__18243\
        );

    \I__3249\ : InMux
    port map (
            O => \N__18273\,
            I => \N__18240\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__18272\,
            I => \N__18237\
        );

    \I__3247\ : Span4Mux_s0_v
    port map (
            O => \N__18269\,
            I => \N__18232\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__18266\,
            I => \N__18232\
        );

    \I__3245\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18229\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__18262\,
            I => \N__18226\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__18261\,
            I => \N__18223\
        );

    \I__3242\ : Span4Mux_h
    port map (
            O => \N__18256\,
            I => \N__18218\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__18253\,
            I => \N__18218\
        );

    \I__3240\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18215\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__18249\,
            I => \N__18212\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__18248\,
            I => \N__18209\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__18243\,
            I => \N__18204\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__18240\,
            I => \N__18204\
        );

    \I__3235\ : InMux
    port map (
            O => \N__18237\,
            I => \N__18201\
        );

    \I__3234\ : Span4Mux_v
    port map (
            O => \N__18232\,
            I => \N__18198\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__18229\,
            I => \N__18195\
        );

    \I__3232\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18192\
        );

    \I__3231\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18189\
        );

    \I__3230\ : Span4Mux_v
    port map (
            O => \N__18218\,
            I => \N__18184\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__18215\,
            I => \N__18184\
        );

    \I__3228\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18181\
        );

    \I__3227\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18177\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__18204\,
            I => \N__18172\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__18201\,
            I => \N__18172\
        );

    \I__3224\ : Sp12to4
    port map (
            O => \N__18198\,
            I => \N__18167\
        );

    \I__3223\ : Sp12to4
    port map (
            O => \N__18195\,
            I => \N__18167\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__18192\,
            I => \N__18162\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__18189\,
            I => \N__18162\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__18184\,
            I => \N__18157\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__18181\,
            I => \N__18157\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__18180\,
            I => \N__18154\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__18177\,
            I => \N__18151\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__18172\,
            I => \N__18148\
        );

    \I__3215\ : Span12Mux_h
    port map (
            O => \N__18167\,
            I => \N__18145\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__18162\,
            I => \N__18140\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__18157\,
            I => \N__18140\
        );

    \I__3212\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18137\
        );

    \I__3211\ : Span12Mux_h
    port map (
            O => \N__18151\,
            I => \N__18134\
        );

    \I__3210\ : Sp12to4
    port map (
            O => \N__18148\,
            I => \N__18131\
        );

    \I__3209\ : Span12Mux_v
    port map (
            O => \N__18145\,
            I => \N__18124\
        );

    \I__3208\ : Sp12to4
    port map (
            O => \N__18140\,
            I => \N__18124\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__18137\,
            I => \N__18124\
        );

    \I__3206\ : Odrv12
    port map (
            O => \N__18134\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__3205\ : Odrv12
    port map (
            O => \N__18131\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__3204\ : Odrv12
    port map (
            O => \N__18124\,
            I => \M_this_ppu_sprites_addr_8\
        );

    \I__3203\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18114\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__3201\ : Span4Mux_v
    port map (
            O => \N__18111\,
            I => \N__18108\
        );

    \I__3200\ : Span4Mux_v
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__3199\ : Span4Mux_h
    port map (
            O => \N__18105\,
            I => \N__18102\
        );

    \I__3198\ : Span4Mux_h
    port map (
            O => \N__18102\,
            I => \N__18099\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__18099\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__18096\,
            I => \N__18093\
        );

    \I__3195\ : InMux
    port map (
            O => \N__18093\,
            I => \N__18089\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__18092\,
            I => \N__18086\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__18089\,
            I => \N__18082\
        );

    \I__3192\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18079\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__18085\,
            I => \N__18076\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__18082\,
            I => \N__18070\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__18079\,
            I => \N__18070\
        );

    \I__3188\ : InMux
    port map (
            O => \N__18076\,
            I => \N__18067\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__18075\,
            I => \N__18064\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__18070\,
            I => \N__18058\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__18067\,
            I => \N__18058\
        );

    \I__3184\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18055\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__18063\,
            I => \N__18052\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__18058\,
            I => \N__18045\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__18055\,
            I => \N__18045\
        );

    \I__3180\ : InMux
    port map (
            O => \N__18052\,
            I => \N__18042\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__18051\,
            I => \N__18039\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \N__18035\
        );

    \I__3177\ : Span4Mux_v
    port map (
            O => \N__18045\,
            I => \N__18029\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__18042\,
            I => \N__18029\
        );

    \I__3175\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18026\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__18038\,
            I => \N__18023\
        );

    \I__3173\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18014\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__18034\,
            I => \N__18011\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__18029\,
            I => \N__18006\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__18026\,
            I => \N__18006\
        );

    \I__3169\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18003\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__18022\,
            I => \N__18000\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__18021\,
            I => \N__17996\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__18020\,
            I => \N__17993\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__18019\,
            I => \N__17990\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__18018\,
            I => \N__17987\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__18017\,
            I => \N__17984\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__18014\,
            I => \N__17981\
        );

    \I__3161\ : InMux
    port map (
            O => \N__18011\,
            I => \N__17978\
        );

    \I__3160\ : Span4Mux_v
    port map (
            O => \N__18006\,
            I => \N__17973\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__18003\,
            I => \N__17973\
        );

    \I__3158\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17970\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__17999\,
            I => \N__17967\
        );

    \I__3156\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17964\
        );

    \I__3155\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17961\
        );

    \I__3154\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17958\
        );

    \I__3153\ : InMux
    port map (
            O => \N__17987\,
            I => \N__17955\
        );

    \I__3152\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17952\
        );

    \I__3151\ : Span4Mux_h
    port map (
            O => \N__17981\,
            I => \N__17947\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__17978\,
            I => \N__17947\
        );

    \I__3149\ : Span4Mux_h
    port map (
            O => \N__17973\,
            I => \N__17942\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__17970\,
            I => \N__17942\
        );

    \I__3147\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17939\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__17964\,
            I => \N__17928\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__17961\,
            I => \N__17928\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__17958\,
            I => \N__17928\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__17955\,
            I => \N__17928\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__17952\,
            I => \N__17928\
        );

    \I__3141\ : Span4Mux_v
    port map (
            O => \N__17947\,
            I => \N__17925\
        );

    \I__3140\ : Span4Mux_v
    port map (
            O => \N__17942\,
            I => \N__17920\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__17939\,
            I => \N__17920\
        );

    \I__3138\ : Span12Mux_v
    port map (
            O => \N__17928\,
            I => \N__17917\
        );

    \I__3137\ : Sp12to4
    port map (
            O => \N__17925\,
            I => \N__17912\
        );

    \I__3136\ : Sp12to4
    port map (
            O => \N__17920\,
            I => \N__17912\
        );

    \I__3135\ : Odrv12
    port map (
            O => \N__17917\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__3134\ : Odrv12
    port map (
            O => \N__17912\,
            I => \M_this_ppu_sprites_addr_7\
        );

    \I__3133\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17901\
        );

    \I__3132\ : InMux
    port map (
            O => \N__17906\,
            I => \N__17901\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__17901\,
            I => \N__17898\
        );

    \I__3130\ : Span12Mux_h
    port map (
            O => \N__17898\,
            I => \N__17895\
        );

    \I__3129\ : Span12Mux_v
    port map (
            O => \N__17895\,
            I => \N__17892\
        );

    \I__3128\ : Odrv12
    port map (
            O => \N__17892\,
            I => port_address_in_7
        );

    \I__3127\ : IoInMux
    port map (
            O => \N__17889\,
            I => \N__17886\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__17886\,
            I => \N__17883\
        );

    \I__3125\ : Span12Mux_s3_h
    port map (
            O => \N__17883\,
            I => \N__17880\
        );

    \I__3124\ : Span12Mux_h
    port map (
            O => \N__17880\,
            I => \N__17876\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__17879\,
            I => \N__17873\
        );

    \I__3122\ : Span12Mux_v
    port map (
            O => \N__17876\,
            I => \N__17869\
        );

    \I__3121\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17864\
        );

    \I__3120\ : InMux
    port map (
            O => \N__17872\,
            I => \N__17864\
        );

    \I__3119\ : Odrv12
    port map (
            O => \N__17869\,
            I => led_c_1
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__17864\,
            I => led_c_1
        );

    \I__3117\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17855\
        );

    \I__3116\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17852\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__17855\,
            I => \N__17849\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__17852\,
            I => \N__17846\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__17849\,
            I => \N__17843\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__17846\,
            I => \N_84\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__17843\,
            I => \N_84\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__17838\,
            I => \N__17833\
        );

    \I__3109\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17828\
        );

    \I__3108\ : InMux
    port map (
            O => \N__17836\,
            I => \N__17823\
        );

    \I__3107\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17823\
        );

    \I__3106\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17819\
        );

    \I__3105\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17816\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17810\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__17823\,
            I => \N__17810\
        );

    \I__3102\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17807\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__17819\,
            I => \N__17804\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17801\
        );

    \I__3099\ : InMux
    port map (
            O => \N__17815\,
            I => \N__17798\
        );

    \I__3098\ : Span4Mux_v
    port map (
            O => \N__17810\,
            I => \N__17795\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__17807\,
            I => \N__17792\
        );

    \I__3096\ : Span4Mux_h
    port map (
            O => \N__17804\,
            I => \N__17785\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__17801\,
            I => \N__17785\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__17798\,
            I => \N__17785\
        );

    \I__3093\ : Span4Mux_v
    port map (
            O => \N__17795\,
            I => \N__17782\
        );

    \I__3092\ : Span4Mux_v
    port map (
            O => \N__17792\,
            I => \N__17777\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__17785\,
            I => \N__17777\
        );

    \I__3090\ : Sp12to4
    port map (
            O => \N__17782\,
            I => \N__17772\
        );

    \I__3089\ : Sp12to4
    port map (
            O => \N__17777\,
            I => \N__17772\
        );

    \I__3088\ : Span12Mux_h
    port map (
            O => \N__17772\,
            I => \N__17769\
        );

    \I__3087\ : Odrv12
    port map (
            O => \N__17769\,
            I => port_address_in_1
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__17766\,
            I => \N__17762\
        );

    \I__3085\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17758\
        );

    \I__3084\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17750\
        );

    \I__3083\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17750\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17747\
        );

    \I__3081\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17744\
        );

    \I__3080\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17741\
        );

    \I__3079\ : InMux
    port map (
            O => \N__17755\,
            I => \N__17738\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__17750\,
            I => \N__17734\
        );

    \I__3077\ : Span4Mux_h
    port map (
            O => \N__17747\,
            I => \N__17727\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__17744\,
            I => \N__17727\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17727\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__17738\,
            I => \N__17724\
        );

    \I__3073\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17721\
        );

    \I__3072\ : Span4Mux_v
    port map (
            O => \N__17734\,
            I => \N__17718\
        );

    \I__3071\ : Span4Mux_v
    port map (
            O => \N__17727\,
            I => \N__17715\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__17724\,
            I => \N__17710\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__17721\,
            I => \N__17710\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__17718\,
            I => \N__17707\
        );

    \I__3067\ : Span4Mux_v
    port map (
            O => \N__17715\,
            I => \N__17704\
        );

    \I__3066\ : Sp12to4
    port map (
            O => \N__17710\,
            I => \N__17701\
        );

    \I__3065\ : Sp12to4
    port map (
            O => \N__17707\,
            I => \N__17698\
        );

    \I__3064\ : Sp12to4
    port map (
            O => \N__17704\,
            I => \N__17693\
        );

    \I__3063\ : Span12Mux_v
    port map (
            O => \N__17701\,
            I => \N__17693\
        );

    \I__3062\ : Span12Mux_h
    port map (
            O => \N__17698\,
            I => \N__17690\
        );

    \I__3061\ : Span12Mux_h
    port map (
            O => \N__17693\,
            I => \N__17687\
        );

    \I__3060\ : Odrv12
    port map (
            O => \N__17690\,
            I => port_address_in_4
        );

    \I__3059\ : Odrv12
    port map (
            O => \N__17687\,
            I => port_address_in_4
        );

    \I__3058\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17677\
        );

    \I__3057\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17672\
        );

    \I__3056\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17672\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__17677\,
            I => \N__17665\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__17672\,
            I => \N__17665\
        );

    \I__3053\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17662\
        );

    \I__3052\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17659\
        );

    \I__3051\ : Span4Mux_v
    port map (
            O => \N__17665\,
            I => \N__17655\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__17662\,
            I => \N__17652\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__17659\,
            I => \N__17649\
        );

    \I__3048\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17646\
        );

    \I__3047\ : Span4Mux_v
    port map (
            O => \N__17655\,
            I => \N__17642\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__17652\,
            I => \N__17635\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__17649\,
            I => \N__17635\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__17646\,
            I => \N__17635\
        );

    \I__3043\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17632\
        );

    \I__3042\ : Sp12to4
    port map (
            O => \N__17642\,
            I => \N__17629\
        );

    \I__3041\ : Span4Mux_v
    port map (
            O => \N__17635\,
            I => \N__17626\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__17632\,
            I => \N__17623\
        );

    \I__3039\ : Span12Mux_h
    port map (
            O => \N__17629\,
            I => \N__17618\
        );

    \I__3038\ : Sp12to4
    port map (
            O => \N__17626\,
            I => \N__17618\
        );

    \I__3037\ : Span12Mux_v
    port map (
            O => \N__17623\,
            I => \N__17615\
        );

    \I__3036\ : Odrv12
    port map (
            O => \N__17618\,
            I => port_address_in_0
        );

    \I__3035\ : Odrv12
    port map (
            O => \N__17615\,
            I => port_address_in_0
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__17610\,
            I => \N__17607\
        );

    \I__3033\ : InMux
    port map (
            O => \N__17607\,
            I => \N__17603\
        );

    \I__3032\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17600\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__17603\,
            I => \N__17597\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__17600\,
            I => \N__17594\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__17597\,
            I => \N__17591\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__17594\,
            I => \N__17588\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__17591\,
            I => \N_36\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__17588\,
            I => \N_36\
        );

    \I__3025\ : InMux
    port map (
            O => \N__17583\,
            I => \N__17569\
        );

    \I__3024\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17569\
        );

    \I__3023\ : InMux
    port map (
            O => \N__17581\,
            I => \N__17560\
        );

    \I__3022\ : InMux
    port map (
            O => \N__17580\,
            I => \N__17560\
        );

    \I__3021\ : InMux
    port map (
            O => \N__17579\,
            I => \N__17560\
        );

    \I__3020\ : InMux
    port map (
            O => \N__17578\,
            I => \N__17560\
        );

    \I__3019\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17551\
        );

    \I__3018\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17551\
        );

    \I__3017\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17551\
        );

    \I__3016\ : InMux
    port map (
            O => \N__17574\,
            I => \N__17551\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__17569\,
            I => \N__17547\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__17560\,
            I => \N__17542\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__17551\,
            I => \N__17542\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__17550\,
            I => \N__17539\
        );

    \I__3011\ : Span4Mux_v
    port map (
            O => \N__17547\,
            I => \N__17534\
        );

    \I__3010\ : Span4Mux_v
    port map (
            O => \N__17542\,
            I => \N__17534\
        );

    \I__3009\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17531\
        );

    \I__3008\ : Sp12to4
    port map (
            O => \N__17534\,
            I => \N__17528\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__17531\,
            I => \N__17525\
        );

    \I__3006\ : Span12Mux_h
    port map (
            O => \N__17528\,
            I => \N__17522\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__17525\,
            I => \N_164\
        );

    \I__3004\ : Odrv12
    port map (
            O => \N__17522\,
            I => \N_164\
        );

    \I__3003\ : InMux
    port map (
            O => \N__17517\,
            I => \N__17514\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__17514\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_8\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__17511\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_8_cascade_\
        );

    \I__3000\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17505\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__17505\,
            I => \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_8\
        );

    \I__2998\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17498\
        );

    \I__2997\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17495\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__17498\,
            I => \N__17492\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__17495\,
            I => \N__17489\
        );

    \I__2994\ : Span4Mux_h
    port map (
            O => \N__17492\,
            I => \N__17486\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__17489\,
            I => \N__17483\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__17486\,
            I => \this_vga_signals.N_124_0\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__17483\,
            I => \this_vga_signals.N_124_0\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__17478\,
            I => \this_vga_signals.N_154_cascade_\
        );

    \I__2989\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17472\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17469\
        );

    \I__2987\ : Span4Mux_h
    port map (
            O => \N__17469\,
            I => \N__17466\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__17466\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__17463\,
            I => \this_vga_signals.N_153_0_cascade_\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__17460\,
            I => \N_686_i_cascade_\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__17457\,
            I => \N__17454\
        );

    \I__2982\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17451\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__17451\,
            I => \this_vga_signals.M_this_state_q_srsts_i_1Z0Z_11\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__17448\,
            I => \N__17445\
        );

    \I__2979\ : InMux
    port map (
            O => \N__17445\,
            I => \N__17442\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__17442\,
            I => \N__17439\
        );

    \I__2977\ : Odrv12
    port map (
            O => \N__17439\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0Z0Z_3\
        );

    \I__2976\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17429\
        );

    \I__2975\ : CEMux
    port map (
            O => \N__17435\,
            I => \N__17424\
        );

    \I__2974\ : CEMux
    port map (
            O => \N__17434\,
            I => \N__17421\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__17433\,
            I => \N__17418\
        );

    \I__2972\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17415\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__17429\,
            I => \N__17412\
        );

    \I__2970\ : InMux
    port map (
            O => \N__17428\,
            I => \N__17407\
        );

    \I__2969\ : InMux
    port map (
            O => \N__17427\,
            I => \N__17407\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__17424\,
            I => \N__17401\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__17421\,
            I => \N__17401\
        );

    \I__2966\ : InMux
    port map (
            O => \N__17418\,
            I => \N__17398\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__17415\,
            I => \N__17394\
        );

    \I__2964\ : Span4Mux_v
    port map (
            O => \N__17412\,
            I => \N__17389\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__17407\,
            I => \N__17389\
        );

    \I__2962\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17386\
        );

    \I__2961\ : Span4Mux_v
    port map (
            O => \N__17401\,
            I => \N__17379\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__17398\,
            I => \N__17379\
        );

    \I__2959\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17376\
        );

    \I__2958\ : Span4Mux_v
    port map (
            O => \N__17394\,
            I => \N__17368\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__17389\,
            I => \N__17368\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__17386\,
            I => \N__17368\
        );

    \I__2955\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17363\
        );

    \I__2954\ : InMux
    port map (
            O => \N__17384\,
            I => \N__17363\
        );

    \I__2953\ : Span4Mux_v
    port map (
            O => \N__17379\,
            I => \N__17360\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__17376\,
            I => \N__17357\
        );

    \I__2951\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17354\
        );

    \I__2950\ : Span4Mux_h
    port map (
            O => \N__17368\,
            I => \N__17349\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__17363\,
            I => \N__17349\
        );

    \I__2948\ : Span4Mux_h
    port map (
            O => \N__17360\,
            I => \N__17346\
        );

    \I__2947\ : Span12Mux_h
    port map (
            O => \N__17357\,
            I => \N__17341\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__17354\,
            I => \N__17341\
        );

    \I__2945\ : Span4Mux_v
    port map (
            O => \N__17349\,
            I => \N__17336\
        );

    \I__2944\ : Span4Mux_h
    port map (
            O => \N__17346\,
            I => \N__17336\
        );

    \I__2943\ : Odrv12
    port map (
            O => \N__17341\,
            I => \M_this_state_d_0_sqmuxa_1\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__17336\,
            I => \M_this_state_d_0_sqmuxa_1\
        );

    \I__2941\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17328\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__17328\,
            I => \N__17325\
        );

    \I__2939\ : Span4Mux_h
    port map (
            O => \N__17325\,
            I => \N__17322\
        );

    \I__2938\ : Span4Mux_h
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__17319\,
            I => \M_this_map_ram_write_data_7\
        );

    \I__2936\ : IoInMux
    port map (
            O => \N__17316\,
            I => \N__17313\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__17313\,
            I => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\
        );

    \I__2934\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17302\
        );

    \I__2933\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17296\
        );

    \I__2932\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17289\
        );

    \I__2931\ : InMux
    port map (
            O => \N__17307\,
            I => \N__17289\
        );

    \I__2930\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17289\
        );

    \I__2929\ : CEMux
    port map (
            O => \N__17305\,
            I => \N__17279\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__17302\,
            I => \N__17276\
        );

    \I__2927\ : InMux
    port map (
            O => \N__17301\,
            I => \N__17273\
        );

    \I__2926\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17263\
        );

    \I__2925\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17263\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__17296\,
            I => \N__17260\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17257\
        );

    \I__2922\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17254\
        );

    \I__2921\ : InMux
    port map (
            O => \N__17287\,
            I => \N__17248\
        );

    \I__2920\ : InMux
    port map (
            O => \N__17286\,
            I => \N__17248\
        );

    \I__2919\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17243\
        );

    \I__2918\ : InMux
    port map (
            O => \N__17284\,
            I => \N__17243\
        );

    \I__2917\ : InMux
    port map (
            O => \N__17283\,
            I => \N__17240\
        );

    \I__2916\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17237\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__17279\,
            I => \N__17234\
        );

    \I__2914\ : Span4Mux_v
    port map (
            O => \N__17276\,
            I => \N__17229\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17229\
        );

    \I__2912\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17226\
        );

    \I__2911\ : InMux
    port map (
            O => \N__17271\,
            I => \N__17217\
        );

    \I__2910\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17217\
        );

    \I__2909\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17217\
        );

    \I__2908\ : InMux
    port map (
            O => \N__17268\,
            I => \N__17217\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__17263\,
            I => \N__17212\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__17260\,
            I => \N__17212\
        );

    \I__2905\ : Span4Mux_h
    port map (
            O => \N__17257\,
            I => \N__17207\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__17254\,
            I => \N__17207\
        );

    \I__2903\ : InMux
    port map (
            O => \N__17253\,
            I => \N__17204\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__17248\,
            I => \N__17195\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__17243\,
            I => \N__17195\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__17240\,
            I => \N__17195\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__17237\,
            I => \N__17195\
        );

    \I__2898\ : Span4Mux_h
    port map (
            O => \N__17234\,
            I => \N__17190\
        );

    \I__2897\ : Span4Mux_h
    port map (
            O => \N__17229\,
            I => \N__17190\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__17226\,
            I => \N__17187\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__17217\,
            I => \N__17184\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__17212\,
            I => \N__17177\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__17207\,
            I => \N__17177\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__17204\,
            I => \N__17177\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__17195\,
            I => \N__17174\
        );

    \I__2890\ : Span4Mux_h
    port map (
            O => \N__17190\,
            I => \N__17169\
        );

    \I__2889\ : Span4Mux_v
    port map (
            O => \N__17187\,
            I => \N__17169\
        );

    \I__2888\ : Odrv12
    port map (
            O => \N__17184\,
            I => \G_425\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__17177\,
            I => \G_425\
        );

    \I__2886\ : Odrv4
    port map (
            O => \N__17174\,
            I => \G_425\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__17169\,
            I => \G_425\
        );

    \I__2884\ : IoInMux
    port map (
            O => \N__17160\,
            I => \N__17157\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__17157\,
            I => \N__17154\
        );

    \I__2882\ : Span12Mux_s1_v
    port map (
            O => \N__17154\,
            I => \N__17151\
        );

    \I__2881\ : Odrv12
    port map (
            O => \N__17151\,
            I => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\
        );

    \I__2880\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17143\
        );

    \I__2879\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17138\
        );

    \I__2878\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17138\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__17143\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__17138\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__2875\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17129\
        );

    \I__2874\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17126\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__17129\,
            I => \N__17123\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__17126\,
            I => \this_vga_signals.M_vcounter_d8\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__17123\,
            I => \this_vga_signals.M_vcounter_d8\
        );

    \I__2870\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17112\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__17117\,
            I => \N__17109\
        );

    \I__2868\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17104\
        );

    \I__2867\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17101\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__17112\,
            I => \N__17098\
        );

    \I__2865\ : InMux
    port map (
            O => \N__17109\,
            I => \N__17095\
        );

    \I__2864\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17088\
        );

    \I__2863\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17088\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__17104\,
            I => \N__17085\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__17101\,
            I => \N__17078\
        );

    \I__2860\ : Span4Mux_v
    port map (
            O => \N__17098\,
            I => \N__17078\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__17095\,
            I => \N__17078\
        );

    \I__2858\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17075\
        );

    \I__2857\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17072\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__17088\,
            I => \N__17068\
        );

    \I__2855\ : Span4Mux_h
    port map (
            O => \N__17085\,
            I => \N__17062\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__17078\,
            I => \N__17062\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__17075\,
            I => \N__17057\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__17072\,
            I => \N__17057\
        );

    \I__2851\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17053\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__17068\,
            I => \N__17050\
        );

    \I__2849\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17047\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__17062\,
            I => \N__17044\
        );

    \I__2847\ : Span12Mux_v
    port map (
            O => \N__17057\,
            I => \N__17041\
        );

    \I__2846\ : InMux
    port map (
            O => \N__17056\,
            I => \N__17038\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__17035\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__17050\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__17047\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__17044\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2841\ : Odrv12
    port map (
            O => \N__17041\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__17038\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__17035\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__17022\,
            I => \N__17019\
        );

    \I__2837\ : InMux
    port map (
            O => \N__17019\,
            I => \N__17016\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__17016\,
            I => \N__17012\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__17015\,
            I => \N__17009\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__17012\,
            I => \N__17006\
        );

    \I__2833\ : InMux
    port map (
            O => \N__17009\,
            I => \N__17003\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__17006\,
            I => \N__16998\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__17003\,
            I => \N__16998\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__16998\,
            I => \this_vga_signals.un1_M_hcounter_d7_1_0\
        );

    \I__2829\ : CEMux
    port map (
            O => \N__16995\,
            I => \N__16992\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__16992\,
            I => \N__16988\
        );

    \I__2827\ : CEMux
    port map (
            O => \N__16991\,
            I => \N__16985\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__16988\,
            I => \N__16980\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__16985\,
            I => \N__16980\
        );

    \I__2824\ : Span4Mux_h
    port map (
            O => \N__16980\,
            I => \N__16977\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__16977\,
            I => \N__16974\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__16974\,
            I => \this_sprites_ram.mem_WE_6\
        );

    \I__2821\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16968\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__16968\,
            I => \N__16965\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__16965\,
            I => \this_vga_signals.M_this_state_q_srsts_i_i_1Z0Z_10\
        );

    \I__2818\ : CEMux
    port map (
            O => \N__16962\,
            I => \N__16959\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__16959\,
            I => \N__16956\
        );

    \I__2816\ : Span4Mux_h
    port map (
            O => \N__16956\,
            I => \N__16952\
        );

    \I__2815\ : CEMux
    port map (
            O => \N__16955\,
            I => \N__16949\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__16952\,
            I => \N__16946\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__16949\,
            I => \N__16943\
        );

    \I__2812\ : Span4Mux_h
    port map (
            O => \N__16946\,
            I => \N__16940\
        );

    \I__2811\ : Span12Mux_v
    port map (
            O => \N__16943\,
            I => \N__16937\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__16940\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__2809\ : Odrv12
    port map (
            O => \N__16937\,
            I => \this_sprites_ram.mem_WE_10\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__16932\,
            I => \N__16929\
        );

    \I__2807\ : InMux
    port map (
            O => \N__16929\,
            I => \N__16925\
        );

    \I__2806\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16922\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__16925\,
            I => \this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__16922\,
            I => \this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__16917\,
            I => \N__16914\
        );

    \I__2802\ : InMux
    port map (
            O => \N__16914\,
            I => \N__16911\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__16911\,
            I => \N__16908\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__16908\,
            I => \N__16905\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__16905\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_6\
        );

    \I__2798\ : InMux
    port map (
            O => \N__16902\,
            I => \N__16893\
        );

    \I__2797\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16893\
        );

    \I__2796\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16888\
        );

    \I__2795\ : InMux
    port map (
            O => \N__16899\,
            I => \N__16888\
        );

    \I__2794\ : InMux
    port map (
            O => \N__16898\,
            I => \N__16885\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__16893\,
            I => \this_vga_signals.N_85\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__16888\,
            I => \this_vga_signals.N_85\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__16885\,
            I => \this_vga_signals.N_85\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__16878\,
            I => \N__16875\
        );

    \I__2789\ : InMux
    port map (
            O => \N__16875\,
            I => \N__16872\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__16872\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_4\
        );

    \I__2787\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16865\
        );

    \I__2786\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16862\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__16865\,
            I => \N__16856\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__16862\,
            I => \N__16856\
        );

    \I__2783\ : InMux
    port map (
            O => \N__16861\,
            I => \N__16853\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__16856\,
            I => \N__16850\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__16853\,
            I => \N__16847\
        );

    \I__2780\ : Span4Mux_h
    port map (
            O => \N__16850\,
            I => \N__16844\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__16847\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2778\ : Odrv4
    port map (
            O => \N__16844\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__2777\ : InMux
    port map (
            O => \N__16839\,
            I => \N__16836\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__16836\,
            I => \N__16833\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__16833\,
            I => \this_vga_signals.CO0\
        );

    \I__2774\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16824\
        );

    \I__2773\ : InMux
    port map (
            O => \N__16829\,
            I => \N__16824\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__16824\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__2771\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16816\
        );

    \I__2770\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16811\
        );

    \I__2769\ : InMux
    port map (
            O => \N__16819\,
            I => \N__16811\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__16816\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__16811\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__16806\,
            I => \this_vga_signals.N_152_0_cascade_\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__16803\,
            I => \N__16800\
        );

    \I__2764\ : InMux
    port map (
            O => \N__16800\,
            I => \N__16797\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__16797\,
            I => \N__16794\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__16794\,
            I => \this_vga_signals.M_vcounter_d7lto8_1\
        );

    \I__2761\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16785\
        );

    \I__2760\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16785\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__16785\,
            I => \this_vga_signals.M_vcounter_d7lt8_0\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__16782\,
            I => \N__16772\
        );

    \I__2757\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16763\
        );

    \I__2756\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16763\
        );

    \I__2755\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16756\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__16778\,
            I => \N__16753\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__16777\,
            I => \N__16750\
        );

    \I__2752\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16747\
        );

    \I__2751\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16743\
        );

    \I__2750\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16738\
        );

    \I__2749\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16738\
        );

    \I__2748\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16731\
        );

    \I__2747\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16731\
        );

    \I__2746\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16731\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__16763\,
            I => \N__16728\
        );

    \I__2744\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16723\
        );

    \I__2743\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16723\
        );

    \I__2742\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16718\
        );

    \I__2741\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16718\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__16756\,
            I => \N__16712\
        );

    \I__2739\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16703\
        );

    \I__2738\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16703\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__16747\,
            I => \N__16700\
        );

    \I__2736\ : InMux
    port map (
            O => \N__16746\,
            I => \N__16697\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__16743\,
            I => \N__16692\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__16738\,
            I => \N__16692\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__16731\,
            I => \N__16689\
        );

    \I__2732\ : Span4Mux_v
    port map (
            O => \N__16728\,
            I => \N__16684\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__16723\,
            I => \N__16684\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__16718\,
            I => \N__16681\
        );

    \I__2729\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16676\
        );

    \I__2728\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16676\
        );

    \I__2727\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16673\
        );

    \I__2726\ : Span4Mux_v
    port map (
            O => \N__16712\,
            I => \N__16670\
        );

    \I__2725\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16665\
        );

    \I__2724\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16665\
        );

    \I__2723\ : InMux
    port map (
            O => \N__16709\,
            I => \N__16660\
        );

    \I__2722\ : InMux
    port map (
            O => \N__16708\,
            I => \N__16660\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__16703\,
            I => \N__16655\
        );

    \I__2720\ : Span12Mux_s9_v
    port map (
            O => \N__16700\,
            I => \N__16655\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__16697\,
            I => \N__16642\
        );

    \I__2718\ : Span4Mux_v
    port map (
            O => \N__16692\,
            I => \N__16642\
        );

    \I__2717\ : Span4Mux_h
    port map (
            O => \N__16689\,
            I => \N__16642\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__16684\,
            I => \N__16642\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__16681\,
            I => \N__16642\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__16676\,
            I => \N__16642\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__16673\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__16670\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__16665\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__16660\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2709\ : Odrv12
    port map (
            O => \N__16655\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__16642\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2707\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16624\
        );

    \I__2706\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16621\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__16627\,
            I => \N__16616\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__16624\,
            I => \N__16611\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__16621\,
            I => \N__16607\
        );

    \I__2702\ : InMux
    port map (
            O => \N__16620\,
            I => \N__16604\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__16619\,
            I => \N__16599\
        );

    \I__2700\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16596\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__16615\,
            I => \N__16593\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__16614\,
            I => \N__16590\
        );

    \I__2697\ : Span4Mux_h
    port map (
            O => \N__16611\,
            I => \N__16587\
        );

    \I__2696\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16584\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__16607\,
            I => \N__16581\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__16604\,
            I => \N__16578\
        );

    \I__2693\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16573\
        );

    \I__2692\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16573\
        );

    \I__2691\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16570\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__16596\,
            I => \N__16567\
        );

    \I__2689\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16564\
        );

    \I__2688\ : InMux
    port map (
            O => \N__16590\,
            I => \N__16561\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__16587\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__16584\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__16581\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__16578\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__16573\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__16570\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__16567\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__16564\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__16561\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2678\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16533\
        );

    \I__2677\ : InMux
    port map (
            O => \N__16541\,
            I => \N__16530\
        );

    \I__2676\ : InMux
    port map (
            O => \N__16540\,
            I => \N__16523\
        );

    \I__2675\ : InMux
    port map (
            O => \N__16539\,
            I => \N__16523\
        );

    \I__2674\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16523\
        );

    \I__2673\ : InMux
    port map (
            O => \N__16537\,
            I => \N__16518\
        );

    \I__2672\ : InMux
    port map (
            O => \N__16536\,
            I => \N__16518\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__16533\,
            I => \N__16512\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__16530\,
            I => \N__16503\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__16523\,
            I => \N__16500\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__16518\,
            I => \N__16497\
        );

    \I__2667\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16494\
        );

    \I__2666\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16491\
        );

    \I__2665\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16488\
        );

    \I__2664\ : Span4Mux_v
    port map (
            O => \N__16512\,
            I => \N__16483\
        );

    \I__2663\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16478\
        );

    \I__2662\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16478\
        );

    \I__2661\ : InMux
    port map (
            O => \N__16509\,
            I => \N__16475\
        );

    \I__2660\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16472\
        );

    \I__2659\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16467\
        );

    \I__2658\ : InMux
    port map (
            O => \N__16506\,
            I => \N__16467\
        );

    \I__2657\ : Span4Mux_v
    port map (
            O => \N__16503\,
            I => \N__16458\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__16500\,
            I => \N__16458\
        );

    \I__2655\ : Span4Mux_v
    port map (
            O => \N__16497\,
            I => \N__16458\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16458\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__16491\,
            I => \N__16453\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__16488\,
            I => \N__16453\
        );

    \I__2651\ : InMux
    port map (
            O => \N__16487\,
            I => \N__16450\
        );

    \I__2650\ : InMux
    port map (
            O => \N__16486\,
            I => \N__16447\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__16483\,
            I => \N__16442\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__16478\,
            I => \N__16442\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__16475\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__16472\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__16467\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__16458\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2643\ : Odrv12
    port map (
            O => \N__16453\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__16450\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__16447\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__16442\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2639\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16420\
        );

    \I__2638\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16413\
        );

    \I__2637\ : InMux
    port map (
            O => \N__16423\,
            I => \N__16413\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__16420\,
            I => \N__16404\
        );

    \I__2635\ : InMux
    port map (
            O => \N__16419\,
            I => \N__16399\
        );

    \I__2634\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16399\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__16413\,
            I => \N__16396\
        );

    \I__2632\ : InMux
    port map (
            O => \N__16412\,
            I => \N__16391\
        );

    \I__2631\ : InMux
    port map (
            O => \N__16411\,
            I => \N__16391\
        );

    \I__2630\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16388\
        );

    \I__2629\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16383\
        );

    \I__2628\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16383\
        );

    \I__2627\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16380\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__16404\,
            I => \N__16371\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__16399\,
            I => \N__16371\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__16396\,
            I => \N__16371\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16391\,
            I => \N__16371\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__16388\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__16383\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__16380\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__16371\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__16362\,
            I => \this_vga_signals.line_clk_1_cascade_\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__16359\,
            I => \M_this_vga_signals_line_clk_0_cascade_\
        );

    \I__2616\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16350\
        );

    \I__2615\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16350\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__16350\,
            I => \this_vga_signals.un4_lvisibility_1\
        );

    \I__2613\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16343\
        );

    \I__2612\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16338\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__16343\,
            I => \N__16332\
        );

    \I__2610\ : InMux
    port map (
            O => \N__16342\,
            I => \N__16327\
        );

    \I__2609\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16327\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__16338\,
            I => \N__16324\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__16337\,
            I => \N__16321\
        );

    \I__2606\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16316\
        );

    \I__2605\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16313\
        );

    \I__2604\ : Span4Mux_v
    port map (
            O => \N__16332\,
            I => \N__16306\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__16327\,
            I => \N__16306\
        );

    \I__2602\ : Span4Mux_v
    port map (
            O => \N__16324\,
            I => \N__16306\
        );

    \I__2601\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16301\
        );

    \I__2600\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16301\
        );

    \I__2599\ : InMux
    port map (
            O => \N__16319\,
            I => \N__16298\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__16316\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__16313\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__16306\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__16301\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__16298\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__16287\,
            I => \N__16284\
        );

    \I__2592\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16281\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__16281\,
            I => \this_vga_signals.line_clk_1\
        );

    \I__2590\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16275\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__16275\,
            I => \N__16263\
        );

    \I__2588\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16258\
        );

    \I__2587\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16258\
        );

    \I__2586\ : InMux
    port map (
            O => \N__16272\,
            I => \N__16255\
        );

    \I__2585\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16250\
        );

    \I__2584\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16250\
        );

    \I__2583\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16245\
        );

    \I__2582\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16245\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16242\
        );

    \I__2580\ : InMux
    port map (
            O => \N__16266\,
            I => \N__16239\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__16263\,
            I => \N__16234\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__16258\,
            I => \N__16234\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__16255\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__16250\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__16245\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__16242\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__16239\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2572\ : Odrv4
    port map (
            O => \N__16234\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__16221\,
            I => \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0Z0Z_2_cascade_\
        );

    \I__2570\ : InMux
    port map (
            O => \N__16218\,
            I => \N__16213\
        );

    \I__2569\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16208\
        );

    \I__2568\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16208\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__16213\,
            I => \M_this_substate_qZ0\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__16208\,
            I => \M_this_substate_qZ0\
        );

    \I__2565\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16200\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__16200\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__2563\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16194\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16191\
        );

    \I__2561\ : Span12Mux_s10_h
    port map (
            O => \N__16191\,
            I => \N__16188\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__16188\,
            I => \M_this_map_ram_write_data_3\
        );

    \I__2559\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16182\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__16182\,
            I => \N__16179\
        );

    \I__2557\ : Odrv12
    port map (
            O => \N__16179\,
            I => \M_this_map_ram_write_data_2\
        );

    \I__2556\ : InMux
    port map (
            O => \N__16176\,
            I => \N__16171\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__16175\,
            I => \N__16167\
        );

    \I__2554\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16164\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__16171\,
            I => \N__16161\
        );

    \I__2552\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16156\
        );

    \I__2551\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16156\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__16164\,
            I => \N__16152\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__16161\,
            I => \N__16148\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__16156\,
            I => \N__16145\
        );

    \I__2547\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16142\
        );

    \I__2546\ : Span4Mux_h
    port map (
            O => \N__16152\,
            I => \N__16138\
        );

    \I__2545\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16135\
        );

    \I__2544\ : Sp12to4
    port map (
            O => \N__16148\,
            I => \N__16128\
        );

    \I__2543\ : Sp12to4
    port map (
            O => \N__16145\,
            I => \N__16128\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__16142\,
            I => \N__16128\
        );

    \I__2541\ : InMux
    port map (
            O => \N__16141\,
            I => \N__16125\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__16138\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__16135\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2538\ : Odrv12
    port map (
            O => \N__16128\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__16125\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2536\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16112\
        );

    \I__2535\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16109\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__16112\,
            I => \N__16106\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__16109\,
            I => \N__16100\
        );

    \I__2532\ : Span4Mux_h
    port map (
            O => \N__16106\,
            I => \N__16100\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16097\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__16100\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__16097\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__16092\,
            I => \N__16086\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__16091\,
            I => \N__16080\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__16090\,
            I => \N__16075\
        );

    \I__2525\ : InMux
    port map (
            O => \N__16089\,
            I => \N__16072\
        );

    \I__2524\ : InMux
    port map (
            O => \N__16086\,
            I => \N__16068\
        );

    \I__2523\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16063\
        );

    \I__2522\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16063\
        );

    \I__2521\ : InMux
    port map (
            O => \N__16083\,
            I => \N__16058\
        );

    \I__2520\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16058\
        );

    \I__2519\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16055\
        );

    \I__2518\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16052\
        );

    \I__2517\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16049\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__16072\,
            I => \N__16044\
        );

    \I__2515\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16041\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__16068\,
            I => \N__16036\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__16063\,
            I => \N__16036\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__16058\,
            I => \N__16027\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__16055\,
            I => \N__16027\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__16052\,
            I => \N__16027\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__16049\,
            I => \N__16027\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__16048\,
            I => \N__16024\
        );

    \I__2507\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16021\
        );

    \I__2506\ : Span4Mux_h
    port map (
            O => \N__16044\,
            I => \N__16018\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__16041\,
            I => \N__16011\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__16036\,
            I => \N__16011\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__16027\,
            I => \N__16011\
        );

    \I__2502\ : InMux
    port map (
            O => \N__16024\,
            I => \N__16008\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__16021\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__16018\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__16011\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__16008\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__15999\,
            I => \N__15995\
        );

    \I__2496\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15976\
        );

    \I__2495\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15971\
        );

    \I__2494\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15971\
        );

    \I__2493\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15968\
        );

    \I__2492\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15965\
        );

    \I__2491\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15962\
        );

    \I__2490\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15953\
        );

    \I__2489\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15953\
        );

    \I__2488\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15953\
        );

    \I__2487\ : InMux
    port map (
            O => \N__15987\,
            I => \N__15953\
        );

    \I__2486\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15950\
        );

    \I__2485\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15947\
        );

    \I__2484\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15942\
        );

    \I__2483\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15942\
        );

    \I__2482\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15936\
        );

    \I__2481\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15936\
        );

    \I__2480\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15931\
        );

    \I__2479\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15931\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__15976\,
            I => \N__15926\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15926\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__15968\,
            I => \N__15915\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__15965\,
            I => \N__15915\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__15962\,
            I => \N__15915\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__15953\,
            I => \N__15915\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__15950\,
            I => \N__15915\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__15947\,
            I => \N__15910\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__15942\,
            I => \N__15910\
        );

    \I__2469\ : InMux
    port map (
            O => \N__15941\,
            I => \N__15906\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__15936\,
            I => \N__15903\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__15931\,
            I => \N__15896\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__15926\,
            I => \N__15896\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__15915\,
            I => \N__15896\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__15910\,
            I => \N__15893\
        );

    \I__2463\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15890\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__15906\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2461\ : Odrv12
    port map (
            O => \N__15903\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__15896\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__15893\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__15890\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2457\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15874\
        );

    \I__2456\ : InMux
    port map (
            O => \N__15878\,
            I => \N__15869\
        );

    \I__2455\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15869\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__15874\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__15869\,
            I => \this_ppu.M_count_qZ0Z_5\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__15864\,
            I => \N__15861\
        );

    \I__2451\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15856\
        );

    \I__2450\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15853\
        );

    \I__2449\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15850\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__15856\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__15853\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__15850\,
            I => \this_ppu.M_count_qZ0Z_4\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__15843\,
            I => \N__15838\
        );

    \I__2444\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15835\
        );

    \I__2443\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15830\
        );

    \I__2442\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15830\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__15835\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__15830\,
            I => \this_ppu.M_count_qZ0Z_6\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__15825\,
            I => \N__15821\
        );

    \I__2438\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15817\
        );

    \I__2437\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15814\
        );

    \I__2436\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15811\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__15817\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__15814\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__15811\,
            I => \this_ppu.M_count_qZ0Z_2\
        );

    \I__2432\ : InMux
    port map (
            O => \N__15804\,
            I => \N__15799\
        );

    \I__2431\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15794\
        );

    \I__2430\ : InMux
    port map (
            O => \N__15802\,
            I => \N__15794\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__15799\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__15794\,
            I => \this_ppu.M_count_qZ0Z_1\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__15789\,
            I => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4_cascade_\
        );

    \I__2426\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15783\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__15783\,
            I => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__15780\,
            I => \N__15776\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__15779\,
            I => \N__15773\
        );

    \I__2422\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15758\
        );

    \I__2421\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15758\
        );

    \I__2420\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15758\
        );

    \I__2419\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15758\
        );

    \I__2418\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15758\
        );

    \I__2417\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15755\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__15758\,
            I => \this_ppu.un16_0\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__15755\,
            I => \this_ppu.un16_0\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__15750\,
            I => \N__15747\
        );

    \I__2413\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15744\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__15744\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\
        );

    \I__2411\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15726\
        );

    \I__2410\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15726\
        );

    \I__2409\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15726\
        );

    \I__2408\ : InMux
    port map (
            O => \N__15738\,
            I => \N__15726\
        );

    \I__2407\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15726\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__15726\,
            I => \this_ppu.N_1195_0\
        );

    \I__2405\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15719\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__15722\,
            I => \N__15716\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15712\
        );

    \I__2402\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15709\
        );

    \I__2401\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15706\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__15712\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__15709\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__15706\,
            I => \this_ppu.M_count_qZ0Z_3\
        );

    \I__2397\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15696\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__15696\,
            I => \this_ppu.M_count_q_RNO_0Z0Z_7\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__15693\,
            I => \N__15690\
        );

    \I__2394\ : InMux
    port map (
            O => \N__15690\,
            I => \N__15687\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__15687\,
            I => \N__15683\
        );

    \I__2392\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15680\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__15683\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__15680\,
            I => \this_ppu.M_count_qZ0Z_7\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__15675\,
            I => \this_vga_signals.N_85_cascade_\
        );

    \I__2388\ : InMux
    port map (
            O => \N__15672\,
            I => \N__15669\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__15669\,
            I => \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_5\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__15666\,
            I => \this_ppu.N_1195_0_cascade_\
        );

    \I__2385\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15660\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__15660\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\
        );

    \I__2383\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15653\
        );

    \I__2382\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15650\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__15653\,
            I => \this_ppu.N_1195_0_1\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__15650\,
            I => \this_ppu.N_1195_0_1\
        );

    \I__2379\ : InMux
    port map (
            O => \N__15645\,
            I => \N__15640\
        );

    \I__2378\ : InMux
    port map (
            O => \N__15644\,
            I => \N__15637\
        );

    \I__2377\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15634\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__15640\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__15637\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__15634\,
            I => \this_ppu.M_count_qZ0Z_0\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__15627\,
            I => \N__15624\
        );

    \I__2372\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15621\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__15621\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\
        );

    \I__2370\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15615\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__15615\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\
        );

    \I__2368\ : InMux
    port map (
            O => \N__15612\,
            I => \N__15609\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__15609\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\
        );

    \I__2366\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15603\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__15603\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\
        );

    \I__2364\ : InMux
    port map (
            O => \N__15600\,
            I => \N__15595\
        );

    \I__2363\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15592\
        );

    \I__2362\ : InMux
    port map (
            O => \N__15598\,
            I => \N__15589\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__15595\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__15592\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__15589\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__2358\ : InMux
    port map (
            O => \N__15582\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__2357\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15573\
        );

    \I__2356\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15573\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__15573\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__2354\ : InMux
    port map (
            O => \N__15570\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__2353\ : InMux
    port map (
            O => \N__15567\,
            I => \N__15562\
        );

    \I__2352\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15557\
        );

    \I__2351\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15557\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__15562\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__15557\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__2348\ : InMux
    port map (
            O => \N__15552\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__2347\ : InMux
    port map (
            O => \N__15549\,
            I => \N__15544\
        );

    \I__2346\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15539\
        );

    \I__2345\ : InMux
    port map (
            O => \N__15547\,
            I => \N__15539\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__15544\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__15539\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__2342\ : InMux
    port map (
            O => \N__15534\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__2341\ : InMux
    port map (
            O => \N__15531\,
            I => \bfn_15_10_0_\
        );

    \I__2340\ : InMux
    port map (
            O => \N__15528\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__2339\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15521\
        );

    \I__2338\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15518\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__15521\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__15518\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__2335\ : CEMux
    port map (
            O => \N__15513\,
            I => \N__15510\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__15510\,
            I => \N__15506\
        );

    \I__2333\ : CEMux
    port map (
            O => \N__15509\,
            I => \N__15501\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__15506\,
            I => \N__15498\
        );

    \I__2331\ : CEMux
    port map (
            O => \N__15505\,
            I => \N__15495\
        );

    \I__2330\ : CEMux
    port map (
            O => \N__15504\,
            I => \N__15492\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__15501\,
            I => \N__15483\
        );

    \I__2328\ : Span4Mux_v
    port map (
            O => \N__15498\,
            I => \N__15483\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__15495\,
            I => \N__15483\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__15492\,
            I => \N__15483\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__15483\,
            I => \this_vga_signals.N_852_0\
        );

    \I__2324\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15477\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__15477\,
            I => \N__15469\
        );

    \I__2322\ : SRMux
    port map (
            O => \N__15476\,
            I => \N__15456\
        );

    \I__2321\ : SRMux
    port map (
            O => \N__15475\,
            I => \N__15456\
        );

    \I__2320\ : SRMux
    port map (
            O => \N__15474\,
            I => \N__15456\
        );

    \I__2319\ : SRMux
    port map (
            O => \N__15473\,
            I => \N__15456\
        );

    \I__2318\ : SRMux
    port map (
            O => \N__15472\,
            I => \N__15456\
        );

    \I__2317\ : Glb2LocalMux
    port map (
            O => \N__15469\,
            I => \N__15456\
        );

    \I__2316\ : GlobalMux
    port map (
            O => \N__15456\,
            I => \N__15453\
        );

    \I__2315\ : gio2CtrlBuf
    port map (
            O => \N__15453\,
            I => \this_vga_signals.N_1098_g\
        );

    \I__2314\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15447\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__15447\,
            I => \N__15444\
        );

    \I__2312\ : Span12Mux_v
    port map (
            O => \N__15444\,
            I => \N__15441\
        );

    \I__2311\ : Span12Mux_h
    port map (
            O => \N__15441\,
            I => \N__15438\
        );

    \I__2310\ : Odrv12
    port map (
            O => \N__15438\,
            I => port_clk_c
        );

    \I__2309\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15432\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__15432\,
            I => \N__15429\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__15429\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__2306\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15423\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__15423\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__2304\ : InMux
    port map (
            O => \N__15420\,
            I => \N__15417\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__15417\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__2302\ : InMux
    port map (
            O => \N__15414\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__2301\ : InMux
    port map (
            O => \N__15411\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__2300\ : InMux
    port map (
            O => \N__15408\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__2299\ : InMux
    port map (
            O => \N__15405\,
            I => \this_ppu.un1_M_count_q_1_cry_0_s1\
        );

    \I__2298\ : InMux
    port map (
            O => \N__15402\,
            I => \this_ppu.un1_M_count_q_1_cry_1_s1\
        );

    \I__2297\ : InMux
    port map (
            O => \N__15399\,
            I => \this_ppu.un1_M_count_q_1_cry_2_s1\
        );

    \I__2296\ : InMux
    port map (
            O => \N__15396\,
            I => \this_ppu.un1_M_count_q_1_cry_3_s1\
        );

    \I__2295\ : InMux
    port map (
            O => \N__15393\,
            I => \this_ppu.un1_M_count_q_1_cry_4_s1\
        );

    \I__2294\ : InMux
    port map (
            O => \N__15390\,
            I => \this_ppu.un1_M_count_q_1_cry_5_s1\
        );

    \I__2293\ : InMux
    port map (
            O => \N__15387\,
            I => \this_ppu.un1_M_count_q_1_cry_6_s1\
        );

    \I__2292\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15381\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__15381\,
            I => \N__15378\
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__15378\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__15375\,
            I => \N__15372\
        );

    \I__2288\ : InMux
    port map (
            O => \N__15372\,
            I => \N__15367\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__15371\,
            I => \N__15361\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__15370\,
            I => \N__15358\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__15367\,
            I => \N__15355\
        );

    \I__2284\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15350\
        );

    \I__2283\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15350\
        );

    \I__2282\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15343\
        );

    \I__2281\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15343\
        );

    \I__2280\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15343\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__15355\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__15350\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__15343\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__15336\,
            I => \this_vga_signals.un6_vvisibilitylto8_0_cascade_\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__15333\,
            I => \this_vga_signals.un6_vvisibilitylt9_0_cascade_\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__15330\,
            I => \this_vga_signals_vvisibility_1_cascade_\
        );

    \I__2273\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15322\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15319\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__15325\,
            I => \N__15316\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15322\,
            I => \N__15313\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__15319\,
            I => \N__15310\
        );

    \I__2268\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15307\
        );

    \I__2267\ : Sp12to4
    port map (
            O => \N__15313\,
            I => \N__15304\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__15310\,
            I => \N__15299\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__15307\,
            I => \N__15299\
        );

    \I__2264\ : Span12Mux_s9_v
    port map (
            O => \N__15304\,
            I => \N__15296\
        );

    \I__2263\ : Span4Mux_h
    port map (
            O => \N__15299\,
            I => \N__15293\
        );

    \I__2262\ : Span12Mux_v
    port map (
            O => \N__15296\,
            I => \N__15290\
        );

    \I__2261\ : Span4Mux_h
    port map (
            O => \N__15293\,
            I => \N__15287\
        );

    \I__2260\ : Odrv12
    port map (
            O => \N__15290\,
            I => \this_vga_signals.vvisibility\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__15287\,
            I => \this_vga_signals.vvisibility\
        );

    \I__2258\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15279\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__15279\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_0\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__15276\,
            I => \this_ppu.N_1195_0_1_cascade_\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__15273\,
            I => \N__15269\
        );

    \I__2254\ : InMux
    port map (
            O => \N__15272\,
            I => \N__15264\
        );

    \I__2253\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15264\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__15264\,
            I => \N__15260\
        );

    \I__2251\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15257\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__15260\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__15257\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__2248\ : InMux
    port map (
            O => \N__15252\,
            I => \N__15249\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__15249\,
            I => \N__15246\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__15246\,
            I => \N__15242\
        );

    \I__2245\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15239\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__15242\,
            I => \this_vga_signals.vaddress_c3_0\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__15239\,
            I => \this_vga_signals.vaddress_c3_0\
        );

    \I__2242\ : InMux
    port map (
            O => \N__15234\,
            I => \N__15229\
        );

    \I__2241\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15224\
        );

    \I__2240\ : InMux
    port map (
            O => \N__15232\,
            I => \N__15224\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__15229\,
            I => \N__15220\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__15224\,
            I => \N__15217\
        );

    \I__2237\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15213\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__15220\,
            I => \N__15209\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__15217\,
            I => \N__15206\
        );

    \I__2234\ : InMux
    port map (
            O => \N__15216\,
            I => \N__15203\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__15213\,
            I => \N__15200\
        );

    \I__2232\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15197\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__15209\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__15206\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__15203\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__15200\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__15197\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__15186\,
            I => \N__15183\
        );

    \I__2225\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15179\
        );

    \I__2224\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15174\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__15179\,
            I => \N__15171\
        );

    \I__2222\ : InMux
    port map (
            O => \N__15178\,
            I => \N__15166\
        );

    \I__2221\ : InMux
    port map (
            O => \N__15177\,
            I => \N__15166\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__15174\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__15171\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__15166\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__2217\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15156\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__15156\,
            I => \N__15153\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__15153\,
            I => \N__15150\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__15150\,
            I => \this_vga_signals.if_m8_0_a3_1_1_1\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__15147\,
            I => \N__15143\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__15146\,
            I => \N__15138\
        );

    \I__2211\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15135\
        );

    \I__2210\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15132\
        );

    \I__2209\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15127\
        );

    \I__2208\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15127\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__15135\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__15132\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__15127\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__2204\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15117\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__15117\,
            I => \this_vga_signals.g2\
        );

    \I__2202\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15111\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__15111\,
            I => \N__15107\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__15110\,
            I => \N__15101\
        );

    \I__2199\ : Span4Mux_h
    port map (
            O => \N__15107\,
            I => \N__15096\
        );

    \I__2198\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15093\
        );

    \I__2197\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15088\
        );

    \I__2196\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15088\
        );

    \I__2195\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15085\
        );

    \I__2194\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15080\
        );

    \I__2193\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15080\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__15096\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__15093\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__15088\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__15085\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__15080\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__15069\,
            I => \N__15066\
        );

    \I__2186\ : InMux
    port map (
            O => \N__15066\,
            I => \N__15063\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__15063\,
            I => \this_vga_signals.g1_3\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__15060\,
            I => \N__15057\
        );

    \I__2183\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15054\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__15054\,
            I => \N__15051\
        );

    \I__2181\ : Span4Mux_h
    port map (
            O => \N__15051\,
            I => \N__15044\
        );

    \I__2180\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15041\
        );

    \I__2179\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15038\
        );

    \I__2178\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15033\
        );

    \I__2177\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15033\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__15044\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__15041\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__15038\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__15033\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__2172\ : InMux
    port map (
            O => \N__15024\,
            I => \N__15020\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__15023\,
            I => \N__15013\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__15020\,
            I => \N__15010\
        );

    \I__2169\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15005\
        );

    \I__2168\ : InMux
    port map (
            O => \N__15018\,
            I => \N__15000\
        );

    \I__2167\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15000\
        );

    \I__2166\ : InMux
    port map (
            O => \N__15016\,
            I => \N__14997\
        );

    \I__2165\ : InMux
    port map (
            O => \N__15013\,
            I => \N__14994\
        );

    \I__2164\ : Span4Mux_h
    port map (
            O => \N__15010\,
            I => \N__14991\
        );

    \I__2163\ : InMux
    port map (
            O => \N__15009\,
            I => \N__14988\
        );

    \I__2162\ : InMux
    port map (
            O => \N__15008\,
            I => \N__14985\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__15005\,
            I => \N__14980\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__15000\,
            I => \N__14980\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__14997\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__14994\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__14991\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__14988\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__14985\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__14980\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__14967\,
            I => \N__14962\
        );

    \I__2152\ : InMux
    port map (
            O => \N__14966\,
            I => \N__14953\
        );

    \I__2151\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14946\
        );

    \I__2150\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14946\
        );

    \I__2149\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14946\
        );

    \I__2148\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14943\
        );

    \I__2147\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14940\
        );

    \I__2146\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14937\
        );

    \I__2145\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14934\
        );

    \I__2144\ : InMux
    port map (
            O => \N__14956\,
            I => \N__14931\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__14953\,
            I => \N__14926\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__14946\,
            I => \N__14921\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__14943\,
            I => \N__14921\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__14940\,
            I => \N__14916\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__14937\,
            I => \N__14909\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__14934\,
            I => \N__14909\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__14931\,
            I => \N__14909\
        );

    \I__2136\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14906\
        );

    \I__2135\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14902\
        );

    \I__2134\ : Span4Mux_h
    port map (
            O => \N__14926\,
            I => \N__14897\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__14921\,
            I => \N__14897\
        );

    \I__2132\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14894\
        );

    \I__2131\ : InMux
    port map (
            O => \N__14919\,
            I => \N__14891\
        );

    \I__2130\ : Span4Mux_v
    port map (
            O => \N__14916\,
            I => \N__14886\
        );

    \I__2129\ : Span4Mux_v
    port map (
            O => \N__14909\,
            I => \N__14886\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__14906\,
            I => \N__14883\
        );

    \I__2127\ : InMux
    port map (
            O => \N__14905\,
            I => \N__14880\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__14902\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__14897\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__14894\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__14891\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__14886\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__14883\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__14880\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2119\ : InMux
    port map (
            O => \N__14865\,
            I => \N__14862\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__14862\,
            I => \N__14859\
        );

    \I__2117\ : Span4Mux_h
    port map (
            O => \N__14859\,
            I => \N__14856\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__14856\,
            I => \this_vga_signals.if_m2\
        );

    \I__2115\ : SRMux
    port map (
            O => \N__14853\,
            I => \N__14850\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__14850\,
            I => \N__14845\
        );

    \I__2113\ : SRMux
    port map (
            O => \N__14849\,
            I => \N__14842\
        );

    \I__2112\ : SRMux
    port map (
            O => \N__14848\,
            I => \N__14839\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__14845\,
            I => \N__14835\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__14842\,
            I => \N__14832\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__14839\,
            I => \N__14829\
        );

    \I__2108\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14826\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__14835\,
            I => \this_vga_signals.N_1098_1\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__14832\,
            I => \this_vga_signals.N_1098_1\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__14829\,
            I => \this_vga_signals.N_1098_1\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__14826\,
            I => \this_vga_signals.N_1098_1\
        );

    \I__2103\ : InMux
    port map (
            O => \N__14817\,
            I => \N__14814\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__14814\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__14811\,
            I => \N__14808\
        );

    \I__2100\ : InMux
    port map (
            O => \N__14808\,
            I => \N__14802\
        );

    \I__2099\ : InMux
    port map (
            O => \N__14807\,
            I => \N__14795\
        );

    \I__2098\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14795\
        );

    \I__2097\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14795\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__14802\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__14795\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__2094\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14787\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__14787\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_N_2L1\
        );

    \I__2092\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14779\
        );

    \I__2091\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14774\
        );

    \I__2090\ : InMux
    port map (
            O => \N__14782\,
            I => \N__14774\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__14779\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__14774\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__14769\,
            I => \this_vga_signals.SUM_2_i_1_2_3_cascade_\
        );

    \I__2086\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14762\
        );

    \I__2085\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14759\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__14762\,
            I => \this_vga_signals.SUM_2_i_1_1_3\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__14759\,
            I => \this_vga_signals.SUM_2_i_1_1_3\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__14754\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_x0_cascade_\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__14751\,
            I => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\
        );

    \I__2080\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14741\
        );

    \I__2079\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14736\
        );

    \I__2078\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14736\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__14745\,
            I => \N__14733\
        );

    \I__2076\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14729\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__14741\,
            I => \N__14724\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__14736\,
            I => \N__14724\
        );

    \I__2073\ : InMux
    port map (
            O => \N__14733\,
            I => \N__14721\
        );

    \I__2072\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14718\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__14729\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__14724\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__14721\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__14718\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__14709\,
            I => \N__14704\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__14708\,
            I => \N__14700\
        );

    \I__2065\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14697\
        );

    \I__2064\ : InMux
    port map (
            O => \N__14704\,
            I => \N__14694\
        );

    \I__2063\ : InMux
    port map (
            O => \N__14703\,
            I => \N__14689\
        );

    \I__2062\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14689\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__14697\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__14694\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__14689\,
            I => \this_vga_signals.mult1_un54_sum_axb2_i\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__14682\,
            I => \N__14679\
        );

    \I__2057\ : InMux
    port map (
            O => \N__14679\,
            I => \N__14673\
        );

    \I__2056\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14673\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__14673\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_N_2L1\
        );

    \I__2054\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14667\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__14667\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_x1\
        );

    \I__2052\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14655\
        );

    \I__2051\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14650\
        );

    \I__2050\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14650\
        );

    \I__2049\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14647\
        );

    \I__2048\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14640\
        );

    \I__2047\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14640\
        );

    \I__2046\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14640\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__14655\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__14650\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__14647\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__14640\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__2041\ : InMux
    port map (
            O => \N__14631\,
            I => \N__14628\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__14628\,
            I => \N__14625\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__14625\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_0\
        );

    \I__2038\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14614\
        );

    \I__2037\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14611\
        );

    \I__2036\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14607\
        );

    \I__2035\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14604\
        );

    \I__2034\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14599\
        );

    \I__2033\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14599\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__14614\,
            I => \N__14594\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__14611\,
            I => \N__14594\
        );

    \I__2030\ : InMux
    port map (
            O => \N__14610\,
            I => \N__14591\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__14607\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__14604\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__14599\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__14594\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__14591\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__2024\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14573\
        );

    \I__2023\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14573\
        );

    \I__2022\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14565\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__14573\,
            I => \N__14562\
        );

    \I__2020\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14555\
        );

    \I__2019\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14555\
        );

    \I__2018\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14555\
        );

    \I__2017\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14550\
        );

    \I__2016\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14550\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__14565\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__14562\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__14555\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__14550\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__14541\,
            I => \this_vga_signals.g2_0_a2_5Z0Z_1_cascade_\
        );

    \I__2010\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14535\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__14535\,
            I => \this_vga_signals.g2_0_a2_2\
        );

    \I__2008\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14529\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__14529\,
            I => \N__14526\
        );

    \I__2006\ : Span4Mux_h
    port map (
            O => \N__14526\,
            I => \N__14523\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__14523\,
            I => \this_vga_signals.g2_0_a2_5\
        );

    \I__2004\ : CEMux
    port map (
            O => \N__14520\,
            I => \N__14517\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__14517\,
            I => \N__14514\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__14514\,
            I => \this_vga_signals.N_852_1\
        );

    \I__2001\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14508\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__14508\,
            I => \N__14502\
        );

    \I__1999\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14495\
        );

    \I__1998\ : InMux
    port map (
            O => \N__14506\,
            I => \N__14495\
        );

    \I__1997\ : InMux
    port map (
            O => \N__14505\,
            I => \N__14492\
        );

    \I__1996\ : Span12Mux_s11_h
    port map (
            O => \N__14502\,
            I => \N__14489\
        );

    \I__1995\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14484\
        );

    \I__1994\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14484\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__14495\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__14492\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1991\ : Odrv12
    port map (
            O => \N__14489\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__14484\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1989\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14472\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__14472\,
            I => \this_vga_signals.un2_hsynclt6_0\
        );

    \I__1987\ : InMux
    port map (
            O => \N__14469\,
            I => \N__14466\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__14466\,
            I => \N__14456\
        );

    \I__1985\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14451\
        );

    \I__1984\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14451\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__14463\,
            I => \N__14445\
        );

    \I__1982\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14442\
        );

    \I__1981\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14439\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__14460\,
            I => \N__14435\
        );

    \I__1979\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14432\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__14456\,
            I => \N__14426\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__14451\,
            I => \N__14426\
        );

    \I__1976\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14423\
        );

    \I__1975\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14416\
        );

    \I__1974\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14416\
        );

    \I__1973\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14416\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__14442\,
            I => \N__14413\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__14439\,
            I => \N__14396\
        );

    \I__1970\ : InMux
    port map (
            O => \N__14438\,
            I => \N__14393\
        );

    \I__1969\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14390\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__14432\,
            I => \N__14387\
        );

    \I__1967\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14384\
        );

    \I__1966\ : Span4Mux_v
    port map (
            O => \N__14426\,
            I => \N__14379\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__14423\,
            I => \N__14379\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__14416\,
            I => \N__14374\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__14413\,
            I => \N__14374\
        );

    \I__1962\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14367\
        );

    \I__1961\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14367\
        );

    \I__1960\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14367\
        );

    \I__1959\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14356\
        );

    \I__1958\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14356\
        );

    \I__1957\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14356\
        );

    \I__1956\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14356\
        );

    \I__1955\ : InMux
    port map (
            O => \N__14405\,
            I => \N__14356\
        );

    \I__1954\ : InMux
    port map (
            O => \N__14404\,
            I => \N__14343\
        );

    \I__1953\ : InMux
    port map (
            O => \N__14403\,
            I => \N__14343\
        );

    \I__1952\ : InMux
    port map (
            O => \N__14402\,
            I => \N__14343\
        );

    \I__1951\ : InMux
    port map (
            O => \N__14401\,
            I => \N__14343\
        );

    \I__1950\ : InMux
    port map (
            O => \N__14400\,
            I => \N__14343\
        );

    \I__1949\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14343\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__14396\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__14393\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__14390\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__14387\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__14384\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__14379\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__14374\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__14367\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__14356\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__14343\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1938\ : InMux
    port map (
            O => \N__14322\,
            I => \N__14319\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__14319\,
            I => \N__14316\
        );

    \I__1936\ : Span4Mux_h
    port map (
            O => \N__14316\,
            I => \N__14313\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__14313\,
            I => \this_vga_signals.un2_hsynclt7\
        );

    \I__1934\ : InMux
    port map (
            O => \N__14310\,
            I => \N__14306\
        );

    \I__1933\ : InMux
    port map (
            O => \N__14309\,
            I => \N__14303\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__14306\,
            I => \this_vga_signals.un2_hsynclto3_0\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__14303\,
            I => \this_vga_signals.un2_hsynclto3_0\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__14298\,
            I => \N__14290\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__14297\,
            I => \N__14285\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__14296\,
            I => \N__14282\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__14295\,
            I => \N__14279\
        );

    \I__1926\ : InMux
    port map (
            O => \N__14294\,
            I => \N__14271\
        );

    \I__1925\ : InMux
    port map (
            O => \N__14293\,
            I => \N__14271\
        );

    \I__1924\ : InMux
    port map (
            O => \N__14290\,
            I => \N__14271\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__14289\,
            I => \N__14267\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__14288\,
            I => \N__14263\
        );

    \I__1921\ : InMux
    port map (
            O => \N__14285\,
            I => \N__14258\
        );

    \I__1920\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14255\
        );

    \I__1919\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14249\
        );

    \I__1918\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14249\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__14271\,
            I => \N__14245\
        );

    \I__1916\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14242\
        );

    \I__1915\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14239\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__14266\,
            I => \N__14234\
        );

    \I__1913\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14229\
        );

    \I__1912\ : InMux
    port map (
            O => \N__14262\,
            I => \N__14229\
        );

    \I__1911\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14226\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__14258\,
            I => \N__14221\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__14255\,
            I => \N__14221\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__14254\,
            I => \N__14212\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__14249\,
            I => \N__14206\
        );

    \I__1906\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14203\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__14245\,
            I => \N__14196\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__14242\,
            I => \N__14196\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__14239\,
            I => \N__14196\
        );

    \I__1902\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14189\
        );

    \I__1901\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14189\
        );

    \I__1900\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14189\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__14229\,
            I => \N__14186\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__14226\,
            I => \N__14181\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__14221\,
            I => \N__14181\
        );

    \I__1896\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14170\
        );

    \I__1895\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14170\
        );

    \I__1894\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14170\
        );

    \I__1893\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14170\
        );

    \I__1892\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14170\
        );

    \I__1891\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14161\
        );

    \I__1890\ : InMux
    port map (
            O => \N__14212\,
            I => \N__14161\
        );

    \I__1889\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14161\
        );

    \I__1888\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14161\
        );

    \I__1887\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14158\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__14206\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__14203\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__14196\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__14189\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__14186\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__14181\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__14170\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__14161\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__14158\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__14139\,
            I => \N__14134\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__14138\,
            I => \N__14129\
        );

    \I__1875\ : InMux
    port map (
            O => \N__14137\,
            I => \N__14118\
        );

    \I__1874\ : InMux
    port map (
            O => \N__14134\,
            I => \N__14118\
        );

    \I__1873\ : InMux
    port map (
            O => \N__14133\,
            I => \N__14115\
        );

    \I__1872\ : InMux
    port map (
            O => \N__14132\,
            I => \N__14108\
        );

    \I__1871\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14108\
        );

    \I__1870\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14108\
        );

    \I__1869\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14105\
        );

    \I__1868\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14100\
        );

    \I__1867\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14100\
        );

    \I__1866\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14095\
        );

    \I__1865\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14095\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__14118\,
            I => \N__14091\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__14115\,
            I => \N__14083\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__14108\,
            I => \N__14080\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__14105\,
            I => \N__14073\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__14100\,
            I => \N__14073\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__14095\,
            I => \N__14073\
        );

    \I__1858\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14070\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__14091\,
            I => \N__14067\
        );

    \I__1856\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14060\
        );

    \I__1855\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14060\
        );

    \I__1854\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14060\
        );

    \I__1853\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14050\
        );

    \I__1852\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14047\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__14083\,
            I => \N__14042\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__14080\,
            I => \N__14042\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__14073\,
            I => \N__14039\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__14070\,
            I => \N__14036\
        );

    \I__1847\ : Sp12to4
    port map (
            O => \N__14067\,
            I => \N__14031\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__14060\,
            I => \N__14031\
        );

    \I__1845\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14026\
        );

    \I__1844\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14026\
        );

    \I__1843\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14019\
        );

    \I__1842\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14019\
        );

    \I__1841\ : InMux
    port map (
            O => \N__14055\,
            I => \N__14019\
        );

    \I__1840\ : InMux
    port map (
            O => \N__14054\,
            I => \N__14016\
        );

    \I__1839\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14013\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__14050\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__14047\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__14042\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__14039\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__14036\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1833\ : Odrv12
    port map (
            O => \N__14031\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__14026\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__14019\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__14016\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__14013\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1828\ : InMux
    port map (
            O => \N__13992\,
            I => \N__13989\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__13989\,
            I => \this_vga_signals.un4_hsynclto7_0\
        );

    \I__1826\ : InMux
    port map (
            O => \N__13986\,
            I => \N__13983\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__13983\,
            I => \N__13980\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__13980\,
            I => \N__13977\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__13977\,
            I => \M_this_map_ram_write_data_1\
        );

    \I__1822\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13971\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__13971\,
            I => \this_vga_signals.SUM_2_i_1_1_1_3\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__13968\,
            I => \this_vga_signals.N_1_3_1_cascade_\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__13965\,
            I => \N__13962\
        );

    \I__1818\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13959\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__13959\,
            I => \this_vga_signals.SUM_2_i_1_2_3\
        );

    \I__1816\ : IoInMux
    port map (
            O => \N__13956\,
            I => \N__13953\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__13953\,
            I => \N__13950\
        );

    \I__1814\ : Span4Mux_s3_v
    port map (
            O => \N__13950\,
            I => \N__13947\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__13947\,
            I => \N__13944\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__13944\,
            I => \N__13941\
        );

    \I__1811\ : Sp12to4
    port map (
            O => \N__13941\,
            I => \N__13938\
        );

    \I__1810\ : Span12Mux_v
    port map (
            O => \N__13938\,
            I => \N__13935\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__13935\,
            I => this_vga_signals_vsync_1_i
        );

    \I__1808\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13929\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__13929\,
            I => \this_vga_signals.un2_vsynclt8\
        );

    \I__1806\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13923\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__13923\,
            I => \N__13917\
        );

    \I__1804\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13914\
        );

    \I__1803\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13909\
        );

    \I__1802\ : InMux
    port map (
            O => \N__13920\,
            I => \N__13909\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__13917\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__13914\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__13909\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d\
        );

    \I__1798\ : InMux
    port map (
            O => \N__13902\,
            I => \N__13898\
        );

    \I__1797\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13895\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__13898\,
            I => \this_vga_signals.mult1_un54_sum_0_3\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__13895\,
            I => \this_vga_signals.mult1_un54_sum_0_3\
        );

    \I__1794\ : InMux
    port map (
            O => \N__13890\,
            I => \N__13887\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__13887\,
            I => \N__13881\
        );

    \I__1792\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13877\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__13885\,
            I => \N__13874\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__13884\,
            I => \N__13871\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__13881\,
            I => \N__13864\
        );

    \I__1788\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13861\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__13877\,
            I => \N__13858\
        );

    \I__1786\ : InMux
    port map (
            O => \N__13874\,
            I => \N__13855\
        );

    \I__1785\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13848\
        );

    \I__1784\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13848\
        );

    \I__1783\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13848\
        );

    \I__1782\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13840\
        );

    \I__1781\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13837\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__13864\,
            I => \N__13832\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__13861\,
            I => \N__13832\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__13858\,
            I => \N__13825\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__13855\,
            I => \N__13825\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__13848\,
            I => \N__13825\
        );

    \I__1775\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13816\
        );

    \I__1774\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13816\
        );

    \I__1773\ : InMux
    port map (
            O => \N__13845\,
            I => \N__13816\
        );

    \I__1772\ : InMux
    port map (
            O => \N__13844\,
            I => \N__13816\
        );

    \I__1771\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13813\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__13840\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__13837\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__13832\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__13825\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__13816\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__13813\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__13800\,
            I => \N__13788\
        );

    \I__1763\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13778\
        );

    \I__1762\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13778\
        );

    \I__1761\ : InMux
    port map (
            O => \N__13797\,
            I => \N__13769\
        );

    \I__1760\ : InMux
    port map (
            O => \N__13796\,
            I => \N__13769\
        );

    \I__1759\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13769\
        );

    \I__1758\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13769\
        );

    \I__1757\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13758\
        );

    \I__1756\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13758\
        );

    \I__1755\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13758\
        );

    \I__1754\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13758\
        );

    \I__1753\ : InMux
    port map (
            O => \N__13787\,
            I => \N__13753\
        );

    \I__1752\ : InMux
    port map (
            O => \N__13786\,
            I => \N__13753\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__13785\,
            I => \N__13749\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__13784\,
            I => \N__13744\
        );

    \I__1749\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13741\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__13778\,
            I => \N__13736\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__13769\,
            I => \N__13736\
        );

    \I__1746\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13731\
        );

    \I__1745\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13731\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__13758\,
            I => \N__13728\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__13753\,
            I => \N__13725\
        );

    \I__1742\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13721\
        );

    \I__1741\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13718\
        );

    \I__1740\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13715\
        );

    \I__1739\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13710\
        );

    \I__1738\ : InMux
    port map (
            O => \N__13744\,
            I => \N__13710\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__13741\,
            I => \N__13705\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__13736\,
            I => \N__13705\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__13731\,
            I => \N__13702\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__13728\,
            I => \N__13697\
        );

    \I__1733\ : Span4Mux_h
    port map (
            O => \N__13725\,
            I => \N__13697\
        );

    \I__1732\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13694\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__13721\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__13718\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__13715\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__13710\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__13705\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__13702\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__13697\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__13694\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__13677\,
            I => \this_vga_signals.un2_hsynclto3_0_cascade_\
        );

    \I__1722\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13671\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__13671\,
            I => \this_vga_signals.M_hcounter_d7lto7_1\
        );

    \I__1720\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13661\
        );

    \I__1719\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13661\
        );

    \I__1718\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13656\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__13661\,
            I => \N__13652\
        );

    \I__1716\ : InMux
    port map (
            O => \N__13660\,
            I => \N__13649\
        );

    \I__1715\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13646\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__13656\,
            I => \N__13640\
        );

    \I__1713\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13637\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__13652\,
            I => \N__13632\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__13649\,
            I => \N__13632\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__13646\,
            I => \N__13624\
        );

    \I__1709\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13621\
        );

    \I__1708\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13616\
        );

    \I__1707\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13616\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__13640\,
            I => \N__13609\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__13637\,
            I => \N__13609\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__13632\,
            I => \N__13609\
        );

    \I__1703\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13606\
        );

    \I__1702\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13597\
        );

    \I__1701\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13597\
        );

    \I__1700\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13597\
        );

    \I__1699\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13597\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__13624\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__13621\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__13616\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__13609\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__13606\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__13597\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__13584\,
            I => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\
        );

    \I__1691\ : InMux
    port map (
            O => \N__13581\,
            I => \N__13574\
        );

    \I__1690\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13574\
        );

    \I__1689\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13571\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__13574\,
            I => \N__13565\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__13571\,
            I => \N__13556\
        );

    \I__1686\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13549\
        );

    \I__1685\ : InMux
    port map (
            O => \N__13569\,
            I => \N__13549\
        );

    \I__1684\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13549\
        );

    \I__1683\ : Span4Mux_h
    port map (
            O => \N__13565\,
            I => \N__13546\
        );

    \I__1682\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13543\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__13563\,
            I => \N__13539\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__13562\,
            I => \N__13536\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__13561\,
            I => \N__13533\
        );

    \I__1678\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13529\
        );

    \I__1677\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13526\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__13556\,
            I => \N__13521\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13521\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__13546\,
            I => \N__13516\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__13543\,
            I => \N__13516\
        );

    \I__1672\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13513\
        );

    \I__1671\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13504\
        );

    \I__1670\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13504\
        );

    \I__1669\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13504\
        );

    \I__1668\ : InMux
    port map (
            O => \N__13532\,
            I => \N__13504\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__13529\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__13526\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__13521\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__13516\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__13513\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__13504\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__13491\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_cascade_\
        );

    \I__1660\ : InMux
    port map (
            O => \N__13488\,
            I => \N__13484\
        );

    \I__1659\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13481\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__13484\,
            I => \N__13478\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__13481\,
            I => \this_vga_signals.g0_0_0_a2_0\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__13478\,
            I => \this_vga_signals.g0_0_0_a2_0\
        );

    \I__1655\ : InMux
    port map (
            O => \N__13473\,
            I => \N__13467\
        );

    \I__1654\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13462\
        );

    \I__1653\ : InMux
    port map (
            O => \N__13471\,
            I => \N__13462\
        );

    \I__1652\ : InMux
    port map (
            O => \N__13470\,
            I => \N__13459\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__13467\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__13462\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__13459\,
            I => \this_vga_signals.mult1_un47_sum_c3\
        );

    \I__1648\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13446\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__13451\,
            I => \N__13438\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__13450\,
            I => \N__13432\
        );

    \I__1645\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13429\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__13446\,
            I => \N__13426\
        );

    \I__1643\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13423\
        );

    \I__1642\ : InMux
    port map (
            O => \N__13444\,
            I => \N__13420\
        );

    \I__1641\ : InMux
    port map (
            O => \N__13443\,
            I => \N__13417\
        );

    \I__1640\ : InMux
    port map (
            O => \N__13442\,
            I => \N__13408\
        );

    \I__1639\ : InMux
    port map (
            O => \N__13441\,
            I => \N__13408\
        );

    \I__1638\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13408\
        );

    \I__1637\ : InMux
    port map (
            O => \N__13437\,
            I => \N__13408\
        );

    \I__1636\ : InMux
    port map (
            O => \N__13436\,
            I => \N__13401\
        );

    \I__1635\ : InMux
    port map (
            O => \N__13435\,
            I => \N__13401\
        );

    \I__1634\ : InMux
    port map (
            O => \N__13432\,
            I => \N__13401\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__13429\,
            I => \N__13398\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__13426\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__13423\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__13420\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__13417\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__13408\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__13401\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__13398\,
            I => \this_vga_signals.mult1_un61_sum_c3\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__13383\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\
        );

    \I__1624\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13371\
        );

    \I__1623\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13368\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__13378\,
            I => \N__13360\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__13377\,
            I => \N__13356\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__13376\,
            I => \N__13353\
        );

    \I__1619\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13350\
        );

    \I__1618\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13347\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__13371\,
            I => \N__13342\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__13368\,
            I => \N__13342\
        );

    \I__1615\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13335\
        );

    \I__1614\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13335\
        );

    \I__1613\ : InMux
    port map (
            O => \N__13365\,
            I => \N__13335\
        );

    \I__1612\ : InMux
    port map (
            O => \N__13364\,
            I => \N__13332\
        );

    \I__1611\ : InMux
    port map (
            O => \N__13363\,
            I => \N__13329\
        );

    \I__1610\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13322\
        );

    \I__1609\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13322\
        );

    \I__1608\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13322\
        );

    \I__1607\ : InMux
    port map (
            O => \N__13353\,
            I => \N__13319\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__13350\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__13347\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__13342\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13335\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__13332\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__13329\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__13322\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__13319\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661\
        );

    \I__1598\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13299\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__13299\,
            I => \this_vga_signals.g0_i_x4_0_a3_2\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__13296\,
            I => \N__13293\
        );

    \I__1595\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13290\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__13290\,
            I => \N__13287\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__13287\,
            I => \this_vga_signals.vaddress_0_6\
        );

    \I__1592\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13281\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__13281\,
            I => \this_vga_signals.g0_i_x4_0_a3_0\
        );

    \I__1590\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13275\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__13275\,
            I => \this_vga_signals.vsync_1_3\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__13272\,
            I => \this_vga_signals.vsync_1_2_cascade_\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__13269\,
            I => \this_vga_signals.mult1_un68_sum_axb1_661_cascade_\
        );

    \I__1586\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13263\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__13263\,
            I => \this_vga_signals.g0_2_0_a2_1\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__13260\,
            I => \this_vga_signals.if_N_5_cascade_\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__13257\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__13254\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_1_cascade_\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__13251\,
            I => \this_vga_signals.mult1_un61_sum_c3_cascade_\
        );

    \I__1580\ : InMux
    port map (
            O => \N__13248\,
            I => \N__13242\
        );

    \I__1579\ : InMux
    port map (
            O => \N__13247\,
            I => \N__13242\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__13242\,
            I => \N__13239\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__13239\,
            I => \this_vga_signals.N_4_0_1_0\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__13236\,
            I => \this_vga_signals.mult1_un47_sum_c3_cascade_\
        );

    \I__1575\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13230\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__13230\,
            I => \this_vga_signals.g1_2\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__13227\,
            I => \this_vga_signals.SUM_3_0_cascade_\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__13224\,
            I => \N__13221\
        );

    \I__1571\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13218\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__13218\,
            I => \this_vga_signals.mult1_un61_sum_axb1_0\
        );

    \I__1569\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13212\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__13212\,
            I => \N__13209\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__13209\,
            I => \N__13206\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__13206\,
            I => \M_this_map_ram_write_data_4\
        );

    \I__1565\ : InMux
    port map (
            O => \N__13203\,
            I => \N__13200\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__13200\,
            I => \this_vga_signals.mult1_un40_sum_axb1_i_0\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__13197\,
            I => \this_vga_signals.N_18_cascade_\
        );

    \I__1562\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__13191\,
            I => \this_vga_signals.g1_0_0_1\
        );

    \I__1560\ : InMux
    port map (
            O => \N__13188\,
            I => \N__13185\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__13185\,
            I => \this_vga_signals.vaddress_1_6\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__13182\,
            I => \this_vga_signals.N_6_cascade_\
        );

    \I__1557\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13173\
        );

    \I__1556\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13173\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__13173\,
            I => \this_vga_signals.g1_1_1\
        );

    \I__1554\ : InMux
    port map (
            O => \N__13170\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1553\ : InMux
    port map (
            O => \N__13167\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1552\ : InMux
    port map (
            O => \N__13164\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1551\ : InMux
    port map (
            O => \N__13161\,
            I => \bfn_11_14_0_\
        );

    \I__1550\ : InMux
    port map (
            O => \N__13158\,
            I => \N__13155\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__13155\,
            I => \this_vga_signals.un4_hsynclt9\
        );

    \I__1548\ : InMux
    port map (
            O => \N__13152\,
            I => \N__13147\
        );

    \I__1547\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13144\
        );

    \I__1546\ : InMux
    port map (
            O => \N__13150\,
            I => \N__13141\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__13147\,
            I => \N__13138\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__13144\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__13141\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__13138\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__13131\,
            I => \N__13127\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__13130\,
            I => \N__13123\
        );

    \I__1539\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13120\
        );

    \I__1538\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13115\
        );

    \I__1537\ : InMux
    port map (
            O => \N__13123\,
            I => \N__13115\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__13120\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__13115\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__13110\,
            I => \this_vga_signals.M_pcounter_q_3_1_cascade_\
        );

    \I__1533\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13101\
        );

    \I__1532\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13101\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__13101\,
            I => \N__13098\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__13098\,
            I => \N_3_0\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__13095\,
            I => \N_3_0_cascade_\
        );

    \I__1528\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13089\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__13089\,
            I => \N__13083\
        );

    \I__1526\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13078\
        );

    \I__1525\ : InMux
    port map (
            O => \N__13087\,
            I => \N__13078\
        );

    \I__1524\ : InMux
    port map (
            O => \N__13086\,
            I => \N__13075\
        );

    \I__1523\ : Span4Mux_h
    port map (
            O => \N__13083\,
            I => \N__13072\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__13078\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__13075\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__13072\,
            I => \this_vga_signals.M_pcounter_q_i_3_1\
        );

    \I__1519\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13062\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__13062\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_1\
        );

    \I__1517\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13056\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__13056\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_a0_0\
        );

    \I__1515\ : InMux
    port map (
            O => \N__13053\,
            I => \N__13046\
        );

    \I__1514\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13042\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__13051\,
            I => \N__13038\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__13050\,
            I => \N__13033\
        );

    \I__1511\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13027\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__13046\,
            I => \N__13024\
        );

    \I__1509\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13021\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__13042\,
            I => \N__13018\
        );

    \I__1507\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13015\
        );

    \I__1506\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13008\
        );

    \I__1505\ : InMux
    port map (
            O => \N__13037\,
            I => \N__13008\
        );

    \I__1504\ : InMux
    port map (
            O => \N__13036\,
            I => \N__13008\
        );

    \I__1503\ : InMux
    port map (
            O => \N__13033\,
            I => \N__12999\
        );

    \I__1502\ : InMux
    port map (
            O => \N__13032\,
            I => \N__12999\
        );

    \I__1501\ : InMux
    port map (
            O => \N__13031\,
            I => \N__12999\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13030\,
            I => \N__12999\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__13027\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__13024\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__13021\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__13018\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__13015\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__13008\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__12999\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__12984\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz_cascade_\
        );

    \I__1491\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12976\
        );

    \I__1490\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12970\
        );

    \I__1489\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12962\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__12976\,
            I => \N__12959\
        );

    \I__1487\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12956\
        );

    \I__1486\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12951\
        );

    \I__1485\ : InMux
    port map (
            O => \N__12973\,
            I => \N__12951\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__12970\,
            I => \N__12948\
        );

    \I__1483\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12945\
        );

    \I__1482\ : InMux
    port map (
            O => \N__12968\,
            I => \N__12936\
        );

    \I__1481\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12936\
        );

    \I__1480\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12936\
        );

    \I__1479\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12936\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__12962\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__12959\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__12956\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__12951\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__12948\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__12945\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__12936\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\
        );

    \I__1471\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12918\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__12918\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__1469\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12912\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__12912\,
            I => \this_vga_signals.if_N_6_0\
        );

    \I__1467\ : InMux
    port map (
            O => \N__12909\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1466\ : InMux
    port map (
            O => \N__12906\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1465\ : InMux
    port map (
            O => \N__12903\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1464\ : InMux
    port map (
            O => \N__12900\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1463\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12894\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__12894\,
            I => \this_vga_signals.g1_0\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__12891\,
            I => \this_vga_signals.g0_i_x4_2_0_0_1_cascade_\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__12888\,
            I => \N__12885\
        );

    \I__1459\ : InMux
    port map (
            O => \N__12885\,
            I => \N__12882\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__12882\,
            I => \this_vga_signals.g0_i_x4_0_0\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__12879\,
            I => \this_vga_signals.N_3_cascade_\
        );

    \I__1456\ : InMux
    port map (
            O => \N__12876\,
            I => \N__12873\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__12873\,
            I => \this_vga_signals.N_4_0_0\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__12870\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_0_cascade_\
        );

    \I__1453\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12864\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__12864\,
            I => \N__12861\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__12861\,
            I => \this_vga_signals.mult1_un75_sum_c2_0_0_0\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__12858\,
            I => \N__12855\
        );

    \I__1449\ : InMux
    port map (
            O => \N__12855\,
            I => \N__12852\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__12852\,
            I => \this_vga_signals.g0_2_1\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__12849\,
            I => \N__12844\
        );

    \I__1446\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12841\
        );

    \I__1445\ : InMux
    port map (
            O => \N__12847\,
            I => \N__12836\
        );

    \I__1444\ : InMux
    port map (
            O => \N__12844\,
            I => \N__12836\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__12841\,
            I => \this_vga_signals.N_5_0_0\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__12836\,
            I => \this_vga_signals.N_5_0_0\
        );

    \I__1441\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12828\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__12828\,
            I => \N__12825\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__12825\,
            I => \N__12822\
        );

    \I__1438\ : Span4Mux_v
    port map (
            O => \N__12822\,
            I => \N__12818\
        );

    \I__1437\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12815\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__12818\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__12815\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1434\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12807\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__12807\,
            I => \this_vga_signals.mult1_un68_sum_ac0_2\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__12804\,
            I => \this_vga_signals.mult1_un68_sum_ac0_2_cascade_\
        );

    \I__1431\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12798\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__12798\,
            I => \this_vga_signals.g1_0_3\
        );

    \I__1429\ : InMux
    port map (
            O => \N__12795\,
            I => \N__12792\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__12792\,
            I => \this_vga_signals.g0_2_0_a2\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__12789\,
            I => \N__12786\
        );

    \I__1426\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12780\
        );

    \I__1425\ : InMux
    port map (
            O => \N__12785\,
            I => \N__12780\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__12780\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__12777\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\
        );

    \I__1422\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12771\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__12771\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__1420\ : InMux
    port map (
            O => \N__12768\,
            I => \N__12765\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__12765\,
            I => \this_vga_signals.g0_1_2\
        );

    \I__1418\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12759\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__12759\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_x1\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__12756\,
            I => \this_vga_signals.g3_0_cascade_\
        );

    \I__1415\ : InMux
    port map (
            O => \N__12753\,
            I => \N__12750\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__12750\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_2\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__12747\,
            I => \this_vga_signals.g0_0_a2_0_0_cascade_\
        );

    \I__1412\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12741\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__12741\,
            I => \this_vga_signals.g1_0_a2_1\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__12738\,
            I => \N__12735\
        );

    \I__1409\ : InMux
    port map (
            O => \N__12735\,
            I => \N__12732\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__12732\,
            I => \this_vga_signals.vaddress_1_5\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__12729\,
            I => \N__12726\
        );

    \I__1406\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12723\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__12723\,
            I => \N__12720\
        );

    \I__1404\ : Span4Mux_h
    port map (
            O => \N__12720\,
            I => \N__12717\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__12717\,
            I => \this_vga_signals.mult1_un47_sum_c3_0_0\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__12714\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_x0_cascade_\
        );

    \I__1401\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12708\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__12708\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_ns\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__12705\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_ns_cascade_\
        );

    \I__1398\ : InMux
    port map (
            O => \N__12702\,
            I => \N__12699\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__12699\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\
        );

    \I__1396\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12693\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__12693\,
            I => \this_vga_signals.g0_i_x4_1\
        );

    \I__1394\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12687\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__12687\,
            I => \this_vga_signals.g0_i_x4_0_1\
        );

    \I__1392\ : InMux
    port map (
            O => \N__12684\,
            I => \N__12681\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__12681\,
            I => \this_vga_signals.mult1_un68_sum_axb1_0\
        );

    \I__1390\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12674\
        );

    \I__1389\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12670\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__12674\,
            I => \N__12666\
        );

    \I__1387\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12663\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__12670\,
            I => \N__12660\
        );

    \I__1385\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12657\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__12666\,
            I => \N__12641\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__12663\,
            I => \N__12641\
        );

    \I__1382\ : Span4Mux_v
    port map (
            O => \N__12660\,
            I => \N__12636\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__12657\,
            I => \N__12636\
        );

    \I__1380\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12631\
        );

    \I__1379\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12631\
        );

    \I__1378\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12624\
        );

    \I__1377\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12624\
        );

    \I__1376\ : InMux
    port map (
            O => \N__12652\,
            I => \N__12624\
        );

    \I__1375\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12619\
        );

    \I__1374\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12619\
        );

    \I__1373\ : InMux
    port map (
            O => \N__12649\,
            I => \N__12616\
        );

    \I__1372\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12609\
        );

    \I__1371\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12609\
        );

    \I__1370\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12609\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__12641\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__12636\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__12631\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__12624\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__12619\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__12616\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__12609\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1362\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12591\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__12591\,
            I => \N__12588\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__12588\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0\
        );

    \I__1359\ : InMux
    port map (
            O => \N__12585\,
            I => \N__12581\
        );

    \I__1358\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12578\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__12581\,
            I => \N__12573\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__12578\,
            I => \N__12573\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__12573\,
            I => \this_vga_signals.SUM_3_0_0\
        );

    \I__1354\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12566\
        );

    \I__1353\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12563\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__12566\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__12563\,
            I => \this_vga_signals.M_pcounter_q_i_3_0\
        );

    \I__1350\ : IoInMux
    port map (
            O => \N__12558\,
            I => \N__12555\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__12555\,
            I => \N__12552\
        );

    \I__1348\ : IoSpan4Mux
    port map (
            O => \N__12552\,
            I => \N__12549\
        );

    \I__1347\ : Span4Mux_s3_v
    port map (
            O => \N__12549\,
            I => \N__12546\
        );

    \I__1346\ : Sp12to4
    port map (
            O => \N__12546\,
            I => \N__12543\
        );

    \I__1345\ : Span12Mux_v
    port map (
            O => \N__12543\,
            I => \N__12540\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__12540\,
            I => this_vga_signals_hsync_1_i
        );

    \I__1343\ : IoInMux
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__12534\,
            I => \N__12531\
        );

    \I__1341\ : Span4Mux_s3_v
    port map (
            O => \N__12531\,
            I => \N__12528\
        );

    \I__1340\ : Sp12to4
    port map (
            O => \N__12528\,
            I => \N__12525\
        );

    \I__1339\ : Span12Mux_s11_h
    port map (
            O => \N__12525\,
            I => \N__12522\
        );

    \I__1338\ : Span12Mux_v
    port map (
            O => \N__12522\,
            I => \N__12519\
        );

    \I__1337\ : Odrv12
    port map (
            O => \N__12519\,
            I => this_vga_signals_hvisibility_i
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__12516\,
            I => \this_vga_signals.g3_0_1_cascade_\
        );

    \I__1335\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12510\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__12510\,
            I => \this_vga_signals.g3_0\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__12507\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\
        );

    \I__1332\ : InMux
    port map (
            O => \N__12504\,
            I => \N__12497\
        );

    \I__1331\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12490\
        );

    \I__1330\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12490\
        );

    \I__1329\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12490\
        );

    \I__1328\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12487\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__12497\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_1\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__12490\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_1\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__12487\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_3_1\
        );

    \I__1324\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12477\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__12477\,
            I => \this_vga_signals.N_6_1_0\
        );

    \I__1322\ : InMux
    port map (
            O => \N__12474\,
            I => \N__12471\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__12471\,
            I => \N__12468\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__12468\,
            I => \N__12464\
        );

    \I__1319\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12461\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__12464\,
            I => \this_vga_signals.N_234\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__12461\,
            I => \this_vga_signals.N_234\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \this_vga_signals.SUM_3_cascade_\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__12453\,
            I => \N__12450\
        );

    \I__1314\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12447\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__12447\,
            I => \this_vga_signals.g0_6_1\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__12444\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9_cascade_\
        );

    \I__1311\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12438\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__12438\,
            I => \this_vga_signals.mult1_un61_sum_axb1_1\
        );

    \I__1309\ : InMux
    port map (
            O => \N__12435\,
            I => \N__12432\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__12432\,
            I => \N__12429\
        );

    \I__1307\ : Span4Mux_h
    port map (
            O => \N__12429\,
            I => \N__12426\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__12426\,
            I => \this_vga_signals.g1_2_0_0\
        );

    \I__1305\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12420\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__12420\,
            I => \N__12415\
        );

    \I__1303\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12410\
        );

    \I__1302\ : InMux
    port map (
            O => \N__12418\,
            I => \N__12410\
        );

    \I__1301\ : Span4Mux_h
    port map (
            O => \N__12415\,
            I => \N__12405\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__12410\,
            I => \N__12405\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__12405\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__1298\ : InMux
    port map (
            O => \N__12402\,
            I => \N__12399\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__12399\,
            I => \this_vga_signals.g1_7\
        );

    \I__1296\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12393\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__12393\,
            I => \this_vga_signals.g0_i_x4_3_0\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__12390\,
            I => \this_vga_signals.mult1_un61_sum_axb1_3_0_cascade_\
        );

    \I__1293\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12384\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__12384\,
            I => \this_vga_signals.g1_1_0\
        );

    \I__1291\ : InMux
    port map (
            O => \N__12381\,
            I => \N__12378\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__12378\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_1\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__12375\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_\
        );

    \I__1288\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12369\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__12369\,
            I => \this_vga_signals.g1_0_1_0\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__12366\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__12363\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_3_cascade_\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__12360\,
            I => \N__12357\
        );

    \I__1283\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12354\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__12354\,
            I => \N__12348\
        );

    \I__1281\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12343\
        );

    \I__1280\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12343\
        );

    \I__1279\ : InMux
    port map (
            O => \N__12351\,
            I => \N__12340\
        );

    \I__1278\ : Odrv12
    port map (
            O => \N__12348\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__12343\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__12340\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__12333\,
            I => \N__12329\
        );

    \I__1274\ : InMux
    port map (
            O => \N__12332\,
            I => \N__12325\
        );

    \I__1273\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12320\
        );

    \I__1272\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12320\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__12325\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__12320\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0
        );

    \I__1269\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__12312\,
            I => \N__12309\
        );

    \I__1267\ : Span4Mux_h
    port map (
            O => \N__12309\,
            I => \N__12306\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__12306\,
            I => \this_vga_signals.d_N_3_1_i\
        );

    \I__1265\ : InMux
    port map (
            O => \N__12303\,
            I => \N__12300\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__12300\,
            I => \this_vga_signals.M_hcounter_q_RNIO08E8Z0Z_3\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__12297\,
            I => \N__12289\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__12296\,
            I => \N__12286\
        );

    \I__1261\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12282\
        );

    \I__1260\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12277\
        );

    \I__1259\ : InMux
    port map (
            O => \N__12293\,
            I => \N__12277\
        );

    \I__1258\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12268\
        );

    \I__1257\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12268\
        );

    \I__1256\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12268\
        );

    \I__1255\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12268\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__12282\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__12277\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__12268\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__12261\,
            I => \this_vga_signals.g1_0_1_cascade_\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__12258\,
            I => \this_vga_signals.g1_2_0_cascade_\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__12255\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_0_0_cascade_\
        );

    \I__1248\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12249\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__12249\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1_0_0_1\
        );

    \I__1246\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12243\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__12243\,
            I => \this_vga_signals.mult1_un89_sum_c3_1_0_0_1\
        );

    \I__1244\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12230\
        );

    \I__1243\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12221\
        );

    \I__1242\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12221\
        );

    \I__1241\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12221\
        );

    \I__1240\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12221\
        );

    \I__1239\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12218\
        );

    \I__1238\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12213\
        );

    \I__1237\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12213\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__12230\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__12221\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__12218\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__12213\,
            I => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0
        );

    \I__1232\ : InMux
    port map (
            O => \N__12204\,
            I => \N__12201\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__12201\,
            I => \this_vga_signals.N_4_2\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__12198\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__12195\,
            I => \N__12192\
        );

    \I__1228\ : InMux
    port map (
            O => \N__12192\,
            I => \N__12189\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__12189\,
            I => \N__12186\
        );

    \I__1226\ : Span4Mux_h
    port map (
            O => \N__12186\,
            I => \N__12183\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__12183\,
            I => \M_this_vga_signals_address_7\
        );

    \I__1224\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12177\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__12177\,
            I => \this_vga_signals.g1\
        );

    \I__1222\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12168\
        );

    \I__1221\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12168\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__12168\,
            I => \N__12165\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__12165\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__1218\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12159\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__12159\,
            I => \this_vga_signals.if_m2_1\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__12156\,
            I => \this_vga_signals.if_m2_1_cascade_\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__12153\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\
        );

    \I__1214\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12142\
        );

    \I__1213\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12137\
        );

    \I__1212\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12137\
        );

    \I__1211\ : InMux
    port map (
            O => \N__12147\,
            I => \N__12134\
        );

    \I__1210\ : InMux
    port map (
            O => \N__12146\,
            I => \N__12131\
        );

    \I__1209\ : InMux
    port map (
            O => \N__12145\,
            I => \N__12128\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__12142\,
            I => \N__12122\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__12137\,
            I => \N__12119\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__12134\,
            I => \N__12116\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__12131\,
            I => \N__12113\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__12128\,
            I => \N__12110\
        );

    \I__1203\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12107\
        );

    \I__1202\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12104\
        );

    \I__1201\ : InMux
    port map (
            O => \N__12125\,
            I => \N__12101\
        );

    \I__1200\ : Odrv12
    port map (
            O => \N__12122\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__12119\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__12116\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__12113\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__12110\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__12107\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__12104\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__12101\,
            I => \M_this_vga_ramdac_en_0\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__12084\,
            I => \N__12081\
        );

    \I__1191\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12078\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__12078\,
            I => \N__12075\
        );

    \I__1189\ : Span4Mux_h
    port map (
            O => \N__12075\,
            I => \N__12072\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__12072\,
            I => \N__12069\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__12069\,
            I => \M_this_vga_signals_address_2\
        );

    \I__1186\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__12063\,
            I => \this_vga_signals.g0_i_x4_0_4\
        );

    \I__1184\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12057\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__12057\,
            I => \N__12054\
        );

    \I__1182\ : Odrv12
    port map (
            O => \N__12054\,
            I => \this_vga_ramdac.m6\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__12051\,
            I => \G_463_cascade_\
        );

    \I__1180\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12045\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__12045\,
            I => \N__12042\
        );

    \I__1178\ : Span4Mux_v
    port map (
            O => \N__12042\,
            I => \N__12038\
        );

    \I__1177\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12035\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__12038\,
            I => \this_vga_ramdac.N_2807_reto\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__12035\,
            I => \this_vga_ramdac.N_2807_reto\
        );

    \I__1174\ : InMux
    port map (
            O => \N__12030\,
            I => \N__12024\
        );

    \I__1173\ : InMux
    port map (
            O => \N__12029\,
            I => \N__12024\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__12024\,
            I => \N_2_0\
        );

    \I__1171\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12018\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__12018\,
            I => \M_this_vga_signals_pixel_clk_0_0\
        );

    \I__1169\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12005\
        );

    \I__1168\ : InMux
    port map (
            O => \N__12014\,
            I => \N__12005\
        );

    \I__1167\ : InMux
    port map (
            O => \N__12013\,
            I => \N__11996\
        );

    \I__1166\ : InMux
    port map (
            O => \N__12012\,
            I => \N__11996\
        );

    \I__1165\ : InMux
    port map (
            O => \N__12011\,
            I => \N__11996\
        );

    \I__1164\ : InMux
    port map (
            O => \N__12010\,
            I => \N__11996\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__12005\,
            I => \G_463\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__11996\,
            I => \G_463\
        );

    \I__1161\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11988\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__11988\,
            I => \N__11985\
        );

    \I__1159\ : Odrv12
    port map (
            O => \N__11985\,
            I => \this_vga_ramdac.m19\
        );

    \I__1158\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11979\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__11979\,
            I => \N__11976\
        );

    \I__1156\ : Span4Mux_v
    port map (
            O => \N__11976\,
            I => \N__11972\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__11975\,
            I => \N__11969\
        );

    \I__1154\ : Span4Mux_h
    port map (
            O => \N__11972\,
            I => \N__11966\
        );

    \I__1153\ : InMux
    port map (
            O => \N__11969\,
            I => \N__11963\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__11966\,
            I => \this_vga_ramdac.N_2810_reto\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__11963\,
            I => \this_vga_ramdac.N_2810_reto\
        );

    \I__1150\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11955\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__11955\,
            I => \M_this_map_ram_write_data_0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11949\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__11949\,
            I => \N__11946\
        );

    \I__1146\ : Span4Mux_h
    port map (
            O => \N__11946\,
            I => \N__11943\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__11943\,
            I => \M_this_map_ram_write_data_5\
        );

    \I__1144\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11937\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__11937\,
            I => \M_this_map_ram_write_data_6\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_\
        );

    \I__1141\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11927\
        );

    \I__1140\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11924\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__11927\,
            I => \this_vga_signals.mult1_un61_sum_axb1_2\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__11924\,
            I => \this_vga_signals.mult1_un61_sum_axb1_2\
        );

    \I__1137\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11916\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__11916\,
            I => \N__11913\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__11913\,
            I => \this_vga_ramdac.N_24_mux\
        );

    \I__1134\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11906\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__11909\,
            I => \N__11903\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__11906\,
            I => \N__11900\
        );

    \I__1131\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11897\
        );

    \I__1130\ : Odrv12
    port map (
            O => \N__11900\,
            I => \this_vga_ramdac.N_2806_reto\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__11897\,
            I => \this_vga_ramdac.N_2806_reto\
        );

    \I__1128\ : InMux
    port map (
            O => \N__11892\,
            I => \N__11886\
        );

    \I__1127\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11883\
        );

    \I__1126\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11878\
        );

    \I__1125\ : InMux
    port map (
            O => \N__11889\,
            I => \N__11875\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__11886\,
            I => \N__11870\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11870\
        );

    \I__1122\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11867\
        );

    \I__1121\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11864\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__11878\,
            I => \N__11858\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__11875\,
            I => \N__11858\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__11870\,
            I => \N__11853\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__11867\,
            I => \N__11853\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__11864\,
            I => \N__11850\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__11863\,
            I => \N__11847\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__11858\,
            I => \N__11844\
        );

    \I__1113\ : Span4Mux_h
    port map (
            O => \N__11853\,
            I => \N__11839\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__11850\,
            I => \N__11839\
        );

    \I__1111\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11836\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__11844\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__11839\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__11836\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__11829\,
            I => \this_vga_signals.M_pcounter_q_3_0_cascade_\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__11826\,
            I => \N_2_0_cascade_\
        );

    \I__1105\ : InMux
    port map (
            O => \N__11823\,
            I => \N__11820\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__11820\,
            I => \N__11817\
        );

    \I__1103\ : Span12Mux_v
    port map (
            O => \N__11817\,
            I => \N__11814\
        );

    \I__1102\ : Odrv12
    port map (
            O => \N__11814\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__1101\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11808\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__11808\,
            I => \N__11804\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__11807\,
            I => \N__11801\
        );

    \I__1098\ : Span4Mux_v
    port map (
            O => \N__11804\,
            I => \N__11798\
        );

    \I__1097\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11795\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__11798\,
            I => \this_vga_ramdac.N_2811_reto\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__11795\,
            I => \this_vga_ramdac.N_2811_reto\
        );

    \I__1094\ : InMux
    port map (
            O => \N__11790\,
            I => \N__11787\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__11787\,
            I => \N__11784\
        );

    \I__1092\ : Span12Mux_v
    port map (
            O => \N__11784\,
            I => \N__11781\
        );

    \I__1091\ : Odrv12
    port map (
            O => \N__11781\,
            I => \this_vga_ramdac.m16\
        );

    \I__1090\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11774\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__11777\,
            I => \N__11771\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__11774\,
            I => \N__11768\
        );

    \I__1087\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11765\
        );

    \I__1086\ : Odrv12
    port map (
            O => \N__11768\,
            I => \this_vga_ramdac.N_2809_reto\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__11765\,
            I => \this_vga_ramdac.N_2809_reto\
        );

    \I__1084\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11757\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__11751\,
            I => \this_vga_ramdac.i2_mux\
        );

    \I__1080\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__11745\,
            I => \N__11741\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__11744\,
            I => \N__11738\
        );

    \I__1077\ : Span4Mux_h
    port map (
            O => \N__11741\,
            I => \N__11735\
        );

    \I__1076\ : InMux
    port map (
            O => \N__11738\,
            I => \N__11732\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__11735\,
            I => \this_vga_ramdac.N_2808_reto\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__11732\,
            I => \this_vga_ramdac.N_2808_reto\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__11727\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_\
        );

    \I__1072\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11721\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11718\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__11718\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__1069\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__11712\,
            I => \this_vga_signals.N_3_2_0_1\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__11709\,
            I => \this_vga_signals.mult1_un61_sum_axb1_3_cascade_\
        );

    \I__1066\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11703\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__11703\,
            I => \this_vga_signals.g1_1\
        );

    \I__1064\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11697\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__11697\,
            I => \this_vga_signals.g0_0\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__11694\,
            I => \this_vga_signals.g0_5_1_cascade_\
        );

    \I__1061\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11688\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__11688\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0_0_0_0\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__11685\,
            I => \N__11682\
        );

    \I__1058\ : InMux
    port map (
            O => \N__11682\,
            I => \N__11679\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__11679\,
            I => \N__11676\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__11676\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__11673\,
            I => \N__11670\
        );

    \I__1054\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11667\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__11667\,
            I => \this_vga_signals.g1_2_1\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__11664\,
            I => \this_vga_signals.if_i4_mux_cascade_\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__11661\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\
        );

    \I__1050\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11655\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__11655\,
            I => \this_vga_signals.g1_0_2\
        );

    \I__1048\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11649\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__11649\,
            I => \this_vga_signals.g0_1\
        );

    \I__1046\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11643\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__11643\,
            I => \this_vga_signals.g1_4_0\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__11640\,
            I => \N__11637\
        );

    \I__1043\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11634\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__11634\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__11631\,
            I => \this_vga_signals.g1_7_cascade_\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__11628\,
            I => \this_vga_signals.N_6_0_cascade_\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__11625\,
            I => \N__11620\
        );

    \I__1038\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11616\
        );

    \I__1037\ : InMux
    port map (
            O => \N__11623\,
            I => \N__11609\
        );

    \I__1036\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11609\
        );

    \I__1035\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11609\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__11616\,
            I => \N__11606\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__11609\,
            I => \N__11601\
        );

    \I__1032\ : Span4Mux_h
    port map (
            O => \N__11606\,
            I => \N__11598\
        );

    \I__1031\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11593\
        );

    \I__1030\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11593\
        );

    \I__1029\ : Span4Mux_h
    port map (
            O => \N__11601\,
            I => \N__11590\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__11598\,
            I => \M_this_vram_read_data_1\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__11593\,
            I => \M_this_vram_read_data_1\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__11590\,
            I => \M_this_vram_read_data_1\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__11583\,
            I => \N__11576\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__11582\,
            I => \N__11572\
        );

    \I__1023\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11569\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__11580\,
            I => \N__11566\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__11579\,
            I => \N__11563\
        );

    \I__1020\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11556\
        );

    \I__1019\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11556\
        );

    \I__1018\ : InMux
    port map (
            O => \N__11572\,
            I => \N__11556\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__11569\,
            I => \N__11553\
        );

    \I__1016\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11548\
        );

    \I__1015\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11548\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__11556\,
            I => \N__11545\
        );

    \I__1013\ : Span4Mux_h
    port map (
            O => \N__11553\,
            I => \N__11542\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__11548\,
            I => \M_this_vram_read_data_3\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__11545\,
            I => \M_this_vram_read_data_3\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__11542\,
            I => \M_this_vram_read_data_3\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__11535\,
            I => \this_vga_signals.g1_1_0_0_0_cascade_\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__11532\,
            I => \this_vga_signals.g1_0_1_0_0_cascade_\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__11529\,
            I => \N__11526\
        );

    \I__1006\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11523\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__11523\,
            I => \N__11520\
        );

    \I__1004\ : Span4Mux_v
    port map (
            O => \N__11520\,
            I => \N__11517\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__11517\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1002\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__11511\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1_0\
        );

    \I__1000\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11505\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__11505\,
            I => \N__11502\
        );

    \I__998\ : Odrv12
    port map (
            O => \N__11502\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \N__11496\
        );

    \I__996\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11493\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__11493\,
            I => \N__11490\
        );

    \I__994\ : Span4Mux_v
    port map (
            O => \N__11490\,
            I => \N__11487\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__11487\,
            I => \M_this_vga_signals_address_3\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__11484\,
            I => \this_vga_signals.mult1_un61_sum_axb1_cascade_\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__11481\,
            I => \this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_cascade_\
        );

    \I__990\ : InMux
    port map (
            O => \N__11478\,
            I => \N__11475\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__11475\,
            I => \N__11472\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__11472\,
            I => \this_vga_signals.if_i4_mux\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__11469\,
            I => \N__11466\
        );

    \I__986\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11463\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__11463\,
            I => \N__11460\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__11460\,
            I => \M_this_vga_signals_address_1\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__982\ : InMux
    port map (
            O => \N__11454\,
            I => \N__11451\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__11451\,
            I => \N__11448\
        );

    \I__980\ : Span4Mux_v
    port map (
            O => \N__11448\,
            I => \N__11445\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__11445\,
            I => \M_this_vga_signals_address_6\
        );

    \I__978\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11439\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__11439\,
            I => \this_vga_signals.mult1_un82_sum_c3\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__11436\,
            I => \N__11433\
        );

    \I__975\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11430\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__11430\,
            I => \this_vga_signals.N_219\
        );

    \I__973\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11418\
        );

    \I__972\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11418\
        );

    \I__971\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11418\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__11418\,
            I => \N__11415\
        );

    \I__969\ : Span4Mux_v
    port map (
            O => \N__11415\,
            I => \N__11410\
        );

    \I__968\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11405\
        );

    \I__967\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11405\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__11410\,
            I => \M_this_vram_read_data_2\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__11405\,
            I => \M_this_vram_read_data_2\
        );

    \I__964\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11392\
        );

    \I__963\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11385\
        );

    \I__962\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11385\
        );

    \I__961\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11385\
        );

    \I__960\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11380\
        );

    \I__959\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11380\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__11392\,
            I => \N__11375\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__11385\,
            I => \N__11375\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__11380\,
            I => \M_this_vram_read_data_0\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__11375\,
            I => \M_this_vram_read_data_0\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__953\ : CascadeBuf
    port map (
            O => \N__11367\,
            I => \N__11364\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__11364\,
            I => \N__11361\
        );

    \I__951\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11358\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__11358\,
            I => \N__11354\
        );

    \I__949\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11351\
        );

    \I__948\ : Span4Mux_v
    port map (
            O => \N__11354\,
            I => \N__11348\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__11351\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__11348\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__945\ : InMux
    port map (
            O => \N__11343\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__11340\,
            I => \N__11337\
        );

    \I__943\ : CascadeBuf
    port map (
            O => \N__11337\,
            I => \N__11334\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__11334\,
            I => \N__11331\
        );

    \I__941\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11328\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__11328\,
            I => \N__11324\
        );

    \I__939\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11321\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__11324\,
            I => \N__11318\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__11321\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__936\ : Odrv4
    port map (
            O => \N__11318\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__935\ : InMux
    port map (
            O => \N__11313\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__11310\,
            I => \N__11307\
        );

    \I__933\ : CascadeBuf
    port map (
            O => \N__11307\,
            I => \N__11304\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__11304\,
            I => \N__11301\
        );

    \I__931\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11298\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__11298\,
            I => \N__11294\
        );

    \I__929\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11291\
        );

    \I__928\ : Span4Mux_v
    port map (
            O => \N__11294\,
            I => \N__11288\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__11291\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__926\ : Odrv4
    port map (
            O => \N__11288\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__925\ : InMux
    port map (
            O => \N__11283\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__11280\,
            I => \N__11277\
        );

    \I__923\ : CascadeBuf
    port map (
            O => \N__11277\,
            I => \N__11274\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__11274\,
            I => \N__11271\
        );

    \I__921\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11268\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__11268\,
            I => \N__11264\
        );

    \I__919\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11261\
        );

    \I__918\ : Span4Mux_v
    port map (
            O => \N__11264\,
            I => \N__11258\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__11261\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__11258\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__915\ : InMux
    port map (
            O => \N__11253\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__11250\,
            I => \N__11247\
        );

    \I__913\ : CascadeBuf
    port map (
            O => \N__11247\,
            I => \N__11244\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__11244\,
            I => \N__11241\
        );

    \I__911\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11238\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__11238\,
            I => \N__11234\
        );

    \I__909\ : InMux
    port map (
            O => \N__11237\,
            I => \N__11231\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__11234\,
            I => \N__11228\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__11231\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__11228\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__905\ : InMux
    port map (
            O => \N__11223\,
            I => \bfn_7_25_0_\
        );

    \I__904\ : InMux
    port map (
            O => \N__11220\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__11217\,
            I => \N__11214\
        );

    \I__902\ : CascadeBuf
    port map (
            O => \N__11214\,
            I => \N__11211\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__11211\,
            I => \N__11208\
        );

    \I__900\ : InMux
    port map (
            O => \N__11208\,
            I => \N__11205\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__11205\,
            I => \N__11201\
        );

    \I__898\ : InMux
    port map (
            O => \N__11204\,
            I => \N__11198\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__11201\,
            I => \N__11195\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__11198\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__11195\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__11190\,
            I => \N__11187\
        );

    \I__893\ : InMux
    port map (
            O => \N__11187\,
            I => \N__11184\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__11184\,
            I => \M_this_vga_signals_address_5\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__11181\,
            I => \N__11178\
        );

    \I__890\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11175\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__11175\,
            I => \M_this_vga_signals_address_4\
        );

    \I__888\ : IoInMux
    port map (
            O => \N__11172\,
            I => \N__11169\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__11169\,
            I => \N__11166\
        );

    \I__886\ : Span4Mux_s2_h
    port map (
            O => \N__11166\,
            I => \N__11163\
        );

    \I__885\ : Sp12to4
    port map (
            O => \N__11163\,
            I => \N__11160\
        );

    \I__884\ : Span12Mux_v
    port map (
            O => \N__11160\,
            I => \N__11157\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__11157\,
            I => rgb_c_3
        );

    \I__882\ : IoInMux
    port map (
            O => \N__11154\,
            I => \N__11151\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__11151\,
            I => \N__11148\
        );

    \I__880\ : Odrv12
    port map (
            O => \N__11148\,
            I => this_vga_signals_vvisibility_i
        );

    \I__879\ : IoInMux
    port map (
            O => \N__11145\,
            I => \N__11142\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11139\
        );

    \I__877\ : IoSpan4Mux
    port map (
            O => \N__11139\,
            I => \N__11136\
        );

    \I__876\ : Span4Mux_s3_h
    port map (
            O => \N__11136\,
            I => \N__11133\
        );

    \I__875\ : Sp12to4
    port map (
            O => \N__11133\,
            I => \N__11130\
        );

    \I__874\ : Span12Mux_v
    port map (
            O => \N__11130\,
            I => \N__11127\
        );

    \I__873\ : Odrv12
    port map (
            O => \N__11127\,
            I => rgb_c_5
        );

    \I__872\ : IoInMux
    port map (
            O => \N__11124\,
            I => \N__11121\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__11121\,
            I => \N__11118\
        );

    \I__870\ : IoSpan4Mux
    port map (
            O => \N__11118\,
            I => \N__11115\
        );

    \I__869\ : Span4Mux_s3_h
    port map (
            O => \N__11115\,
            I => \N__11112\
        );

    \I__868\ : Odrv4
    port map (
            O => \N__11112\,
            I => rgb_c_1
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__11109\,
            I => \N__11106\
        );

    \I__866\ : CascadeBuf
    port map (
            O => \N__11106\,
            I => \N__11103\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__11103\,
            I => \N__11100\
        );

    \I__864\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11097\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__11097\,
            I => \N__11093\
        );

    \I__862\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11090\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__11093\,
            I => \N__11087\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__11090\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__859\ : Odrv4
    port map (
            O => \N__11087\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__11082\,
            I => \N__11079\
        );

    \I__857\ : CascadeBuf
    port map (
            O => \N__11079\,
            I => \N__11076\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__11076\,
            I => \N__11073\
        );

    \I__855\ : InMux
    port map (
            O => \N__11073\,
            I => \N__11070\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__11070\,
            I => \N__11066\
        );

    \I__853\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11063\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__11066\,
            I => \N__11060\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__11063\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__11060\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__849\ : InMux
    port map (
            O => \N__11055\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__11052\,
            I => \N__11049\
        );

    \I__847\ : CascadeBuf
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__11046\,
            I => \N__11043\
        );

    \I__845\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11040\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__11040\,
            I => \N__11036\
        );

    \I__843\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11033\
        );

    \I__842\ : Span4Mux_v
    port map (
            O => \N__11036\,
            I => \N__11030\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__11033\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__11030\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__839\ : InMux
    port map (
            O => \N__11025\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__11022\,
            I => \N__11019\
        );

    \I__837\ : CascadeBuf
    port map (
            O => \N__11019\,
            I => \N__11016\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__11016\,
            I => \N__11013\
        );

    \I__835\ : InMux
    port map (
            O => \N__11013\,
            I => \N__11010\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__11010\,
            I => \N__11006\
        );

    \I__833\ : InMux
    port map (
            O => \N__11009\,
            I => \N__11003\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__11006\,
            I => \N__11000\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__11003\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__11000\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__829\ : InMux
    port map (
            O => \N__10995\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__828\ : IoInMux
    port map (
            O => \N__10992\,
            I => \N__10989\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__10989\,
            I => \N__10986\
        );

    \I__826\ : Span4Mux_s0_h
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__825\ : Sp12to4
    port map (
            O => \N__10983\,
            I => \N__10980\
        );

    \I__824\ : Odrv12
    port map (
            O => \N__10980\,
            I => port_data_rw_0_i
        );

    \I__823\ : IoInMux
    port map (
            O => \N__10977\,
            I => \N__10974\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10971\
        );

    \I__821\ : Span4Mux_s3_h
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__820\ : Sp12to4
    port map (
            O => \N__10968\,
            I => \N__10965\
        );

    \I__819\ : Odrv12
    port map (
            O => \N__10965\,
            I => rgb_c_0
        );

    \I__818\ : IoInMux
    port map (
            O => \N__10962\,
            I => \N__10959\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__10959\,
            I => \N__10956\
        );

    \I__816\ : Span4Mux_s3_h
    port map (
            O => \N__10956\,
            I => \N__10953\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__10953\,
            I => rgb_c_2
        );

    \I__814\ : IoInMux
    port map (
            O => \N__10950\,
            I => \N__10947\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__10947\,
            I => \N__10944\
        );

    \I__812\ : Span4Mux_s3_h
    port map (
            O => \N__10944\,
            I => \N__10941\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__10941\,
            I => \N__10938\
        );

    \I__810\ : Sp12to4
    port map (
            O => \N__10938\,
            I => \N__10935\
        );

    \I__809\ : Odrv12
    port map (
            O => \N__10935\,
            I => rgb_c_4
        );

    \I__808\ : IoInMux
    port map (
            O => \N__10932\,
            I => \N__10929\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__10929\,
            I => \N__10926\
        );

    \I__806\ : Odrv12
    port map (
            O => \N__10926\,
            I => port_nmib_0_i
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_20_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_19_0_\
        );

    \IN_MUX_bfv_20_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_vaddress_q_cry_7\,
            carryinitout => \bfn_20_20_0_\
        );

    \IN_MUX_bfv_19_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_19_0_\
        );

    \IN_MUX_bfv_19_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_haddress_q_cry_7\,
            carryinitout => \bfn_19_20_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_24_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_16_0_\
        );

    \IN_MUX_bfv_24_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_19_0_\
        );

    \IN_MUX_bfv_19_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_17_0_\
        );

    \IN_MUX_bfv_19_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_vaddress_q_3_cry_7\,
            carryinitout => \bfn_19_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_haddress_q_2_cry_7\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_28_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_28_21_0_\
        );

    \IN_MUX_bfv_28_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_external_address_q_cry_7\,
            carryinitout => \bfn_28_22_0_\
        );

    \IN_MUX_bfv_21_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_13_0_\
        );

    \IN_MUX_bfv_21_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_sprites_address_q_cry_7\,
            carryinitout => \bfn_21_14_0_\
        );

    \IN_MUX_bfv_7_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_24_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_7_25_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17160\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_1098_g\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34657\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17316\,
            GLOBALBUFFEROUTPUT => \N_515_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_ppu.port_data_rw_0_i_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__21404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26567\,
            lcout => port_data_rw_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11910\,
            in2 => \_gnd_net_\,
            in3 => \N__11882\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11891\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11982\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI497S8_9_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21408\,
            in2 => \_gnd_net_\,
            in3 => \N__15326\,
            lcout => port_nmib_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11889\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIM8094_0_9_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15327\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11890\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11881\,
            in2 => \_gnd_net_\,
            in3 => \N__12048\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_0_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17574\,
            in1 => \N__11096\,
            in2 => \N__17433\,
            in3 => \N__17436\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_24_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_1_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17578\,
            in1 => \N__11069\,
            in2 => \_gnd_net_\,
            in3 => \N__11055\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_2_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17575\,
            in1 => \N__11039\,
            in2 => \_gnd_net_\,
            in3 => \N__11025\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_3_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17579\,
            in1 => \N__11009\,
            in2 => \_gnd_net_\,
            in3 => \N__10995\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_4_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17576\,
            in1 => \N__11357\,
            in2 => \_gnd_net_\,
            in3 => \N__11343\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_5_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17580\,
            in1 => \N__11327\,
            in2 => \_gnd_net_\,
            in3 => \N__11313\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_6_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17577\,
            in1 => \N__11297\,
            in2 => \_gnd_net_\,
            in3 => \N__11283\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_7_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17581\,
            in1 => \N__11267\,
            in2 => \_gnd_net_\,
            in3 => \N__11253\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \N__34632\,
            ce => 'H',
            sr => \N__28662\
        );

    \M_this_map_address_q_8_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__17582\,
            in1 => \N__11237\,
            in2 => \_gnd_net_\,
            in3 => \N__11223\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \N__34639\,
            ce => 'H',
            sr => \N__28659\
        );

    \M_this_map_address_q_9_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11204\,
            in1 => \N__17583\,
            in2 => \_gnd_net_\,
            in3 => \N__11220\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34639\,
            ce => 'H',
            sr => \N__28659\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3J5O7_9_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12148\,
            in2 => \_gnd_net_\,
            in3 => \N__12831\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI7VUTC_9_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__12149\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12677\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101001101"
        )
    port map (
            in0 => \N__11605\,
            in1 => \N__11414\,
            in2 => \N__11580\,
            in3 => \N__11396\,
            lcout => \this_vga_ramdac.m19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010110010111"
        )
    port map (
            in0 => \N__11604\,
            in1 => \N__11413\,
            in2 => \N__11579\,
            in3 => \N__11395\,
            lcout => \this_vga_ramdac.m16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIEDCEO4_9_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__12146\,
            in1 => \N__11508\,
            in2 => \_gnd_net_\,
            in3 => \N__11442\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__11581\,
            in1 => \N__11624\,
            in2 => \_gnd_net_\,
            in3 => \N__11400\,
            lcout => \this_vga_ramdac.N_24_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIF2OJ6_6_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__12126\,
            in1 => \N__14469\,
            in2 => \N__11436\,
            in3 => \N__12474\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_ac0_3_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__11478\,
            in1 => \N__12315\,
            in2 => \N__12360\,
            in3 => \N__12423\,
            lcout => \this_vga_signals.mult1_un82_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000111111"
        )
    port map (
            in0 => \N__11399\,
            in1 => \N__11427\,
            in2 => \N__11583\,
            in3 => \N__11623\,
            lcout => \this_vga_ramdac.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__13668\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13581\,
            lcout => \this_vga_signals.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIKHT15_9_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__13667\,
            in1 => \N__13580\,
            in2 => \N__15325\,
            in3 => \N__13890\,
            lcout => \M_this_vga_ramdac_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101001011"
        )
    port map (
            in0 => \N__11397\,
            in1 => \N__11426\,
            in2 => \N__11582\,
            in3 => \N__11619\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110101"
        )
    port map (
            in0 => \N__11425\,
            in1 => \N__11398\,
            in2 => \N__11625\,
            in3 => \N__11575\,
            lcout => \this_vga_ramdac.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_18_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001011"
        )
    port map (
            in0 => \N__14961\,
            in1 => \N__12162\,
            in2 => \N__11685\,
            in3 => \N__12678\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNITO6PD6_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110000010"
        )
    port map (
            in0 => \N__14958\,
            in1 => \N__12396\,
            in2 => \N__11535\,
            in3 => \N__12246\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIAQLVLB_2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__12125\,
            in1 => \N__11514\,
            in2 => \N__11532\,
            in3 => \N__11658\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_16_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__12174\,
            in1 => \N__14965\,
            in2 => \N__12333\,
            in3 => \N__12353\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_2_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__12352\,
            in1 => \N__12328\,
            in2 => \N__14967\,
            in3 => \N__12173\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIG45VS_9_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__12145\,
            in1 => \N__12295\,
            in2 => \_gnd_net_\,
            in3 => \N__12240\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000110000011"
        )
    port map (
            in0 => \N__13052\,
            in1 => \N__12980\,
            in2 => \N__14296\,
            in3 => \N__14462\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1\,
            ltout => \this_vga_signals.mult1_un61_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011111000001"
        )
    port map (
            in0 => \N__13794\,
            in1 => \N__14123\,
            in2 => \N__11484\,
            in3 => \N__12652\,
            lcout => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0,
            ltout => \this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m4_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__14865\,
            in1 => \N__13797\,
            in2 => \N__11481\,
            in3 => \N__12293\,
            lcout => \this_vga_signals.if_i4_mux\,
            ltout => \this_vga_signals.if_i4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__12294\,
            in1 => \N__11706\,
            in2 => \N__11664\,
            in3 => \N__11652\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIQSM9K2_2_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11724\,
            in1 => \N__12594\,
            in2 => \N__11661\,
            in3 => \N__11646\,
            lcout => \this_vga_signals.g1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIAJMMB_2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13796\,
            in1 => \N__14957\,
            in2 => \_gnd_net_\,
            in3 => \N__12235\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI2BF2A_2_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12654\,
            in1 => \N__12435\,
            in2 => \_gnd_net_\,
            in3 => \N__12585\,
            lcout => \this_vga_signals.g1_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111100001"
        )
    port map (
            in0 => \N__13795\,
            in1 => \N__14124\,
            in2 => \N__11640\,
            in3 => \N__12653\,
            lcout => this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_7_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000101"
        )
    port map (
            in0 => \N__13786\,
            in1 => \_gnd_net_\,
            in2 => \N__14138\,
            in3 => \N__12646\,
            lcout => \this_vga_signals.g1_7\,
            ltout => \this_vga_signals.g1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_7_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14956\,
            in2 => \N__11631\,
            in3 => \N__11930\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_m2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000100"
        )
    port map (
            in0 => \N__11715\,
            in1 => \N__12372\,
            in2 => \N__11628\,
            in3 => \N__11691\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_4_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101011011010"
        )
    port map (
            in0 => \N__14465\,
            in1 => \N__12584\,
            in2 => \N__11673\,
            in3 => \N__14293\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_10_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001011111"
        )
    port map (
            in0 => \N__14294\,
            in1 => \_gnd_net_\,
            in2 => \N__11727\,
            in3 => \N__14133\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_20_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12647\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14128\,
            lcout => \this_vga_signals.N_3_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_2_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000110000011"
        )
    port map (
            in0 => \N__13049\,
            in1 => \N__12979\,
            in2 => \N__14298\,
            in3 => \N__14464\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axb1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000101101"
        )
    port map (
            in0 => \N__12648\,
            in1 => \N__14132\,
            in2 => \N__11709\,
            in3 => \N__13787\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_6_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111101111"
        )
    port map (
            in0 => \N__14088\,
            in1 => \N__14270\,
            in2 => \N__12453\,
            in3 => \N__12973\,
            lcout => \this_vga_signals.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_5_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001000100"
        )
    port map (
            in0 => \N__14089\,
            in1 => \N__13767\,
            in2 => \_gnd_net_\,
            in3 => \N__12649\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_5_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111000110"
        )
    port map (
            in0 => \N__11931\,
            in1 => \N__11700\,
            in2 => \N__11694\,
            in3 => \N__12504\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_0_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14090\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13768\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_1_9_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110111011"
        )
    port map (
            in0 => \N__13660\,
            in1 => \N__13564\,
            in2 => \_gnd_net_\,
            in3 => \N__13880\,
            lcout => \this_vga_signals.g1_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000110000011"
        )
    port map (
            in0 => \N__13045\,
            in1 => \N__12974\,
            in2 => \N__14289\,
            in3 => \N__14450\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__11919\,
            in1 => \N__34733\,
            in2 => \N__11909\,
            in3 => \N__12014\,
            lcout => \this_vga_ramdac.N_2806_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__12015\,
            in1 => \N__34734\,
            in2 => \N__11863\,
            in3 => \N__12150\,
            lcout => \this_vga_ramdac.M_this_vga_ramdac_en_reto_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_RNIEKLV2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13092\,
            in1 => \N__12569\,
            in2 => \_gnd_net_\,
            in3 => \N__17071\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNITGFO3_0_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13150\,
            in2 => \N__11829\,
            in3 => \N__17310\,
            lcout => \N_2_0\,
            ltout => \N_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_1_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11826\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34594\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__34726\,
            in1 => \N__11823\,
            in2 => \N__11807\,
            in3 => \N__12013\,
            lcout => \this_vga_ramdac.N_2811_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__12011\,
            in1 => \N__11790\,
            in2 => \N__11777\,
            in3 => \N__34724\,
            lcout => \this_vga_ramdac.N_2809_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__34723\,
            in1 => \N__11760\,
            in2 => \N__11744\,
            in3 => \N__12010\,
            lcout => \this_vga_ramdac.N_2808_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.G_463_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12021\,
            in1 => \N__13106\,
            in2 => \_gnd_net_\,
            in3 => \N__12029\,
            lcout => \G_463\,
            ltout => \G_463_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__12041\,
            in1 => \N__12060\,
            in2 => \N__12051\,
            in3 => \N__34722\,
            lcout => \this_vga_ramdac.N_2807_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13107\,
            in2 => \_gnd_net_\,
            in3 => \N__12030\,
            lcout => \M_this_vga_signals_pixel_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__12012\,
            in1 => \N__11991\,
            in2 => \N__11975\,
            in3 => \N__34725\,
            lcout => \this_vga_ramdac.N_2810_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_0_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34158\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17427\,
            lcout => \M_this_map_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_5_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33459\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17428\,
            lcout => \M_this_map_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_6_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35439\,
            in2 => \_gnd_net_\,
            in3 => \N__17397\,
            lcout => \M_this_map_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12795\,
            in1 => \N__12684\,
            in2 => \N__16092\,
            in3 => \N__12702\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_m2_0_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110101000001"
        )
    port map (
            in0 => \N__16170\,
            in1 => \N__12066\,
            in2 => \N__11934\,
            in3 => \N__12180\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI8AIVHV_9_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__12867\,
            in1 => \N__12127\,
            in2 => \N__12198\,
            in3 => \N__12744\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011101000"
        )
    port map (
            in0 => \N__16116\,
            in1 => \N__12696\,
            in2 => \N__16175\,
            in3 => \N__12801\,
            lcout => \this_vga_signals.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16776\,
            in2 => \_gnd_net_\,
            in3 => \N__16542\,
            lcout => \this_vga_signals.vaddress_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011000101010"
        )
    port map (
            in0 => \N__16861\,
            in1 => \N__17309\,
            in2 => \N__17022\,
            in3 => \N__17116\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m2_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \N__12239\,
            in1 => \N__13791\,
            in2 => \N__12297\,
            in3 => \N__12419\,
            lcout => \this_vga_signals.if_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m2_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__12418\,
            in1 => \N__12285\,
            in2 => \N__13800\,
            in3 => \N__12236\,
            lcout => \this_vga_signals.if_m2_1\,
            ltout => \this_vga_signals.if_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110010100011"
        )
    port map (
            in0 => \N__14966\,
            in1 => \N__12303\,
            in2 => \N__12156\,
            in3 => \N__12332\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI43G6H2_9_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12153\,
            in3 => \N__12147\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_4_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12690\,
            in1 => \N__12774\,
            in2 => \N__12729\,
            in3 => \N__13452\,
            lcout => \this_vga_signals.g0_i_x4_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \d_m1_2_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12351\,
            in1 => \N__12292\,
            in2 => \_gnd_net_\,
            in3 => \N__12238\,
            lcout => this_vga_signals_un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIV3EFO_2_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12237\,
            in1 => \N__13793\,
            in2 => \N__12296\,
            in3 => \N__14960\,
            lcout => \this_vga_signals.d_N_3_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIO08E8_3_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13792\,
            in1 => \N__14127\,
            in2 => \_gnd_net_\,
            in3 => \N__12669\,
            lcout => \this_vga_signals.M_hcounter_q_RNIO08E8Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__14125\,
            in1 => \N__12821\,
            in2 => \N__14297\,
            in3 => \N__12501\,
            lcout => this_vga_signals_un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_0_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14930\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13798\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_2_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12234\,
            in1 => \N__12847\,
            in2 => \N__12261\,
            in3 => \N__12503\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_2_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001011"
        )
    port map (
            in0 => \N__12387\,
            in1 => \N__12915\,
            in2 => \N__12258\,
            in3 => \N__12204\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_o2_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101110001"
        )
    port map (
            in0 => \N__15024\,
            in1 => \N__14511\,
            in2 => \N__12255\,
            in3 => \N__12252\,
            lcout => \this_vga_signals.mult1_un89_sum_c3_1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g1_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12502\,
            in1 => \N__13799\,
            in2 => \N__12849\,
            in3 => \N__12233\,
            lcout => \this_vga_signals.N_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__14126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12655\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIMID621_5_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12656\,
            in1 => \N__12381\,
            in2 => \N__12888\,
            in3 => \N__12402\,
            lcout => \this_vga_signals.g0_i_x4_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_4_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000010011"
        )
    port map (
            in0 => \N__14412\,
            in1 => \N__14220\,
            in2 => \N__13051\,
            in3 => \N__12975\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axb1_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_17_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111100001"
        )
    port map (
            in0 => \N__12651\,
            in1 => \N__13747\,
            in2 => \N__12390\,
            in3 => \N__14057\,
            lcout => \this_vga_signals.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_8_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101110001001"
        )
    port map (
            in0 => \N__14056\,
            in1 => \N__12441\,
            in2 => \N__13784\,
            in3 => \N__12650\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_1\,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_0_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13748\,
            in1 => \N__12897\,
            in2 => \N__12375\,
            in3 => \N__12500\,
            lcout => \this_vga_signals.g1_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_1_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__14055\,
            in1 => \N__12467\,
            in2 => \_gnd_net_\,
            in3 => \N__14216\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_3_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110010"
        )
    port map (
            in0 => \N__14217\,
            in1 => \N__13036\,
            in2 => \N__12366\,
            in3 => \N__14410\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__12921\,
            in1 => \N__12480\,
            in2 => \N__12363\,
            in3 => \N__14218\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_3_1_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14219\,
            in1 => \N__13037\,
            in2 => \N__12507\,
            in3 => \N__14411\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__13847\,
            in1 => \N__14401\,
            in2 => \N__13563\,
            in3 => \N__13630\,
            lcout => \this_vga_signals.N_6_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_2_9_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__13629\,
            in1 => \N__13532\,
            in2 => \_gnd_net_\,
            in3 => \N__13846\,
            lcout => \this_vga_signals.N_234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011100011111"
        )
    port map (
            in0 => \N__13844\,
            in1 => \N__14400\,
            in2 => \N__13562\,
            in3 => \N__13627\,
            lcout => \this_vga_signals.SUM_3\,
            ltout => \this_vga_signals.SUM_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_6_1_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101011111"
        )
    port map (
            in0 => \N__14402\,
            in1 => \_gnd_net_\,
            in2 => \N__12456\,
            in3 => \N__14058\,
            lcout => \this_vga_signals.g0_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_2_9_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100101100011"
        )
    port map (
            in0 => \N__13845\,
            in1 => \N__14399\,
            in2 => \N__13561\,
            in3 => \N__13628\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIAA7K1_4_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14059\,
            in2 => \N__12444\,
            in3 => \N__14237\,
            lcout => \this_vga_signals.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000110000011"
        )
    port map (
            in0 => \N__13041\,
            in1 => \N__12969\,
            in2 => \N__14266\,
            in3 => \N__14403\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIC8D41_2_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14404\,
            in1 => \N__14920\,
            in2 => \N__13785\,
            in3 => \N__14238\,
            lcout => \this_vga_signals.g1_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_3_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011111000001"
        )
    port map (
            in0 => \N__13752\,
            in1 => \N__14086\,
            in2 => \N__13224\,
            in3 => \N__12673\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101100110111"
        )
    port map (
            in0 => \N__13645\,
            in1 => \N__13542\,
            in2 => \N__14460\,
            in3 => \N__13867\,
            lcout => \this_vga_signals.SUM_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13087\,
            in1 => \N__12570\,
            in2 => \_gnd_net_\,
            in3 => \N__17107\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34588\,
            ce => \N__17305\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__17108\,
            in1 => \N__13088\,
            in2 => \N__13131\,
            in3 => \N__13151\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34588\,
            ce => \N__17305\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__13158\,
            in1 => \N__14322\,
            in2 => \N__13885\,
            in3 => \N__13659\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__13666\,
            in1 => \N__13579\,
            in2 => \_gnd_net_\,
            in3 => \N__13886\,
            lcout => this_vga_signals_hvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011001000100"
        )
    port map (
            in0 => \N__13248\,
            in1 => \N__12711\,
            in2 => \N__15999\,
            in3 => \N__12513\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI5NOID_3_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13364\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIC44JP1_2_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__16089\,
            in1 => \N__13488\,
            in2 => \N__12516\,
            in3 => \N__13449\,
            lcout => \this_vga_signals.g3_0\,
            ltout => \this_vga_signals.g3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIGG1CK4_2_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001011010"
        )
    port map (
            in0 => \N__13247\,
            in1 => \_gnd_net_\,
            in2 => \N__12756\,
            in3 => \N__12810\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI90GQ8D_1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100111110000"
        )
    port map (
            in0 => \N__14532\,
            in1 => \N__12753\,
            in2 => \N__12747\,
            in3 => \N__13194\,
            lcout => \this_vga_signals.g1_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000110111001"
        )
    port map (
            in0 => \N__13203\,
            in1 => \N__13188\,
            in2 => \N__12738\,
            in3 => \N__15114\,
            lcout => \this_vga_signals.mult1_un47_sum_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__14619\,
            in1 => \N__14579\,
            in2 => \N__13377\,
            in3 => \N__13926\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_ns_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13437\,
            in2 => \N__12714\,
            in3 => \N__12762\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_ns\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111011010"
        )
    port map (
            in0 => \N__13441\,
            in1 => \N__15982\,
            in2 => \N__12705\,
            in3 => \N__13266\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14580\,
            in1 => \N__16779\,
            in2 => \_gnd_net_\,
            in3 => \N__13178\,
            lcout => \this_vga_signals.g0_i_x4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_1_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__16541\,
            in1 => \_gnd_net_\,
            in2 => \N__13378\,
            in3 => \N__16084\,
            lcout => \this_vga_signals.g0_i_x4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_0_a2_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13375\,
            in1 => \N__15998\,
            in2 => \N__12789\,
            in3 => \N__13442\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_ac0_2_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000100001"
        )
    port map (
            in0 => \N__13359\,
            in1 => \N__15981\,
            in2 => \N__13451\,
            in3 => \N__12785\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_2\,
            ltout => \this_vga_signals.mult1_un68_sum_ac0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000111"
        )
    port map (
            in0 => \N__16085\,
            in1 => \N__13179\,
            in2 => \N__12804\,
            in3 => \N__12768\,
            lcout => \this_vga_signals.g1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13367\,
            in1 => \N__15990\,
            in2 => \N__16778\,
            in3 => \N__13436\,
            lcout => \this_vga_signals.g0_2_0_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110011001"
        )
    port map (
            in0 => \N__14618\,
            in1 => \N__14571\,
            in2 => \_gnd_net_\,
            in3 => \N__13921\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15989\,
            in2 => \N__12777\,
            in3 => \N__16762\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_2_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15987\,
            in1 => \N__14572\,
            in2 => \N__13450\,
            in3 => \N__13365\,
            lcout => \this_vga_signals.g0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_a3_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13366\,
            in1 => \N__15988\,
            in2 => \N__16777\,
            in3 => \N__13435\,
            lcout => \this_vga_signals.N_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_x1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__14617\,
            in1 => \N__14570\,
            in2 => \N__13376\,
            in3 => \N__13920\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__16620\,
            in1 => \N__16761\,
            in2 => \_gnd_net_\,
            in3 => \N__16515\,
            lcout => \this_vga_signals.vaddress_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_11_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110111011"
        )
    port map (
            in0 => \N__13065\,
            in1 => \N__14094\,
            in2 => \_gnd_net_\,
            in3 => \N__14262\,
            lcout => \this_vga_signals.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIF18M2_5_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010011011001"
        )
    port map (
            in0 => \N__13053\,
            in1 => \N__12981\,
            in2 => \N__14288\,
            in3 => \N__14459\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x4_2_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI42KN6_5_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12891\,
            in3 => \N__12848\,
            lcout => \this_vga_signals.g0_i_x4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_0_a2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13380\,
            in1 => \N__13902\,
            in2 => \_gnd_net_\,
            in3 => \N__13445\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010000001111"
        )
    port map (
            in0 => \N__16078\,
            in1 => \N__15992\,
            in2 => \N__12879\,
            in3 => \N__12876\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000101011"
        )
    port map (
            in0 => \N__16079\,
            in1 => \N__16174\,
            in2 => \N__12870\,
            in3 => \N__13302\,
            lcout => \this_vga_signals.mult1_un75_sum_c2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIL0C14_6_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111001110000"
        )
    port map (
            in0 => \N__14408\,
            in1 => \N__13032\,
            in2 => \N__12858\,
            in3 => \N__12968\,
            lcout => \this_vga_signals.N_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_a0_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14210\,
            in2 => \_gnd_net_\,
            in3 => \N__14406\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_a0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010100010"
        )
    port map (
            in0 => \N__12967\,
            in1 => \N__14215\,
            in2 => \N__13050\,
            in3 => \N__14409\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_13_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100001000"
        )
    port map (
            in0 => \N__14407\,
            in1 => \N__13031\,
            in2 => \N__14254\,
            in3 => \N__12966\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_tz_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__14054\,
            in1 => \N__14211\,
            in2 => \_gnd_net_\,
            in3 => \N__14405\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_0_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__13059\,
            in1 => \N__13030\,
            in2 => \N__12984\,
            in3 => \N__12965\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_19_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15009\,
            in2 => \_gnd_net_\,
            in3 => \N__14919\,
            lcout => \this_vga_signals.if_N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14505\,
            in2 => \N__15023\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17268\,
            in1 => \N__14929\,
            in2 => \_gnd_net_\,
            in3 => \N__12909\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__34566\,
            ce => 'H',
            sr => \N__14849\
        );

    \this_vga_signals.M_hcounter_q_3_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17306\,
            in1 => \N__13783\,
            in2 => \_gnd_net_\,
            in3 => \N__12906\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__34566\,
            ce => 'H',
            sr => \N__14849\
        );

    \this_vga_signals.M_hcounter_q_4_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17269\,
            in1 => \N__14087\,
            in2 => \_gnd_net_\,
            in3 => \N__12903\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__34566\,
            ce => 'H',
            sr => \N__14849\
        );

    \this_vga_signals.M_hcounter_q_5_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17307\,
            in1 => \N__14248\,
            in2 => \_gnd_net_\,
            in3 => \N__12900\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__34566\,
            ce => 'H',
            sr => \N__14849\
        );

    \this_vga_signals.M_hcounter_q_6_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17270\,
            in1 => \N__14438\,
            in2 => \_gnd_net_\,
            in3 => \N__13170\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__34566\,
            ce => 'H',
            sr => \N__14849\
        );

    \this_vga_signals.M_hcounter_q_7_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17308\,
            in1 => \N__13868\,
            in2 => \_gnd_net_\,
            in3 => \N__13167\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__34566\,
            ce => 'H',
            sr => \N__14849\
        );

    \this_vga_signals.M_hcounter_q_8_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17271\,
            in1 => \N__13560\,
            in2 => \_gnd_net_\,
            in3 => \N__13164\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__34566\,
            ce => 'H',
            sr => \N__14849\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13655\,
            in2 => \_gnd_net_\,
            in3 => \N__13161\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34574\,
            ce => \N__14520\,
            sr => \N__14853\
        );

    \this_vga_signals.M_hcounter_q_RNISKQ82_7_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__13570\,
            in1 => \N__13992\,
            in2 => \N__13884\,
            in3 => \N__14449\,
            lcout => \this_vga_signals.un4_hsynclt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110111011"
        )
    port map (
            in0 => \N__13643\,
            in1 => \N__13569\,
            in2 => \_gnd_net_\,
            in3 => \N__13869\,
            lcout => \this_vga_signals.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNIAOTU3_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__13086\,
            in1 => \N__13152\,
            in2 => \N__13130\,
            in3 => \N__17056\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_pcounter_q_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNIQLNN4_1_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13126\,
            in2 => \N__13110\,
            in3 => \N__17301\,
            lcout => \N_3_0\,
            ltout => \N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13095\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101100110111"
        )
    port map (
            in0 => \N__13644\,
            in1 => \N__13568\,
            in2 => \N__14463\,
            in3 => \N__13870\,
            lcout => OPEN,
            ltout => \this_vga_signals.SUM_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_g0_i_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011010010001"
        )
    port map (
            in0 => \N__14261\,
            in1 => \N__13233\,
            in2 => \N__13227\,
            in3 => \N__14448\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_4_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33574\,
            in2 => \_gnd_net_\,
            in3 => \N__17432\,
            lcout => \M_this_map_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__16346\,
            in1 => \N__15252\,
            in2 => \N__13965\,
            in3 => \N__14766\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_a2_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15980\,
            in1 => \N__13444\,
            in2 => \_gnd_net_\,
            in3 => \N__13374\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQJ81Q1_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000110"
        )
    port map (
            in0 => \N__16071\,
            in1 => \N__16155\,
            in2 => \N__13197\,
            in3 => \N__13487\,
            lcout => \this_vga_signals.g1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_0_6_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__16760\,
            in1 => \N__16628\,
            in2 => \_gnd_net_\,
            in3 => \N__16536\,
            lcout => \this_vga_signals.vaddress_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_0_m2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010100101"
        )
    port map (
            in0 => \N__16537\,
            in1 => \N__15106\,
            in2 => \N__15060\,
            in3 => \N__14744\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110101"
        )
    port map (
            in0 => \N__14622\,
            in1 => \N__16780\,
            in2 => \N__13182\,
            in3 => \N__14703\,
            lcout => \this_vga_signals.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_661_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111001111000"
        )
    port map (
            in0 => \N__14664\,
            in1 => \N__16759\,
            in2 => \N__14708\,
            in3 => \N__13470\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1_661\,
            ltout => \this_vga_signals.mult1_un68_sum_axb1_661_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_0_a2_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15979\,
            in2 => \N__13269\,
            in3 => \N__16781\,
            lcout => \this_vga_signals.g0_2_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000010100"
        )
    port map (
            in0 => \N__15159\,
            in1 => \N__15232\,
            in2 => \N__15375\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001110"
        )
    port map (
            in0 => \N__15048\,
            in1 => \N__14659\,
            in2 => \N__13260\,
            in3 => \N__15100\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010000001"
        )
    port map (
            in0 => \N__15983\,
            in1 => \N__15233\,
            in2 => \N__13257\,
            in3 => \N__14568\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010101001"
        )
    port map (
            in0 => \N__16769\,
            in1 => \N__14660\,
            in2 => \N__13254\,
            in3 => \N__13473\,
            lcout => \this_vga_signals.mult1_un61_sum_c3\,
            ltout => \this_vga_signals.mult1_un61_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_0_a2_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15984\,
            in1 => \N__16770\,
            in2 => \N__13251\,
            in3 => \N__13363\,
            lcout => \this_vga_signals.N_4_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010111100101"
        )
    port map (
            in0 => \N__15047\,
            in1 => \N__14658\,
            in2 => \N__14745\,
            in3 => \N__15099\,
            lcout => \this_vga_signals.mult1_un47_sum_c3\,
            ltout => \this_vga_signals.mult1_un47_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16517\,
            in1 => \N__16768\,
            in2 => \N__13236\,
            in3 => \N__14707\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d_0\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_3_d_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_a2_0_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001010101"
        )
    port map (
            in0 => \N__14569\,
            in1 => \_gnd_net_\,
            in2 => \N__13491\,
            in3 => \N__14610\,
            lcout => \this_vga_signals.g0_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIEQV87_2_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13472\,
            in1 => \N__15986\,
            in2 => \N__16090\,
            in3 => \N__16538\,
            lcout => \this_vga_signals.g2_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_d_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__15234\,
            in1 => \N__14663\,
            in2 => \N__14709\,
            in3 => \N__13471\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111101"
        )
    port map (
            in0 => \N__14662\,
            in1 => \N__15050\,
            in2 => \N__15110\,
            in3 => \N__14746\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__16771\,
            in1 => \N__15991\,
            in2 => \_gnd_net_\,
            in3 => \N__13901\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_2_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13284\,
            in1 => \N__13443\,
            in2 => \N__13383\,
            in3 => \N__13379\,
            lcout => \this_vga_signals.g0_i_x4_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_a3_0_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011000011"
        )
    port map (
            in0 => \N__15120\,
            in1 => \N__16539\,
            in2 => \N__13296\,
            in3 => \N__14747\,
            lcout => \this_vga_signals.g0_i_x4_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__16540\,
            in1 => \N__16278\,
            in2 => \N__16782\,
            in3 => \N__16425\,
            lcout => \this_vga_signals.vsync_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICSHP_7_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16083\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16347\,
            lcout => OPEN,
            ltout => \this_vga_signals.vsync_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI1FF84_6_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__13932\,
            in1 => \N__13278\,
            in2 => \N__13272\,
            in3 => \N__16629\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI7QQL1_1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__16775\,
            in1 => \N__16176\,
            in2 => \N__16091\,
            in3 => \N__15993\,
            lcout => \this_vga_signals.un2_vsynclt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_10_1_i_o3_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101001"
        )
    port map (
            in0 => \N__14621\,
            in1 => \N__14748\,
            in2 => \N__15069\,
            in3 => \N__13922\,
            lcout => \this_vga_signals.mult1_un54_sum_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__15016\,
            in1 => \N__14507\,
            in2 => \_gnd_net_\,
            in3 => \N__17300\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34560\,
            ce => 'H',
            sr => \N__14848\
        );

    \this_vga_signals.M_hcounter_q_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14506\,
            in2 => \_gnd_net_\,
            in3 => \N__17299\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34560\,
            ce => 'H',
            sr => \N__14848\
        );

    \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14209\,
            in1 => \N__14431\,
            in2 => \_gnd_net_\,
            in3 => \N__13843\,
            lcout => \this_vga_signals.M_hcounter_d7lto7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13724\,
            in2 => \_gnd_net_\,
            in3 => \N__14905\,
            lcout => \this_vga_signals.un2_hsynclto3_0\,
            ltout => \this_vga_signals.un2_hsynclto3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__15017\,
            in1 => \N__14500\,
            in2 => \N__13677\,
            in3 => \N__14053\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hcounter_d7lt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__13674\,
            in1 => \N__13631\,
            in2 => \N__13584\,
            in3 => \N__13559\,
            lcout => \this_vga_signals.M_hcounter_d7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14838\,
            in2 => \_gnd_net_\,
            in3 => \N__17288\,
            lcout => \this_vga_signals.N_852_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14501\,
            in1 => \N__14309\,
            in2 => \_gnd_net_\,
            in3 => \N__15018\,
            lcout => \this_vga_signals.un2_hsynclt6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIEVMV1_4_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14475\,
            in1 => \N__14137\,
            in2 => \N__14295\,
            in3 => \N__14461\,
            lcout => \this_vga_signals.un2_hsynclt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIADGD1_1_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__14310\,
            in1 => \N__14278\,
            in2 => \N__14139\,
            in3 => \N__15019\,
            lcout => \this_vga_signals.un4_hsynclto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_1_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33979\,
            in2 => \_gnd_net_\,
            in3 => \N__17406\,
            lcout => \M_this_map_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIT6RN_8_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111010011"
        )
    port map (
            in0 => \N__15142\,
            in1 => \N__16423\,
            in2 => \N__15273\,
            in3 => \N__13974\,
            lcout => \this_vga_signals.SUM_2_i_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_6_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14783\,
            in2 => \N__15371\,
            in3 => \N__14806\,
            lcout => \this_vga_signals.SUM_2_i_1_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIPKB1_7_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__14807\,
            in1 => \N__15364\,
            in2 => \_gnd_net_\,
            in3 => \N__14817\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_1_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNITUMI_8_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001111"
        )
    port map (
            in0 => \N__16424\,
            in1 => \N__15182\,
            in2 => \N__13968\,
            in3 => \N__15272\,
            lcout => \this_vga_signals.SUM_2_i_1_2_3\,
            ltout => \this_vga_signals.SUM_2_i_1_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__16319\,
            in1 => \N__15245\,
            in2 => \N__14769\,
            in3 => \N__14765\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_N_2L1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14782\,
            in2 => \N__15370\,
            in3 => \N__14805\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010011001"
        )
    port map (
            in0 => \N__16274\,
            in1 => \N__15141\,
            in2 => \N__14682\,
            in3 => \N__16412\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_ns_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14790\,
            in2 => \N__14754\,
            in3 => \N__14670\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un40_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100011000011"
        )
    port map (
            in0 => \N__15049\,
            in1 => \N__14661\,
            in2 => \N__14751\,
            in3 => \N__14732\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_x1_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100010011"
        )
    port map (
            in0 => \N__16411\,
            in1 => \N__16273\,
            in2 => \N__15146\,
            in3 => \N__14678\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15216\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.g2_0_a2_5_1_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__14631\,
            in1 => \N__14620\,
            in2 => \_gnd_net_\,
            in3 => \N__14578\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_0_a2_5Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIUR0A01_3_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100011100111"
        )
    port map (
            in0 => \N__15985\,
            in1 => \N__16746\,
            in2 => \N__14541\,
            in3 => \N__14538\,
            lcout => \this_vga_signals.g2_0_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101001101"
        )
    port map (
            in0 => \N__15105\,
            in1 => \N__16508\,
            in2 => \N__16619\,
            in3 => \N__16709\,
            lcout => \this_vga_signals.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010011111"
        )
    port map (
            in0 => \N__16708\,
            in1 => \N__16511\,
            in2 => \N__16614\,
            in3 => \N__15104\,
            lcout => \this_vga_signals.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNID73S_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100001111"
        )
    port map (
            in0 => \N__15223\,
            in1 => \_gnd_net_\,
            in2 => \N__15186\,
            in3 => \N__16510\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m2_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15008\,
            in2 => \_gnd_net_\,
            in3 => \N__14959\,
            lcout => \this_vga_signals.if_m2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17253\,
            in2 => \_gnd_net_\,
            in3 => \N__17067\,
            lcout => \this_vga_signals.N_1098_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15600\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__15504\,
            sr => \N__15472\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15549\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34515\,
            ce => \N__15504\,
            sr => \N__15472\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_N_2L1_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101111111"
        )
    port map (
            in0 => \N__14784\,
            in1 => \N__15366\,
            in2 => \N__14811\,
            in3 => \N__15263\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15566\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34521\,
            ce => \N__15513\,
            sr => \N__15474\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15525\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34521\,
            ce => \N__15513\,
            sr => \N__15474\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIQE4H_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__15177\,
            in1 => \N__15212\,
            in2 => \_gnd_net_\,
            in3 => \N__15365\,
            lcout => \this_vga_signals.vaddress_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15565\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34521\,
            ce => \N__15513\,
            sr => \N__15474\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15598\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34521\,
            ce => \N__15513\,
            sr => \N__15474\
        );

    \this_vga_signals.un5_vaddress_if_m8_0_a3_1_1_1_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110110110111"
        )
    port map (
            in0 => \N__16407\,
            in1 => \N__16266\,
            in2 => \N__15147\,
            in3 => \N__15178\,
            lcout => \this_vga_signals.if_m8_0_a3_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15599\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__15509\,
            sr => \N__15476\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15578\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__15509\,
            sr => \N__15476\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15547\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__15509\,
            sr => \N__15476\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15548\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__15509\,
            sr => \N__15476\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15567\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__15509\,
            sr => \N__15476\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15579\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34525\,
            ce => \N__15509\,
            sr => \N__15476\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16320\,
            in2 => \_gnd_net_\,
            in3 => \N__16269\,
            lcout => OPEN,
            ltout => \this_vga_signals.un6_vvisibilitylto8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__16506\,
            in1 => \N__16603\,
            in2 => \N__15336\,
            in3 => \N__16710\,
            lcout => OPEN,
            ltout => \this_vga_signals.un6_vvisibilitylt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNINQIT3_5_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000011"
        )
    port map (
            in0 => \N__16711\,
            in1 => \N__15282\,
            in2 => \N__15333\,
            in3 => \N__16507\,
            lcout => this_vga_signals_vvisibility_1,
            ltout => \this_vga_signals_vvisibility_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIM8094_9_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16409\,
            in2 => \N__15330\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.vvisibility\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16268\,
            in1 => \N__16408\,
            in2 => \N__16337\,
            in3 => \N__16602\,
            lcout => \this_vga_signals.vaddress_ac0_9_0_a0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI01PG1_0_1_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__20977\,
            in1 => \N__18442\,
            in2 => \_gnd_net_\,
            in3 => \N__35075\,
            lcout => \this_ppu.N_1195_0_1\,
            ltout => \this_ppu.N_1195_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_0_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__15645\,
            in1 => \N__20978\,
            in2 => \N__15276\,
            in3 => \N__21527\,
            lcout => \this_ppu.M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34537\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15644\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15804\,
            in2 => \N__20081\,
            in3 => \N__15405\,
            lcout => \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_0_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20030\,
            in2 => \N__15825\,
            in3 => \N__15402\,
            lcout => \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_1_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20034\,
            in2 => \N__15722\,
            in3 => \N__15399\,
            lcout => \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_2_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15860\,
            in2 => \N__20083\,
            in3 => \N__15396\,
            lcout => \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_3_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15879\,
            in2 => \N__20082\,
            in3 => \N__15393\,
            lcout => \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_4_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15842\,
            in2 => \N__20084\,
            in3 => \N__15390\,
            lcout => \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_count_q_1_cry_5_s1\,
            carryout => \this_ppu.un1_M_count_q_1_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNO_0_7_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000011110"
        )
    port map (
            in0 => \N__21012\,
            in1 => \N__21533\,
            in2 => \N__15693\,
            in3 => \N__15387\,
            lcout => \this_ppu.M_count_q_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34816\,
            in2 => \_gnd_net_\,
            in3 => \N__17475\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34553\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34829\,
            in2 => \_gnd_net_\,
            in3 => \N__15384\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15450\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15420\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__34837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15435\,
            lcout => \this_reset_cond.M_stage_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15426\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17282\,
            in2 => \_gnd_net_\,
            in3 => \N__15480\,
            lcout => \this_vga_signals.N_852_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17284\,
            in1 => \N__16115\,
            in2 => \N__17117\,
            in3 => \N__17115\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__34516\,
            ce => 'H',
            sr => \N__15473\
        );

    \this_vga_signals.M_vcounter_q_1_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17286\,
            in1 => \N__16151\,
            in2 => \_gnd_net_\,
            in3 => \N__15414\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__34516\,
            ce => 'H',
            sr => \N__15473\
        );

    \this_vga_signals.M_vcounter_q_2_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17285\,
            in1 => \N__16047\,
            in2 => \_gnd_net_\,
            in3 => \N__15411\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__34516\,
            ce => 'H',
            sr => \N__15473\
        );

    \this_vga_signals.M_vcounter_q_3_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__17287\,
            in1 => \N__15941\,
            in2 => \_gnd_net_\,
            in3 => \N__15408\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__34516\,
            ce => 'H',
            sr => \N__15473\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16715\,
            in2 => \_gnd_net_\,
            in3 => \N__15582\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16509\,
            in2 => \_gnd_net_\,
            in3 => \N__15570\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16610\,
            in2 => \_gnd_net_\,
            in3 => \N__15552\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16336\,
            in2 => \_gnd_net_\,
            in3 => \N__15534\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16272\,
            in2 => \_gnd_net_\,
            in3 => \N__15531\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16410\,
            in2 => \_gnd_net_\,
            in3 => \N__15528\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34522\,
            ce => \N__15505\,
            sr => \N__15475\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15524\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34522\,
            ce => \N__15505\,
            sr => \N__15475\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16487\,
            in1 => \N__16335\,
            in2 => \N__16615\,
            in3 => \N__16267\,
            lcout => \this_vga_signals.M_vcounter_d7lto8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI4GQN4_0_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21575\,
            in1 => \N__21661\,
            in2 => \_gnd_net_\,
            in3 => \N__21616\,
            lcout => \this_ppu.N_132_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI4L615_0_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__21628\,
            in1 => \N__21591\,
            in2 => \N__20995\,
            in3 => \N__21663\,
            lcout => \this_ppu.un16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI4HJ86_0_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__21627\,
            in1 => \N__21662\,
            in2 => \N__21602\,
            in3 => \N__15656\,
            lcout => \this_ppu.N_1195_0\,
            ltout => \this_ppu.N_1195_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_2_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010010000"
        )
    port map (
            in0 => \N__15824\,
            in1 => \N__15769\,
            in2 => \N__15666\,
            in3 => \N__15663\,
            lcout => \this_ppu.M_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_0_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001111110011"
        )
    port map (
            in0 => \N__21592\,
            in1 => \N__15657\,
            in2 => \N__21673\,
            in3 => \N__21629\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIL508_7_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15686\,
            in2 => \_gnd_net_\,
            in3 => \N__15643\,
            lcout => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_1_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__15803\,
            in1 => \N__15770\,
            in2 => \N__15627\,
            in3 => \N__15737\,
            lcout => \this_ppu.M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_5_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__15740\,
            in1 => \N__15618\,
            in2 => \N__15779\,
            in3 => \N__15878\,
            lcout => \this_ppu.M_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_4_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000100000000"
        )
    port map (
            in0 => \N__15612\,
            in1 => \N__15772\,
            in2 => \N__15864\,
            in3 => \N__15739\,
            lcout => \this_ppu.M_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_6_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000000010"
        )
    port map (
            in0 => \N__15741\,
            in1 => \N__15606\,
            in2 => \N__15780\,
            in3 => \N__15841\,
            lcout => \this_ppu.M_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIDE0G_2_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15877\,
            in1 => \N__15859\,
            in2 => \N__15843\,
            in3 => \N__15820\,
            lcout => OPEN,
            ltout => \this_ppu.M_count_d_1_sqmuxa_1_i_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_RNIKM001_1_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15715\,
            in1 => \N__15802\,
            in2 => \N__15789\,
            in3 => \N__15786\,
            lcout => \this_ppu.M_count_d_0_sqmuxa_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_count_q_3_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100100000000"
        )
    port map (
            in0 => \N__15723\,
            in1 => \N__15771\,
            in2 => \N__15750\,
            in3 => \N__15738\,
            lcout => \this_ppu.M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34538\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16821\,
            lcout => \this_pixel_clk_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34546\,
            ce => 'H',
            sr => \N__34994\
        );

    \this_ppu.M_count_q_7_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__18448\,
            in1 => \N__15699\,
            in2 => \N__21020\,
            in3 => \N__21534\,
            lcout => \this_ppu.M_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34546\,
            ce => 'H',
            sr => \N__34994\
        );

    \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_2_1_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17859\,
            in2 => \_gnd_net_\,
            in3 => \N__35088\,
            lcout => \this_vga_signals.N_85\,
            ltout => \this_vga_signals.N_85_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__15672\,
            in1 => \N__21476\,
            in2 => \N__15675\,
            in3 => \N__22981\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_i_1_5_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__17837\,
            in1 => \N__17765\,
            in2 => \_gnd_net_\,
            in3 => \N__17682\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_444_i_i_o2_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__20898\,
            in1 => \_gnd_net_\,
            in2 => \N__21765\,
            in3 => \N__23144\,
            lcout => \this_vga_signals.N_124_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_1_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__17761\,
            in1 => \N__16216\,
            in2 => \N__17838\,
            in3 => \N__17680\,
            lcout => \this_vga_signals_M_this_state_q_srsts_0_1_i_a2_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0_2_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__17836\,
            in1 => \N__16217\,
            in2 => \N__17766\,
            in3 => \N__17681\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_0_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__21492\,
            in1 => \N__16898\,
            in2 => \N__16221\,
            in3 => \N__27607\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34561\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010101010"
        )
    port map (
            in0 => \N__16218\,
            in1 => \N__16928\,
            in2 => \N__17610\,
            in3 => \N__17858\,
            lcout => \M_this_substate_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34568\,
            ce => 'H',
            sr => \N__34990\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_i_1_6_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__17832\,
            in1 => \N__17755\,
            in2 => \_gnd_net_\,
            in3 => \N__17671\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16203\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34575\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_3_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33730\,
            in2 => \_gnd_net_\,
            in3 => \N__17385\,
            lcout => \M_this_map_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_2_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33845\,
            in2 => \_gnd_net_\,
            in3 => \N__17384\,
            lcout => \M_this_map_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__16141\,
            in1 => \N__16105\,
            in2 => \N__16048\,
            in3 => \N__15909\,
            lcout => \this_vga_signals.M_vcounter_d7lt8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__16716\,
            in1 => \N__16791\,
            in2 => \N__16803\,
            in3 => \N__16418\,
            lcout => \this_vga_signals.M_vcounter_d8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__16790\,
            in1 => \N__16717\,
            in2 => \N__16627\,
            in3 => \N__16516\,
            lcout => \this_vga_signals.un4_lvisibility_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16868\,
            in1 => \N__17146\,
            in2 => \_gnd_net_\,
            in3 => \N__16419\,
            lcout => \this_vga_signals.line_clk_1\,
            ltout => \this_vga_signals.line_clk_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICHRV3_7_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__16355\,
            in1 => \N__16341\,
            in2 => \N__16362\,
            in3 => \N__16270\,
            lcout => \M_this_vga_signals_line_clk_0\,
            ltout => \M_this_vga_signals_line_clk_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIGL6V4_0_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__21576\,
            in1 => \N__21674\,
            in2 => \N__16359\,
            in3 => \N__35083\,
            lcout => \this_ppu.M_state_q_RNIGL6V4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__16356\,
            in1 => \N__16342\,
            in2 => \N__16287\,
            in3 => \N__16271\,
            lcout => \this_ppu.M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_1_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100001000"
        )
    port map (
            in0 => \N__17283\,
            in1 => \N__16839\,
            in2 => \N__17015\,
            in3 => \N__17147\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_1_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__29792\,
            in1 => \N__29951\,
            in2 => \_gnd_net_\,
            in3 => \N__20723\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34520\,
            ce => 'H',
            sr => \N__19139\
        );

    \this_ppu.M_haddress_q_0_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110111110010"
        )
    port map (
            in0 => \N__21078\,
            in1 => \N__21114\,
            in2 => \N__31503\,
            in3 => \N__29950\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34520\,
            ce => 'H',
            sr => \N__19139\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_1_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16869\,
            in2 => \_gnd_net_\,
            in3 => \N__17118\,
            lcout => \this_vga_signals.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_10_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000000010000"
        )
    port map (
            in0 => \N__16971\,
            in1 => \N__23222\,
            in2 => \N__21444\,
            in3 => \N__27549\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__16830\,
            in1 => \N__16820\,
            in2 => \_gnd_net_\,
            in3 => \N__35071\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.G_425_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__16829\,
            in1 => \N__16819\,
            in2 => \_gnd_net_\,
            in3 => \N__35070\,
            lcout => \G_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_1_i_a2_1_1_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__27550\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35079\,
            lcout => \this_vga_signals.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_i_o2_8_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23431\,
            in1 => \N__23148\,
            in2 => \_gnd_net_\,
            in3 => \N__21729\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_152_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_8_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__35080\,
            in1 => \N__27551\,
            in2 => \N__16806\,
            in3 => \N__22928\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__16899\,
            in1 => \N__21469\,
            in2 => \N__17448\,
            in3 => \N__24422\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_0_a2_2_0_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24421\,
            in2 => \_gnd_net_\,
            in3 => \N__28914\,
            lcout => \this_vga_signals.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_4_0_wclke_3_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__30318\,
            in1 => \N__30239\,
            in2 => \N__30162\,
            in3 => \N__30048\,
            lcout => \this_sprites_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__21470\,
            in1 => \N__16900\,
            in2 => \N__16878\,
            in3 => \N__25225\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_i_1_10_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010101"
        )
    port map (
            in0 => \N__20899\,
            in1 => \N__27537\,
            in2 => \N__22992\,
            in3 => \N__21728\,
            lcout => \this_vga_signals.M_this_state_q_srsts_i_i_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_wclke_3_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__30317\,
            in1 => \N__30238\,
            in2 => \N__30161\,
            in3 => \N__30047\,
            lcout => \this_sprites_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_3_sn_m2_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27584\,
            in2 => \_gnd_net_\,
            in3 => \N__22881\,
            lcout => \N_383_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__21483\,
            in1 => \N__16901\,
            in2 => \N__16932\,
            in3 => \N__22882\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__21484\,
            in1 => \N__23315\,
            in2 => \N__16917\,
            in3 => \N__16902\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_i_1_4_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17831\,
            in1 => \N__17757\,
            in2 => \_gnd_net_\,
            in3 => \N__17670\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_i_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_11_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__23203\,
            in1 => \N__20901\,
            in2 => \N__17457\,
            in3 => \N__21730\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_d_4_sqmuxa_0_a3_0_a2_0_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22991\,
            in2 => \_gnd_net_\,
            in3 => \N__27519\,
            lcout => \N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_1_11_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110010"
        )
    port map (
            in0 => \N__23202\,
            in1 => \N__27520\,
            in2 => \N__23433\,
            in3 => \N__35089\,
            lcout => \this_vga_signals.M_this_state_q_srsts_i_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0_3_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17822\,
            in1 => \N__17756\,
            in2 => \_gnd_net_\,
            in3 => \N__17658\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_en_0_a3_0_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23210\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27536\,
            lcout => \M_this_state_d_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_map_ram_write_data_7_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35226\,
            in2 => \_gnd_net_\,
            in3 => \N__17375\,
            lcout => \M_this_map_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35076\,
            lcout => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17133\,
            in1 => \N__17272\,
            in2 => \_gnd_net_\,
            in3 => \N__17093\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_7_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__20454\,
            in1 => \N__20528\,
            in2 => \N__20401\,
            in3 => \N__18909\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34517\,
            ce => 'H',
            sr => \N__19141\
        );

    \this_ppu.M_haddress_q_5_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20527\,
            in2 => \_gnd_net_\,
            in3 => \N__18907\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34523\,
            ce => 'H',
            sr => \N__19140\
        );

    \this_vga_signals.M_lcounter_q_RNIL33N6_1_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__17148\,
            in1 => \N__17132\,
            in2 => \_gnd_net_\,
            in3 => \N__17094\,
            lcout => \this_vga_signals.un1_M_hcounter_d7_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__19293\,
            in1 => \N__19461\,
            in2 => \_gnd_net_\,
            in3 => \N__19315\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34526\,
            ce => \N__19401\,
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__19456\,
            in1 => \N__19227\,
            in2 => \_gnd_net_\,
            in3 => \N__21301\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34539\,
            ce => \N__19394\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_o2_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__21721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23430\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_153_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_qlde_i_i_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__35084\,
            in1 => \N__35261\,
            in2 => \N__17463\,
            in3 => \N__17502\,
            lcout => \M_this_data_count_qlde_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_9_8_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19316\,
            in1 => \N__19342\,
            in2 => \N__19271\,
            in3 => \N__19360\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__19361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19446\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34547\,
            ce => \N__19393\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_686_i_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__21722\,
            in1 => \N__23253\,
            in2 => \_gnd_net_\,
            in3 => \N__35085\,
            lcout => \N_686_i\,
            ltout => \N_686_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__19343\,
            in1 => \_gnd_net_\,
            in2 => \N__17460\,
            in3 => \N__19329\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34547\,
            ce => \N__19393\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__19454\,
            in1 => \N__20160\,
            in2 => \N__17550\,
            in3 => \N__35096\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34555\,
            ce => \N__19395\,
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_6_8_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19183\,
            in2 => \_gnd_net_\,
            in3 => \N__19211\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_8_8_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20113\,
            in1 => \N__20143\,
            in2 => \N__19514\,
            in3 => \N__20171\,
            lcout => OPEN,
            ltout => \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_8_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17517\,
            in1 => \N__21240\,
            in2 => \N__17511\,
            in3 => \N__17508\,
            lcout => \N_848\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__20114\,
            in1 => \N__19524\,
            in2 => \_gnd_net_\,
            in3 => \N__19452\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34555\,
            ce => \N__19395\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__19455\,
            in1 => \N__19200\,
            in2 => \N__26499\,
            in3 => \N__35097\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34555\,
            ce => \N__19395\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__19170\,
            in1 => \N__19453\,
            in2 => \_gnd_net_\,
            in3 => \N__19184\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34555\,
            ce => \N__19395\,
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_0_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__23760\,
            in1 => \N__29111\,
            in2 => \N__28946\,
            in3 => \N__19485\,
            lcout => \M_this_sprites_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34562\,
            ce => 'H',
            sr => \N__28660\
        );

    \this_vga_signals.N_444_i_i_a2_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17501\,
            in2 => \_gnd_net_\,
            in3 => \N__21720\,
            lcout => \this_vga_signals.N_154\,
            ltout => \this_vga_signals.N_154_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_3_0_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__17606\,
            in1 => \N__18377\,
            in2 => \N__17478\,
            in3 => \N__34695\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_5_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__35091\,
            in1 => \N__20367\,
            in2 => \_gnd_net_\,
            in3 => \N__20325\,
            lcout => \this_ppu.M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0_0_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__18384\,
            in1 => \N__27521\,
            in2 => \N__17879\,
            in3 => \N__35090\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_0_a2_0_0_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17906\,
            in1 => \N__23361\,
            in2 => \N__26540\,
            in3 => \N__18366\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001111"
        )
    port map (
            in0 => \N__18360\,
            in1 => \_gnd_net_\,
            in2 => \N__18354\,
            in3 => \N__18351\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_0_6_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__18345\,
            in1 => \N__32010\,
            in2 => \N__31667\,
            in3 => \N__31452\,
            lcout => \M_this_ppu_sprites_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_1_6_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__31453\,
            in1 => \N__18117\,
            in2 => \N__31986\,
            in3 => \N__31642\,
            lcout => \M_this_ppu_sprites_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_substate_d_0_sqmuxa_0_a3_0_a2_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17907\,
            in1 => \N__17872\,
            in2 => \N__26541\,
            in3 => \N__23360\,
            lcout => \N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_0_m2_0_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__17815\,
            in1 => \N__17737\,
            in2 => \_gnd_net_\,
            in3 => \N__17645\,
            lcout => \N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI01PG1_1_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__21011\,
            in1 => \N__18456\,
            in2 => \_gnd_net_\,
            in3 => \N__35086\,
            lcout => \this_ppu.N_1156_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIE07J4_0_1_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => port_dmab_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_2_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__18420\,
            in1 => \N__18995\,
            in2 => \N__19046\,
            in3 => \N__18410\,
            lcout => \M_this_ppu_oam_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIGJUB2_3_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__20361\,
            in1 => \N__18937\,
            in2 => \_gnd_net_\,
            in3 => \N__20319\,
            lcout => \this_ppu.un1_M_oam_idx_q_1_c1\,
            ltout => \this_ppu.un1_M_oam_idx_q_1_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_RNIHI6C2_2_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19038\,
            in2 => \N__18462\,
            in3 => \N__18993\,
            lcout => \this_ppu.un1_M_oam_idx_q_1_c3\,
            ltout => \this_ppu.un1_M_oam_idx_q_1_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_3_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20838\,
            in2 => \N__18459\,
            in3 => \N__18405\,
            lcout => \M_this_ppu_oam_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_2_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__20362\,
            in1 => \N__21016\,
            in2 => \_gnd_net_\,
            in3 => \N__18455\,
            lcout => \this_ppu.N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_4_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__18406\,
            in1 => \N__18968\,
            in2 => \N__20846\,
            in3 => \N__18426\,
            lcout => \this_ppu.M_oam_idx_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_1_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__18994\,
            in1 => \N__18404\,
            in2 => \_gnd_net_\,
            in3 => \N__18419\,
            lcout => \M_this_ppu_oam_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34589\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_0_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000101000"
        )
    port map (
            in0 => \N__18411\,
            in1 => \N__20366\,
            in2 => \N__18941\,
            in3 => \N__20324\,
            lcout => \M_this_ppu_oam_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34595\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_idx_q_RNI3VF_4_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19045\,
            in1 => \N__18992\,
            in2 => \N__18969\,
            in3 => \N__18933\,
            lcout => \this_ppu.N_144_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_6_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20453\,
            in1 => \N__20529\,
            in2 => \_gnd_net_\,
            in3 => \N__18908\,
            lcout => \M_this_ppu_map_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34524\,
            ce => 'H',
            sr => \N__19155\
        );

    \this_ppu.M_haddress_q_RNIRHU1G_1_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__29826\,
            in1 => \N__29961\,
            in2 => \_gnd_net_\,
            in3 => \N__20715\,
            lcout => \this_ppu.un1_M_haddress_q_3_c2\,
            ltout => \this_ppu.un1_M_haddress_q_3_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI81A2G_4_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20597\,
            in1 => \N__20230\,
            in2 => \N__18912\,
            in3 => \N__29726\,
            lcout => \this_ppu.un1_M_haddress_q_3_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18891\,
            in1 => \N__18873\,
            in2 => \_gnd_net_\,
            in3 => \N__29630\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_6_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__34721\,
            in1 => \N__20781\,
            in2 => \N__21087\,
            in3 => \N__21110\,
            lcout => \this_ppu.M_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_2_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__29949\,
            in1 => \N__29804\,
            in2 => \N__29742\,
            in3 => \N__20722\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34533\,
            ce => 'H',
            sr => \N__19154\
        );

    \this_ppu.M_haddress_q_RNI88B5_0_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29896\,
            in2 => \_gnd_net_\,
            in3 => \N__29947\,
            lcout => OPEN,
            ltout => \this_ppu.un2_hscroll_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNIVK7O_0_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001011"
        )
    port map (
            in0 => \N__29948\,
            in1 => \N__31552\,
            in2 => \N__18861\,
            in3 => \N__31480\,
            lcout => \M_this_ppu_sprites_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_3_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20231\,
            in1 => \N__29727\,
            in2 => \_gnd_net_\,
            in3 => \N__19163\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34533\,
            ce => 'H',
            sr => \N__19154\
        );

    \this_ppu.M_haddress_q_4_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__19164\,
            in1 => \N__20598\,
            in2 => \N__29743\,
            in3 => \N__20232\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34533\,
            ce => 'H',
            sr => \N__19154\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29628\,
            in1 => \N__19116\,
            in2 => \_gnd_net_\,
            in3 => \N__19101\,
            lcout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_wclke_3_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__30243\,
            in1 => \N__30294\,
            in2 => \N__30157\,
            in3 => \N__30054\,
            lcout => \this_sprites_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__19248\,
            in1 => \N__19457\,
            in2 => \_gnd_net_\,
            in3 => \N__19270\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34548\,
            ce => \N__19397\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__19449\,
            in1 => \N__19236\,
            in2 => \_gnd_net_\,
            in3 => \N__21258\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34556\,
            ce => \N__19396\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__20184\,
            in1 => \N__19451\,
            in2 => \_gnd_net_\,
            in3 => \N__21280\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34556\,
            ce => \N__19396\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__20127\,
            in1 => \N__19447\,
            in2 => \_gnd_net_\,
            in3 => \N__20147\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34556\,
            ce => \N__19396\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19448\,
            in1 => \N__19494\,
            in2 => \N__22839\,
            in3 => \N__25245\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34556\,
            ce => \N__19396\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__19450\,
            in1 => \N__20196\,
            in2 => \_gnd_net_\,
            in3 => \N__21332\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34556\,
            ce => \N__19396\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_c_0_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19362\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_0_THRU_LUT4_0_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19841\,
            in2 => \N__19347\,
            in3 => \N__19323\,
            lcout => \M_this_data_count_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_1_THRU_LUT4_0_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19320\,
            in2 => \N__19911\,
            in3 => \N__19281\,
            lcout => \M_this_data_count_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_2_THRU_LUT4_0_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19845\,
            in2 => \N__19278\,
            in3 => \N__19239\,
            lcout => \M_this_data_count_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_3_THRU_LUT4_0_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21257\,
            in2 => \N__19912\,
            in3 => \N__19230\,
            lcout => \M_this_data_count_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_4_THRU_LUT4_0_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19849\,
            in2 => \N__21312\,
            in3 => \N__19215\,
            lcout => \M_this_data_count_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_6_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19212\,
            in2 => \N__19910\,
            in3 => \N__19194\,
            lcout => \M_this_data_count_q_s_6\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_6_THRU_LUT4_0_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19850\,
            in2 => \N__19191\,
            in3 => \N__20199\,
            lcout => \M_this_data_count_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_7_THRU_LUT4_0_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21333\,
            in2 => \N__19837\,
            in3 => \N__20187\,
            lcout => \M_this_data_count_q_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_8_THRU_LUT4_0_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19765\,
            in2 => \N__21285\,
            in3 => \N__20175\,
            lcout => \M_this_data_count_q_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_10_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20172\,
            in2 => \N__19835\,
            in3 => \N__20154\,
            lcout => \M_this_data_count_q_s_10\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_10_THRU_LUT4_0_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19758\,
            in2 => \N__20151\,
            in3 => \N__20118\,
            lcout => \M_this_data_count_q_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_11_THRU_LUT4_0_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20115\,
            in2 => \N__19836\,
            in3 => \N__19518\,
            lcout => \M_this_data_count_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_13_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19515\,
            in2 => \_gnd_net_\,
            in3 => \N__19497\,
            lcout => \M_this_data_count_q_s_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_0_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__23801\,
            in1 => \N__34173\,
            in2 => \N__27667\,
            in3 => \N__27554\,
            lcout => \N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNILG0GD_0_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__35081\,
            in1 => \N__21371\,
            in2 => \N__19479\,
            in3 => \N__21549\,
            lcout => \this_ppu.M_state_q_RNILG0GDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIPG425_1_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21550\,
            in1 => \N__30683\,
            in2 => \_gnd_net_\,
            in3 => \N__30821\,
            lcout => \this_ppu.un1_M_vaddress_q_2_c2\,
            ltout => \this_ppu.un1_M_vaddress_q_2_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21892\,
            in1 => \N__21933\,
            in2 => \N__20286\,
            in3 => \N__30631\,
            lcout => \this_ppu.un1_M_vaddress_q_2_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_5_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21843\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34582\,
            ce => 'H',
            sr => \N__21981\
        );

    \this_ppu.M_vaddress_q_7_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__21845\,
            in1 => \N__20281\,
            in2 => \N__21809\,
            in3 => \N__22124\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34582\,
            ce => 'H',
            sr => \N__21981\
        );

    \this_ppu.M_vaddress_q_6_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20283\,
            in1 => \N__21802\,
            in2 => \_gnd_net_\,
            in3 => \N__21844\,
            lcout => \M_this_ppu_map_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34582\,
            ce => 'H',
            sr => \N__21981\
        );

    \this_ppu.un1_M_haddress_q_2_cry_0_c_inv_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22080\,
            in2 => \N__29901\,
            in3 => \N__29965\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_0\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_1_c_inv_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22068\,
            in2 => \N__31794\,
            in3 => \N__29820\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_0\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_2_c_inv_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31835\,
            in2 => \N__22056\,
            in3 => \N__29734\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_1\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_3_c_inv_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22037\,
            in2 => \N__24924\,
            in3 => \N__20248\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_2\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_4_c_inv_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22022\,
            in2 => \N__20343\,
            in3 => \N__20614\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_3\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_5_c_inv_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22007\,
            in2 => \N__20298\,
            in3 => \N__20545\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_4\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_6_c_inv_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20467\,
            in1 => \N__22281\,
            in2 => \N__30897\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_5\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_7_c_inv_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20411\,
            in1 => \N__24885\,
            in2 => \N__22269\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_2_cry_6\,
            carryout => \this_ppu.un1_M_haddress_q_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_2_cry_7_c_RNIFEE22_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22101\,
            in1 => \N__22251\,
            in2 => \_gnd_net_\,
            in3 => \N__20370\,
            lcout => \this_ppu.vscroll8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_3_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20868\,
            in2 => \_gnd_net_\,
            in3 => \N__35094\,
            lcout => \this_ppu.M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc1_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31021\,
            in2 => \_gnd_net_\,
            in3 => \N__30944\,
            lcout => \this_ppu.un1_M_haddress_q_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_2_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__20331\,
            in1 => \N__20323\,
            in2 => \N__21024\,
            in3 => \N__35093\,
            lcout => \this_ppu.M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc2_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__30945\,
            in1 => \_gnd_net_\,
            in2 => \N__31026\,
            in3 => \N__31068\,
            lcout => \this_ppu.un1_M_haddress_q_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_4_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__20842\,
            in1 => \N__20811\,
            in2 => \N__20799\,
            in3 => \N__35095\,
            lcout => \this_ppu.M_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_6_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20837\,
            in1 => \N__20810\,
            in2 => \N__20798\,
            in3 => \N__35077\,
            lcout => \this_ppu.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_7_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__35078\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31671\,
            lcout => \this_ppu.M_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__20769\,
            in1 => \N__24033\,
            in2 => \N__23700\,
            in3 => \N__21228\,
            lcout => \M_this_ppu_vram_data_0\,
            ltout => \M_this_ppu_vram_data_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.vram_en_i_a2_0_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21125\,
            in1 => \N__22571\,
            in2 => \N__20742\,
            in3 => \N__22703\,
            lcout => \this_ppu.N_156\,
            ltout => \this_ppu.N_156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI22N1G_5_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31478\,
            in2 => \N__20739\,
            in3 => \N__21077\,
            lcout => \M_this_ppu_vram_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29629\,
            in1 => \N__20697\,
            in2 => \_gnd_net_\,
            in3 => \N__20679\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29633\,
            in1 => \N__20667\,
            in2 => \_gnd_net_\,
            in3 => \N__20652\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__22624\,
            in1 => \N__23691\,
            in2 => \N__21231\,
            in3 => \N__26850\,
            lcout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_13_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__31582\,
            in1 => \N__31479\,
            in2 => \N__21222\,
            in3 => \N__32211\,
            lcout => \this_sprites_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21198\,
            in1 => \N__21177\,
            in2 => \_gnd_net_\,
            in3 => \N__29632\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNO_0_1_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__31481\,
            in1 => \N__21079\,
            in2 => \_gnd_net_\,
            in3 => \N__21548\,
            lcout => \this_ppu.N_150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__23697\,
            in1 => \N__21159\,
            in2 => \N__22632\,
            in3 => \N__21153\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__23699\,
            in1 => \N__21147\,
            in2 => \N__21141\,
            in3 => \N__20907\,
            lcout => \M_this_ppu_vram_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_1_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__21109\,
            in1 => \N__21093\,
            in2 => \N__21086\,
            in3 => \N__34701\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20940\,
            in1 => \N__20925\,
            in2 => \_gnd_net_\,
            in3 => \N__29631\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIH92S_10_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24476\,
            in1 => \N__21756\,
            in2 => \N__23620\,
            in3 => \N__20900\,
            lcout => OPEN,
            ltout => \M_this_state_q_RNIH92SZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI373A1_8_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23221\,
            in2 => \N__21495\,
            in3 => \N__22938\,
            lcout => \M_this_state_q_RNI373A1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_13_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__21687\,
            in1 => \N__23429\,
            in2 => \N__21491\,
            in3 => \N__23618\,
            lcout => \M_this_state_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_12_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__21686\,
            in1 => \N__21426\,
            in2 => \N__23345\,
            in3 => \N__23619\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34563\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_7_i_a2_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22929\,
            in1 => \N__24433\,
            in2 => \_gnd_net_\,
            in3 => \N__25244\,
            lcout => \this_vga_signals.N_485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_a2_0_i_o2_7_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23428\,
            in2 => \_gnd_net_\,
            in3 => \N__35082\,
            lcout => \this_vga_signals.N_94_0\,
            ltout => \this_vga_signals.N_94_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_i_0_12_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__23617\,
            in1 => \N__21758\,
            in2 => \N__21429\,
            in3 => \N__27514\,
            lcout => \this_vga_signals.M_this_state_q_srsts_i_i_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un21_i_a3_1_1_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24432\,
            in1 => \N__23139\,
            in2 => \N__23344\,
            in3 => \N__27636\,
            lcout => OPEN,
            ltout => \this_vga_signals_un21_i_a3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIE07J4_1_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__21420\,
            in1 => \N__21774\,
            in2 => \N__21411\,
            in3 => \N__23106\,
            lcout => port_dmab_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_this_state_q_srsts_i_a2_7_8_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21328\,
            in1 => \N__21308\,
            in2 => \N__21281\,
            in3 => \N__21256\,
            lcout => \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_a3_0_0_7_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__23140\,
            in1 => \N__23432\,
            in2 => \_gnd_net_\,
            in3 => \N__24484\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_srsts_i_a3_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_0_7_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000101"
        )
    port map (
            in0 => \N__35092\,
            in1 => \N__27518\,
            in2 => \N__21780\,
            in3 => \N__25233\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_srsts_i_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__25234\,
            in1 => \N__24485\,
            in2 => \N__21777\,
            in3 => \N__21732\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI6Q0S_5_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22994\,
            in1 => \N__23138\,
            in2 => \N__23343\,
            in3 => \N__25232\,
            lcout => \M_this_state_q_RNI6Q0SZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_i_o2_12_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21757\,
            in2 => \_gnd_net_\,
            in3 => \N__21731\,
            lcout => \this_vga_signals.N_93_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_1_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100001111000"
        )
    port map (
            in0 => \N__30823\,
            in1 => \N__21551\,
            in2 => \N__30695\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_vaddress_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34576\,
            ce => 'H',
            sr => \N__21974\
        );

    \this_ppu.M_vaddress_q_0_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__21678\,
            in1 => \N__21636\,
            in2 => \N__21603\,
            in3 => \N__30822\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34576\,
            ce => 'H',
            sr => \N__21974\
        );

    \this_ppu.M_vaddress_q_2_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__30824\,
            in1 => \N__30633\,
            in2 => \N__30694\,
            in3 => \N__21552\,
            lcout => \this_ppu.M_vaddress_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34576\,
            ce => 'H',
            sr => \N__21974\
        );

    \this_ppu.M_vaddress_q_3_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21992\,
            in1 => \N__21934\,
            in2 => \_gnd_net_\,
            in3 => \N__30634\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34576\,
            ce => 'H',
            sr => \N__21974\
        );

    \this_ppu.M_vaddress_q_4_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__30632\,
            in1 => \N__21993\,
            in2 => \N__21941\,
            in3 => \N__21893\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34576\,
            ce => 'H',
            sr => \N__21974\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_0_c_inv_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23567\,
            in2 => \N__30780\,
            in3 => \N__30812\,
            lcout => \this_ppu.M_this_ppu_vram_addr_i_7\,
            ltout => OPEN,
            carryin => \bfn_19_17_0_\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_1_c_inv_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23552\,
            in2 => \N__31899\,
            in3 => \N__30676\,
            lcout => \this_ppu.M_vaddress_q_i_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_0\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_2_c_inv_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23537\,
            in2 => \N__30597\,
            in3 => \N__30624\,
            lcout => \this_ppu.M_vaddress_q_i_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_1\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_3_c_inv_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23519\,
            in2 => \N__24936\,
            in3 => \N__21932\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_2\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_4_c_inv_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23501\,
            in2 => \N__22245\,
            in3 => \N__21891\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_3\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_5_c_inv_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23483\,
            in2 => \N__33123\,
            in3 => \N__21842\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_7\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_4\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_6_c_inv_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23465\,
            in2 => \N__32910\,
            in3 => \N__21801\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_8\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_5\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_7_c_inv_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32094\,
            in2 => \N__23451\,
            in3 => \N__22123\,
            lcout => \this_ppu.M_this_ppu_map_addr_i_9\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_3_cry_6\,
            carryout => \this_ppu.un1_M_vaddress_q_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_LUT4_0_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22104\,
            lcout => \this_ppu.un1_M_vaddress_q_3_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_4_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__34830\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22092\,
            lcout => \this_reset_cond.M_stage_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_0_c_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22079\,
            in2 => \N__29897\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_19_19_0_\,
            carryout => \this_ppu.un1_M_haddress_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_1_c_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22067\,
            in2 => \N__31790\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_0\,
            carryout => \this_ppu.un1_M_haddress_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_2_c_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22049\,
            in2 => \N__31836\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_1\,
            carryout => \this_ppu.un1_M_haddress_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_3_c_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30943\,
            in2 => \N__22038\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_2\,
            carryout => \this_ppu.un1_M_haddress_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_4_c_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31025\,
            in2 => \N__22023\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_3\,
            carryout => \this_ppu.un1_M_haddress_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_5_c_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31067\,
            in2 => \N__22008\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_4\,
            carryout => \this_ppu.un1_M_haddress_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_6_c_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22280\,
            in2 => \N__30978\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_5\,
            carryout => \this_ppu.un1_M_haddress_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_haddress_q_cry_7_c_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22265\,
            in2 => \N__24912\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_haddress_q_cry_6\,
            carryout => \this_ppu.un1_M_haddress_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_7_c_RNI6VRP1_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__32157\,
            in1 => \N__31914\,
            in2 => \N__23733\,
            in3 => \N__22254\,
            lcout => \this_ppu.vscroll8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_4_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24853\,
            in1 => \N__26483\,
            in2 => \_gnd_net_\,
            in3 => \N__24833\,
            lcout => \M_this_oam_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34605\,
            ce => 'H',
            sr => \N__28657\
        );

    \this_ppu.un1_oam_data_axbxc1_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33041\,
            in2 => \_gnd_net_\,
            in3 => \N__32966\,
            lcout => \this_ppu.un1_M_vaddress_q_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29648\,
            in1 => \N__22227\,
            in2 => \_gnd_net_\,
            in3 => \N__22212\,
            lcout => \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22194\,
            in1 => \N__22176\,
            in2 => \_gnd_net_\,
            in3 => \N__29649\,
            lcout => \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_12_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__31501\,
            in1 => \N__31578\,
            in2 => \N__22164\,
            in3 => \N__32259\,
            lcout => \this_sprites_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34541\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__23695\,
            in1 => \N__24099\,
            in2 => \N__22628\,
            in3 => \N__22146\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__23696\,
            in1 => \N__22722\,
            in2 => \N__22716\,
            in3 => \N__29559\,
            lcout => \M_this_ppu_vram_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22692\,
            in1 => \N__22674\,
            in2 => \_gnd_net_\,
            in3 => \N__29627\,
            lcout => \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22659\,
            in1 => \_gnd_net_\,
            in2 => \N__29650\,
            in3 => \N__22647\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_mem_0_1_RNIL62PZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__23681\,
            in1 => \N__22620\,
            in2 => \N__22593\,
            in3 => \N__22287\,
            lcout => OPEN,
            ltout => \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__23698\,
            in1 => \N__22590\,
            in2 => \N__22584\,
            in3 => \N__24069\,
            lcout => \M_this_ppu_vram_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_2_6_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__22560\,
            in1 => \N__31492\,
            in2 => \N__31663\,
            in3 => \N__31941\,
            lcout => \M_this_ppu_sprites_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29623\,
            in1 => \N__22314\,
            in2 => \_gnd_net_\,
            in3 => \N__22299\,
            lcout => \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_10_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__24024\,
            in1 => \N__24153\,
            in2 => \N__22848\,
            in3 => \N__29007\,
            lcout => \M_this_sprites_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34557\,
            ce => 'H',
            sr => \N__28665\
        );

    \M_this_sprites_address_q_11_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__22854\,
            in1 => \N__24141\,
            in2 => \N__22863\,
            in3 => \N__29008\,
            lcout => \M_this_sprites_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34557\,
            ce => 'H',
            sr => \N__28665\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_11_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__27552\,
            in1 => \N__33608\,
            in2 => \N__29021\,
            in3 => \N__27681\,
            lcout => \N_792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_11_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__26298\,
            in1 => \N__30279\,
            in2 => \_gnd_net_\,
            in3 => \N__29091\,
            lcout => \M_this_sprites_address_qc_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_10_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27680\,
            in1 => \N__29003\,
            in2 => \N__33753\,
            in3 => \N__27553\,
            lcout => \N_795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_13_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__26310\,
            in1 => \N__29114\,
            in2 => \N__23157\,
            in3 => \N__30084\,
            lcout => \M_this_sprites_address_qc_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27504\,
            in2 => \_gnd_net_\,
            in3 => \N__35087\,
            lcout => \N_773_0\,
            ltout => \N_773_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_9_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22827\,
            in3 => \N__22930\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_443_i_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110011"
        )
    port map (
            in0 => \N__22824\,
            in1 => \N__28947\,
            in2 => \N__24489\,
            in3 => \N__27503\,
            lcout => \N_443_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_0_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__27297\,
            in1 => \N__34193\,
            in2 => \N__33609\,
            in3 => \N__27328\,
            lcout => \N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_13_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__28993\,
            in1 => \N__27668\,
            in2 => \N__35425\,
            in3 => \N__27505\,
            lcout => \N_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_en_0_i_0_0_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__27296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24483\,
            lcout => \N_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIUK1S_3_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23217\,
            in1 => \N__22993\,
            in2 => \N__24437\,
            in3 => \N__23608\,
            lcout => OPEN,
            ltout => \port_dmab_ac0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNI392H1_1_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24490\,
            in1 => \N__23137\,
            in2 => \N__23109\,
            in3 => \N__22893\,
            lcout => port_dmab_ac0_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_2_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__27329\,
            in1 => \N__35410\,
            in2 => \N__33908\,
            in3 => \N__27298\,
            lcout => \N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_2_13_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27418\,
            in1 => \N__25247\,
            in2 => \_gnd_net_\,
            in3 => \N__28941\,
            lcout => \N_809\,
            ltout => \N_809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_8_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001111"
        )
    port map (
            in0 => \N__24525\,
            in1 => \_gnd_net_\,
            in2 => \N__22998\,
            in3 => \N__26285\,
            lcout => \M_this_sprites_address_qc_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_394_0_i_i_o2_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__22995\,
            in1 => \N__25246\,
            in2 => \N__23346\,
            in3 => \N__27417\,
            lcout => \N_749_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2_0_a3_0_a2_0_a2_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22937\,
            in2 => \_gnd_net_\,
            in3 => \N__27416\,
            lcout => \this_vga_signals.M_this_sprites_address_d_0_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_4_13_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__27625\,
            in1 => \N__22892\,
            in2 => \_gnd_net_\,
            in3 => \N__27419\,
            lcout => \N_813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_address_delay.M_this_start_address_delay_out_i_0_i2_i_o2_0_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__23283\,
            in1 => \N__23245\,
            in2 => \_gnd_net_\,
            in3 => \N__23581\,
            lcout => \N_775_0\,
            ltout => \N_775_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_1_0_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23382\,
            in3 => \N__23379\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_en_1_sqmuxa_i_o2_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__23643\,
            in1 => \N__23246\,
            in2 => \N__23289\,
            in3 => \N__23582\,
            lcout => \N_122_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a2_i_o2_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__23285\,
            in1 => \N__23244\,
            in2 => \_gnd_net_\,
            in3 => \N__23580\,
            lcout => \N_87_0\,
            ltout => \N_87_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_data_count_d_5_sqmuxa_0_a3_0_a2_0_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23349\,
            in3 => \N__23342\,
            lcout => \N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__23284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23583\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_5_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34831\,
            in2 => \_gnd_net_\,
            in3 => \N__23229\,
            lcout => \this_reset_cond.M_stage_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_9_0_i_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__23223\,
            in1 => \N__24495\,
            in2 => \N__23638\,
            in3 => \N__27457\,
            lcout => \un1_M_this_state_q_9_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_0_c_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23568\,
            in2 => \N__30779\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_19_0_\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_1_c_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23553\,
            in2 => \N__31895\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_0\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_2_c_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23538\,
            in2 => \N__30590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_1\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_3_c_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32965\,
            in2 => \N__23523\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_2\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_4_c_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33042\,
            in2 => \N__23505\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_3\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_5_c_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33075\,
            in2 => \N__23487\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_4\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_6_c_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32997\,
            in2 => \N__23469\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_5\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_7_c_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23450\,
            in2 => \N__32124\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_vaddress_q_cry_6\,
            carryout => \this_ppu.un1_M_vaddress_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_vaddress_q_cry_7_THRU_LUT4_0_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23736\,
            lcout => \this_ppu.un1_M_vaddress_q_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_radreg_11_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__31672\,
            in1 => \N__31477\,
            in2 => \N__23724\,
            in3 => \N__32232\,
            lcout => \this_sprites_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIMU531_13_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32769\,
            in1 => \N__23639\,
            in2 => \N__32691\,
            in3 => \N__27527\,
            lcout => \un1_M_this_oam_address_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_1_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__32665\,
            in1 => \N__32774\,
            in2 => \N__32384\,
            in3 => \N__35074\,
            lcout => \N_1174_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_1_1_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__35072\,
            in1 => \N__32336\,
            in2 => \N__32844\,
            in3 => \N__32664\,
            lcout => \N_1190_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_0_1_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__32335\,
            in1 => \N__32773\,
            in2 => \N__32692\,
            in3 => \N__35073\,
            lcout => \N_1182_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNILNG41_3_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24772\,
            in1 => \N__26411\,
            in2 => \_gnd_net_\,
            in3 => \N__26437\,
            lcout => \un1_M_this_oam_address_q_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_23_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35222\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34623\,
            ce => \N__28325\,
            sr => \N__34995\
        );

    \M_this_data_tmp_q_esr_18_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34623\,
            ce => \N__28325\,
            sr => \N__34995\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29651\,
            in1 => \N__24126\,
            in2 => \_gnd_net_\,
            in3 => \N__24111\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24093\,
            in1 => \N__24081\,
            in2 => \_gnd_net_\,
            in3 => \N__29656\,
            lcout => \this_sprites_ram.mem_mem_1_1_RNINA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29657\,
            in1 => \_gnd_net_\,
            in2 => \N__24063\,
            in3 => \N__24048\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_10_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__24181\,
            in1 => \N__26308\,
            in2 => \_gnd_net_\,
            in3 => \N__29112\,
            lcout => \M_this_sprites_address_qc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_0_0_wclke_3_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30219\,
            in1 => \N__30280\,
            in2 => \N__30123\,
            in3 => \N__30053\,
            lcout => \this_sprites_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_0_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23824\,
            in2 => \N__23775\,
            in3 => \N__23774\,
            lcout => \M_this_sprites_address_q_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_21_13_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_sprites_address_q_cry_0_THRU_LUT4_0_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27740\,
            in2 => \_gnd_net_\,
            in3 => \N__23745\,
            lcout => \un1_M_this_sprites_address_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_0\,
            carryout => \un1_M_this_sprites_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_2_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25410\,
            in2 => \_gnd_net_\,
            in3 => \N__23742\,
            lcout => \M_this_sprites_address_q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_1\,
            carryout => \un1_M_this_sprites_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_3_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25828\,
            in2 => \_gnd_net_\,
            in3 => \N__23739\,
            lcout => \M_this_sprites_address_q_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_2\,
            carryout => \un1_M_this_sprites_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_4_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26654\,
            in2 => \_gnd_net_\,
            in3 => \N__24384\,
            lcout => \M_this_sprites_address_q_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_3\,
            carryout => \un1_M_this_sprites_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_5_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28764\,
            in2 => \_gnd_net_\,
            in3 => \N__24381\,
            lcout => \M_this_sprites_address_q_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_4\,
            carryout => \un1_M_this_sprites_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_6_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27928\,
            in2 => \_gnd_net_\,
            in3 => \N__24378\,
            lcout => \M_this_sprites_address_q_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_5\,
            carryout => \un1_M_this_sprites_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_7_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25018\,
            in2 => \_gnd_net_\,
            in3 => \N__24375\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_6\,
            carryout => \un1_M_this_sprites_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_8_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24524\,
            in2 => \_gnd_net_\,
            in3 => \N__24372\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_21_14_0_\,
            carryout => \un1_M_this_sprites_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_9_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26050\,
            in2 => \_gnd_net_\,
            in3 => \N__24369\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_8\,
            carryout => \un1_M_this_sprites_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_10_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24194\,
            in2 => \_gnd_net_\,
            in3 => \N__24144\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_9\,
            carryout => \un1_M_this_sprites_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_1_11_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30293\,
            in2 => \_gnd_net_\,
            in3 => \N__24132\,
            lcout => \M_this_sprites_address_q_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_10\,
            carryout => \un1_M_this_sprites_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_12_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30198\,
            in2 => \_gnd_net_\,
            in3 => \N__24129\,
            lcout => \M_this_sprites_address_q_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_sprites_address_q_cry_11\,
            carryout => \un1_M_this_sprites_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_13_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010001100"
        )
    port map (
            in0 => \N__30102\,
            in1 => \N__24753\,
            in2 => \N__29022\,
            in3 => \N__24747\,
            lcout => \M_this_sprites_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34577\,
            ce => 'H',
            sr => \N__28664\
        );

    \M_this_sprites_address_q_12_LC_21_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__29087\,
            in1 => \N__24744\,
            in2 => \N__29020\,
            in3 => \N__24501\,
            lcout => \M_this_sprites_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34583\,
            ce => 'H',
            sr => \N__28663\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_7_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27678\,
            in1 => \N__28994\,
            in2 => \N__34197\,
            in3 => \N__27544\,
            lcout => OPEN,
            ltout => \N_807_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_7_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__24942\,
            in1 => \N__28999\,
            in2 => \N__24738\,
            in3 => \N__24735\,
            lcout => \M_this_sprites_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34583\,
            ce => 'H',
            sr => \N__28663\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_8_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27679\,
            in1 => \N__34016\,
            in2 => \N__29019\,
            in3 => \N__27545\,
            lcout => OPEN,
            ltout => \N_803_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_8_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__28995\,
            in1 => \N__24726\,
            in2 => \N__24720\,
            in3 => \N__24717\,
            lcout => \M_this_sprites_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34583\,
            ce => 'H',
            sr => \N__28663\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_a2_1_9_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__27459\,
            in1 => \N__33904\,
            in2 => \N__27666\,
            in3 => \N__28942\,
            lcout => \N_799\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_3_0_12_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__27632\,
            in1 => \N__30197\,
            in2 => \N__33457\,
            in3 => \N__27460\,
            lcout => \N_602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_this_state_q_3_0_i_0_o2_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__24494\,
            in1 => \N__24438\,
            in2 => \_gnd_net_\,
            in3 => \N__27458\,
            lcout => \this_vga_signals.un1_M_this_state_q_3_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_RNO_0_7_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__25001\,
            in1 => \N__26286\,
            in2 => \_gnd_net_\,
            in3 => \N__29071\,
            lcout => \M_this_sprites_address_qc_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32967\,
            lcout => \M_this_oam_ram_read_data_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_0_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30942\,
            lcout => \M_this_oam_ram_read_data_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc4_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__30974\,
            in1 => \N__31063\,
            in2 => \N__24908\,
            in3 => \N__26505\,
            lcout => \this_ppu.un1_M_haddress_q_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_2_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34609\,
            ce => \N__26374\,
            sr => \N__34987\
        );

    \M_this_data_tmp_q_esr_1_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34609\,
            ce => \N__26374\,
            sr => \N__34987\
        );

    \M_this_oam_address_q_0_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__32383\,
            in1 => \N__26496\,
            in2 => \_gnd_net_\,
            in3 => \N__32842\,
            lcout => \M_this_oam_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34612\,
            ce => 'H',
            sr => \N__28658\
        );

    \M_this_oam_address_q_5_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__24860\,
            in1 => \N__24834\,
            in2 => \N__24809\,
            in3 => \N__26498\,
            lcout => \M_this_oam_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34612\,
            ce => 'H',
            sr => \N__28658\
        );

    \M_this_oam_address_q_3_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__26497\,
            in1 => \N__26407\,
            in2 => \N__24779\,
            in3 => \N__26441\,
            lcout => \M_this_oam_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34612\,
            ce => 'H',
            sr => \N__28658\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_2_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32376\,
            in1 => \N__32778\,
            in2 => \N__25290\,
            in3 => \N__32571\,
            lcout => \N_746_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_5_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33463\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34617\,
            ce => \N__26381\,
            sr => \N__34991\
        );

    \M_this_data_tmp_q_esr_0_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34123\,
            lcout => \M_this_data_tmp_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34617\,
            ce => \N__26381\,
            sr => \N__34991\
        );

    \M_this_data_tmp_q_esr_4_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34617\,
            ce => \N__26381\,
            sr => \N__34991\
        );

    \M_this_data_tmp_q_esr_7_LC_21_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35200\,
            lcout => \M_this_data_tmp_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34617\,
            ce => \N__26381\,
            sr => \N__34991\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a2_28_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32377\,
            in1 => \N__32689\,
            in2 => \N__33606\,
            in3 => \N__32845\,
            lcout => \M_this_oam_ram_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_21_LC_21_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34624\,
            ce => \N__28327\,
            sr => \N__34993\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_4_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__26647\,
            in1 => \N__27682\,
            in2 => \N__33607\,
            in3 => \N__27546\,
            lcout => \N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_3_bm_1_LC_22_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__25251\,
            in1 => \N__27547\,
            in2 => \N__27770\,
            in3 => \N__25182\,
            lcout => \this_vga_signals.M_this_sprites_address_q_3_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_2_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__29115\,
            in1 => \N__26316\,
            in2 => \N__25380\,
            in3 => \N__29010\,
            lcout => \M_this_sprites_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__28666\
        );

    \M_this_sprites_address_q_RNO_0_9_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__26051\,
            in1 => \N__26309\,
            in2 => \_gnd_net_\,
            in3 => \N__29113\,
            lcout => OPEN,
            ltout => \M_this_sprites_address_qc_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_9_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__29009\,
            in1 => \N__26259\,
            in2 => \N__26247\,
            in3 => \N__26244\,
            lcout => \M_this_sprites_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__28666\
        );

    \M_this_sprites_address_q_3_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__29116\,
            in1 => \N__26028\,
            in2 => \N__25794\,
            in3 => \N__29011\,
            lcout => \M_this_sprites_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__28666\
        );

    \this_vga_signals.M_this_sprites_address_q_3_0_i_m2_3_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__25874\,
            in1 => \N__27677\,
            in2 => \N__33749\,
            in3 => \N__27543\,
            lcout => \N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIS5A21_0_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__27186\,
            in1 => \N__31457\,
            in2 => \N__31653\,
            in3 => \N__30842\,
            lcout => \M_this_ppu_sprites_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_2_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__25411\,
            in1 => \N__27676\,
            in2 => \N__33909\,
            in3 => \N__27542\,
            lcout => \N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_1_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__33416\,
            in1 => \N__27327\,
            in2 => \N__34050\,
            in3 => \N__27305\,
            lcout => \M_this_sprites_ram_write_data_iv_i_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_15_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35168\,
            lcout => \M_this_data_tmp_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34610\,
            ce => \N__28217\,
            sr => \N__34984\
        );

    \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_5_0_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26616\,
            in1 => \N__26598\,
            in2 => \N__26586\,
            in3 => \N__26556\,
            lcout => \this_vga_signals.M_this_state_q_srsts_0_0_a2_1_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_8_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32375\,
            in1 => \N__32572\,
            in2 => \N__28227\,
            in3 => \N__32779\,
            lcout => \N_54_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_ac0_1_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31012\,
            in2 => \_gnd_net_\,
            in3 => \N__30930\,
            lcout => \this_ppu.un1_oam_data_1_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_1_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__26492\,
            in1 => \N__32426\,
            in2 => \N__32690\,
            in3 => \N__32843\,
            lcout => \M_this_oam_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34615\,
            ce => 'H',
            sr => \N__28661\
        );

    \M_this_oam_address_q_2_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26406\,
            in1 => \N__26491\,
            in2 => \_gnd_net_\,
            in3 => \N__26445\,
            lcout => \M_this_oam_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34615\,
            ce => 'H',
            sr => \N__28661\
        );

    \M_this_data_tmp_q_esr_6_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34618\,
            ce => \N__26382\,
            sr => \N__34988\
        );

    \M_this_data_tmp_q_esr_3_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34618\,
            ce => \N__26382\,
            sr => \N__34988\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_6_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32437\,
            in1 => \N__32853\,
            in2 => \N__26352\,
            in3 => \N__32587\,
            lcout => \N_742_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_26_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32435\,
            in1 => \N__32850\,
            in2 => \N__33896\,
            in3 => \N__32582\,
            lcout => \N_34_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_4_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32436\,
            in1 => \N__32851\,
            in2 => \N__26961\,
            in3 => \N__32586\,
            lcout => \N_744_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_7_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32852\,
            in1 => \N__26940\,
            in2 => \N__32657\,
            in3 => \N__32438\,
            lcout => \N_56_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_16_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34159\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34625\,
            ce => \N__28328\,
            sr => \N__34992\
        );

    \M_this_data_tmp_q_esr_22_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35437\,
            lcout => \M_this_data_tmp_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34625\,
            ce => \N__28328\,
            sr => \N__34992\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_16_LC_22_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32453\,
            in1 => \N__32652\,
            in2 => \N__26919\,
            in3 => \N__32880\,
            lcout => \N_738_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_22_LC_22_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32454\,
            in1 => \N__32653\,
            in2 => \N__26898\,
            in3 => \N__32881\,
            lcout => \N_40_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29652\,
            in1 => \N__26877\,
            in2 => \_gnd_net_\,
            in3 => \N__26862\,
            lcout => \this_sprites_ram.mem_mem_2_0_RNINE6PZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_4_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__29016\,
            in1 => \N__29125\,
            in2 => \N__26841\,
            in3 => \N__26832\,
            lcout => \M_this_sprites_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__28667\
        );

    \this_vga_signals.M_this_sprites_address_q_0_i_m2_0_6_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__27921\,
            in1 => \N__27684\,
            in2 => \N__35406\,
            in3 => \N__27548\,
            lcout => OPEN,
            ltout => \N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_6_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__29017\,
            in1 => \N__29126\,
            in2 => \N__28113\,
            in3 => \N__28110\,
            lcout => \M_this_sprites_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__28667\
        );

    \M_this_sprites_address_q_1_LC_23_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27345\,
            in1 => \N__29018\,
            in2 => \_gnd_net_\,
            in3 => \N__27897\,
            lcout => \M_this_sprites_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => 'H',
            sr => \N__28667\
        );

    \this_vga_signals.M_this_sprites_address_q_3_0_5_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__28701\,
            in1 => \N__27683\,
            in2 => \N__33468\,
            in3 => \N__27555\,
            lcout => \N_595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_address_q_3_am_1_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__27766\,
            in1 => \N__27669\,
            in2 => \N__34036\,
            in3 => \N__27538\,
            lcout => \this_vga_signals.M_this_sprites_address_q_3_amZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_sprites_ram_write_data_iv_i_i_3_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__33742\,
            in1 => \N__27336\,
            in2 => \N__35211\,
            in3 => \N__27309\,
            lcout => \M_this_sprites_ram_write_data_iv_i_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNINGCA_0_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30778\,
            in2 => \_gnd_net_\,
            in3 => \N__30841\,
            lcout => \this_ppu.un2_vscroll_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_19_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33732\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34611\,
            ce => \N__28326\,
            sr => \N__34983\
        );

    \this_ppu.M_haddress_q_RNI4S061_1_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__31500\,
            in1 => \N__29766\,
            in2 => \N__31683\,
            in3 => \N__29838\,
            lcout => \M_this_ppu_sprites_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_10_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33897\,
            lcout => \M_this_data_tmp_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34616\,
            ce => \N__28213\,
            sr => \N__34985\
        );

    \M_this_data_tmp_q_esr_12_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34616\,
            ce => \N__28213\,
            sr => \N__34985\
        );

    \M_this_data_tmp_q_esr_13_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33447\,
            lcout => \M_this_data_tmp_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34616\,
            ce => \N__28213\,
            sr => \N__34985\
        );

    \M_this_data_tmp_q_esr_14_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35426\,
            lcout => \M_this_data_tmp_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34616\,
            ce => \N__28213\,
            sr => \N__34985\
        );

    \M_this_data_tmp_q_esr_8_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34166\,
            lcout => \M_this_data_tmp_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34616\,
            ce => \N__28213\,
            sr => \N__34985\
        );

    \M_this_data_tmp_q_esr_9_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34037\,
            lcout => \M_this_data_tmp_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34619\,
            ce => \N__28218\,
            sr => \N__34986\
        );

    \M_this_data_tmp_q_esr_11_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33731\,
            lcout => \M_this_data_tmp_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34619\,
            ce => \N__28218\,
            sr => \N__34986\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_3_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32459\,
            in1 => \N__32574\,
            in2 => \N__28182\,
            in3 => \N__32893\,
            lcout => \N_745_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_14_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32458\,
            in1 => \N__32573\,
            in2 => \N__28161\,
            in3 => \N__32892\,
            lcout => \N_739_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_5_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32859\,
            in1 => \N__32441\,
            in2 => \N__28137\,
            in3 => \N__32679\,
            lcout => \N_743_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_27_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32439\,
            in1 => \N__32667\,
            in2 => \N__33701\,
            in3 => \N__32860\,
            lcout => \N_32_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_11_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32442\,
            in1 => \N__32668\,
            in2 => \N__28395\,
            in3 => \N__32861\,
            lcout => \M_this_oam_ram_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_0_LC_23_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32858\,
            in1 => \N__32440\,
            in2 => \N__28374\,
            in3 => \N__32678\,
            lcout => \N_748_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_17_LC_23_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32666\,
            in1 => \N__32443\,
            in2 => \N__28338\,
            in3 => \N__32862\,
            lcout => \N_44_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_17_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34628\,
            ce => \N__28329\,
            sr => \N__34989\
        );

    \M_this_data_tmp_q_esr_20_LC_23_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33585\,
            lcout => \M_this_data_tmp_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34628\,
            ce => \N__28329\,
            sr => \N__34989\
        );

    \this_vga_signals.M_this_oam_ram_write_data_23_LC_23_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32863\,
            in1 => \N__28269\,
            in2 => \N__32693\,
            in3 => \N__32456\,
            lcout => \M_this_oam_ram_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_20_LC_23_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32455\,
            in1 => \N__32669\,
            in2 => \N__28248\,
            in3 => \N__32864\,
            lcout => \N_42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a2_30_LC_23_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32865\,
            in1 => \N__35438\,
            in2 => \N__32694\,
            in3 => \N__32457\,
            lcout => \M_this_oam_ram_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29676\,
            in1 => \N__29670\,
            in2 => \_gnd_net_\,
            in3 => \N__29658\,
            lcout => \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_haddress_q_RNI70261_2_LC_24_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__31502\,
            in1 => \N__31803\,
            in2 => \N__31678\,
            in3 => \N__29741\,
            lcout => \M_this_ppu_sprites_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30241\,
            in1 => \N__30295\,
            in2 => \N__30158\,
            in3 => \N__30051\,
            lcout => \this_sprites_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__30319\,
            in1 => \N__30240\,
            in2 => \N__30144\,
            in3 => \N__30050\,
            lcout => \this_sprites_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIIL4G1_2_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__31464\,
            in1 => \N__30552\,
            in2 => \N__31652\,
            in3 => \N__30642\,
            lcout => \M_this_ppu_sprites_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_sprites_address_q_5_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__29127\,
            in1 => \N__29043\,
            in2 => \N__29031\,
            in3 => \N__29012\,
            lcout => \M_this_sprites_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34598\,
            ce => 'H',
            sr => \N__28668\
        );

    \this_sprites_ram.mem_mem_7_0_wclke_3_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30320\,
            in1 => \N__30220\,
            in2 => \N__30159\,
            in3 => \N__30049\,
            lcout => \this_sprites_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_vaddress_q_RNIFH3G1_1_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__31499\,
            in1 => \N__30651\,
            in2 => \N__31677\,
            in3 => \N__30699\,
            lcout => \M_this_ppu_sprites_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_0_c_inv_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30840\,
            in2 => \N__30708\,
            in3 => \N__30765\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_24_16_0_\,
            carryout => \this_ppu.un2_vscroll_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_0_c_RNI9R5O_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30690\,
            in2 => \N__31848\,
            in3 => \N__30645\,
            lcout => \this_ppu.un2_vscroll_cry_0_c_RNI9R5OZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un2_vscroll_cry_0\,
            carryout => \this_ppu.un2_vscroll_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_vscroll_cry_1_c_RNIBU6O_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__30635\,
            in1 => \N__30589\,
            in2 => \_gnd_net_\,
            in3 => \N__30555\,
            lcout => \this_ppu.un2_vscroll_cry_1_c_RNIBU6OZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI53UU_6_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__30543\,
            in1 => \N__31482\,
            in2 => \N__31673\,
            in3 => \N__32178\,
            lcout => \M_this_ppu_sprites_addr_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30324\,
            in1 => \N__30242\,
            in2 => \N__30160\,
            in3 => \N__30052\,
            lcout => \this_sprites_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_0_c_inv_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29973\,
            in2 => \N__29847\,
            in3 => \N__29895\,
            lcout => \this_ppu.M_this_oam_ram_read_data_iZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_24_19_0_\,
            carryout => \this_ppu.un2_hscroll_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_0_c_RNICE4J_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29837\,
            in2 => \N__31755\,
            in3 => \N__29760\,
            lcout => \this_ppu.un2_hscroll_cry_0_c_RNICE4JZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un2_hscroll_cry_0\,
            carryout => \this_ppu.un2_hscroll_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un2_hscroll_cry_1_c_RNIEH5J_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__29753\,
            in1 => \N__31825\,
            in2 => \_gnd_net_\,
            in3 => \N__31806\,
            lcout => \this_ppu.un2_hscroll_cry_1_c_RNIEH5JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_0_RNISG75_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31789\,
            lcout => \M_this_oam_ram_read_data_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_1_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32373\,
            in1 => \N__32687\,
            in2 => \N__31746\,
            in3 => \N__32854\,
            lcout => \N_747_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_10_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32374\,
            in1 => \N__32688\,
            in2 => \N__31722\,
            in3 => \N__32855\,
            lcout => \M_this_oam_ram_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI43UU_6_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__31959\,
            in1 => \N__31704\,
            in2 => \N__31682\,
            in3 => \N__31437\,
            lcout => \M_this_ppu_sprites_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_12_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32857\,
            in1 => \N__32432\,
            in2 => \N__31089\,
            in3 => \N__32677\,
            lcout => \N_740_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_axbxc3_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__31050\,
            in1 => \N__31002\,
            in2 => \N__30970\,
            in3 => \N__30918\,
            lcout => \this_ppu.un1_M_haddress_q_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_19_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32856\,
            in1 => \N__32431\,
            in2 => \N__30882\,
            in3 => \N__32676\,
            lcout => \M_this_oam_ram_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un9lto7_4_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32255\,
            in1 => \N__32225\,
            in2 => \N__32201\,
            in3 => \N__32174\,
            lcout => \this_ppu.un9lto7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_9_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32429\,
            in1 => \N__32656\,
            in2 => \N__32142\,
            in3 => \N__32849\,
            lcout => \N_741_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_ac0_1_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33030\,
            in2 => \_gnd_net_\,
            in3 => \N__32943\,
            lcout => OPEN,
            ltout => \this_ppu.un1_oam_data_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc4_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__33071\,
            in1 => \N__32111\,
            in2 => \N__32097\,
            in3 => \N__32996\,
            lcout => \this_ppu.un1_M_vaddress_q_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_13_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32847\,
            in1 => \N__32430\,
            in2 => \N__32079\,
            in3 => \N__32686\,
            lcout => \M_this_oam_ram_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_15_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32428\,
            in1 => \N__32655\,
            in2 => \N__32061\,
            in3 => \N__32848\,
            lcout => \M_this_oam_ram_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_sqmuxa_i_o2_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32427\,
            in1 => \N__32654\,
            in2 => \_gnd_net_\,
            in3 => \N__32846\,
            lcout => \N_123_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un9lto7_5_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32009\,
            in1 => \N__31973\,
            in2 => \N__31958\,
            in3 => \N__31925\,
            lcout => \this_ppu.un9lto7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_oam_ram_read_data_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_18_LC_24_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32433\,
            in1 => \N__32680\,
            in2 => \N__33147\,
            in3 => \N__32876\,
            lcout => \M_this_oam_ram_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc2_LC_24_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__33067\,
            in1 => \N__33034\,
            in2 => \_gnd_net_\,
            in3 => \N__32949\,
            lcout => \this_ppu.un1_M_vaddress_q_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_24_LC_24_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32434\,
            in1 => \N__32681\,
            in2 => \N__34191\,
            in3 => \N__32877\,
            lcout => \N_38_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_0_a2_31_LC_24_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32460\,
            in1 => \N__32682\,
            in2 => \N__35221\,
            in3 => \N__32878\,
            lcout => \M_this_oam_ram_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_29_LC_24_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32895\,
            in1 => \N__32685\,
            in2 => \N__33467\,
            in3 => \N__32463\,
            lcout => \N_736_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_i_25_LC_24_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32461\,
            in1 => \N__32683\,
            in2 => \N__34041\,
            in3 => \N__32879\,
            lcout => \N_737_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_axbxc3_LC_24_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__33066\,
            in1 => \N__33029\,
            in2 => \N__32995\,
            in3 => \N__32942\,
            lcout => \this_ppu.un1_M_vaddress_q_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_oam_ram_write_data_21_LC_24_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32894\,
            in1 => \N__32684\,
            in2 => \N__32475\,
            in3 => \N__32462\,
            lcout => \M_this_oam_ram_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_8_LC_26_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34850\,
            in2 => \_gnd_net_\,
            in3 => \N__33312\,
            lcout => \this_reset_cond.M_stage_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_6_LC_26_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__34848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33327\,
            lcout => \this_reset_cond.M_stage_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_7_LC_26_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__34849\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33318\,
            lcout => \this_reset_cond.M_stage_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_external_address_q_0_LC_28_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35302\,
            in1 => \N__33269\,
            in2 => \N__33306\,
            in3 => \N__33305\,
            lcout => \M_this_external_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_28_21_0_\,
            carryout => \un1_M_this_external_address_q_cry_0\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_1_LC_28_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35311\,
            in1 => \N__33245\,
            in2 => \_gnd_net_\,
            in3 => \N__33234\,
            lcout => \M_this_external_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_0\,
            carryout => \un1_M_this_external_address_q_cry_1\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_2_LC_28_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35303\,
            in1 => \N__33224\,
            in2 => \_gnd_net_\,
            in3 => \N__33213\,
            lcout => \M_this_external_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_1\,
            carryout => \un1_M_this_external_address_q_cry_2\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_3_LC_28_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35312\,
            in1 => \N__33200\,
            in2 => \_gnd_net_\,
            in3 => \N__33189\,
            lcout => \M_this_external_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_2\,
            carryout => \un1_M_this_external_address_q_cry_3\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_4_LC_28_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35304\,
            in1 => \N__33179\,
            in2 => \_gnd_net_\,
            in3 => \N__33168\,
            lcout => \M_this_external_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_3\,
            carryout => \un1_M_this_external_address_q_cry_4\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_5_LC_28_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35313\,
            in1 => \N__33161\,
            in2 => \_gnd_net_\,
            in3 => \N__33150\,
            lcout => \M_this_external_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_4\,
            carryout => \un1_M_this_external_address_q_cry_5\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_6_LC_28_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35305\,
            in1 => \N__34241\,
            in2 => \_gnd_net_\,
            in3 => \N__34230\,
            lcout => \M_this_external_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_5\,
            carryout => \un1_M_this_external_address_q_cry_6\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_7_LC_28_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35310\,
            in1 => \N__34211\,
            in2 => \_gnd_net_\,
            in3 => \N__34200\,
            lcout => \M_this_external_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_6\,
            carryout => \un1_M_this_external_address_q_cry_7\,
            clk => \N__34631\,
            ce => 'H',
            sr => \N__34981\
        );

    \M_this_external_address_q_8_LC_28_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__35298\,
            in2 => \N__34070\,
            in3 => \N__34053\,
            lcout => \M_this_external_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_28_22_0_\,
            carryout => \un1_M_this_external_address_q_cry_8\,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \M_this_external_address_q_9_LC_28_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__34046\,
            in1 => \N__35306\,
            in2 => \N__33929\,
            in3 => \N__33912\,
            lcout => \M_this_external_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_8\,
            carryout => \un1_M_this_external_address_q_cry_9\,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \M_this_external_address_q_10_LC_28_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__33879\,
            in1 => \N__35299\,
            in2 => \N__33773\,
            in3 => \N__33756\,
            lcout => \M_this_external_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_9\,
            carryout => \un1_M_this_external_address_q_cry_10\,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \M_this_external_address_q_11_LC_28_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__33697\,
            in1 => \N__35307\,
            in2 => \N__33629\,
            in3 => \N__33612\,
            lcout => \M_this_external_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_10\,
            carryout => \un1_M_this_external_address_q_cry_11\,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \M_this_external_address_q_12_LC_28_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__33584\,
            in1 => \N__35300\,
            in2 => \N__33488\,
            in3 => \N__33471\,
            lcout => \M_this_external_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_11\,
            carryout => \un1_M_this_external_address_q_cry_12\,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \M_this_external_address_q_13_LC_28_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__33405\,
            in1 => \N__35308\,
            in2 => \N__33344\,
            in3 => \N__35442\,
            lcout => \M_this_external_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_12\,
            carryout => \un1_M_this_external_address_q_cry_13\,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \M_this_external_address_q_14_LC_28_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__35383\,
            in1 => \N__35301\,
            in2 => \N__35333\,
            in3 => \N__35316\,
            lcout => \M_this_external_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_M_this_external_address_q_cry_13\,
            carryout => \un1_M_this_external_address_q_cry_14\,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \M_this_external_address_q_15_LC_28_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__35108\,
            in1 => \N__35309\,
            in2 => \N__35201\,
            in3 => \N__35127\,
            lcout => \M_this_external_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34637\,
            ce => 'H',
            sr => \N__34982\
        );

    \this_reset_cond.M_stage_q_9_LC_32_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__34854\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34746\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34638\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
