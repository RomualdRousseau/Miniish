-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Jun 20 2021 15:53:16

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    write_address : in std_logic_vector(14 downto 0);
    write_data : in std_logic_vector(5 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    write_en : in std_logic;
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__15245\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal write_data_c_5 : std_logic;
signal write_data_c_4 : std_logic;
signal write_data_c_3 : std_logic;
signal write_data_c_2 : std_logic;
signal write_data_c_1 : std_logic;
signal write_data_c_0 : std_logic;
signal write_address_c_9 : std_logic;
signal write_address_c_8 : std_logic;
signal write_address_c_7 : std_logic;
signal write_address_c_6 : std_logic;
signal write_address_c_5 : std_logic;
signal write_address_c_4 : std_logic;
signal write_address_c_3 : std_logic;
signal write_address_c_2 : std_logic;
signal write_address_c_10 : std_logic;
signal write_address_c_1 : std_logic;
signal write_address_c_0 : std_logic;
signal \VCCG0\ : std_logic;
signal \this_vga_signals_N_170_i\ : std_logic;
signal \this_vga_signals_N_171_i\ : std_logic;
signal rgb5_i : std_logic;
signal vsync_c : std_logic;
signal \this_vga_signals_N_94_i\ : std_logic;
signal \this_vram.mem_out_bus0_0\ : std_logic;
signal \this_vram.mem_out_bus1_0\ : std_logic;
signal \this_vram.mem_out_bus0_2\ : std_logic;
signal \this_vram.mem_out_bus1_2\ : std_logic;
signal \this_vram.mem_out_bus0_3\ : std_logic;
signal \this_vram.mem_out_bus1_3\ : std_logic;
signal \this_vram.mem_out_bus0_4\ : std_logic;
signal \this_vram.mem_out_bus1_4\ : std_logic;
signal \this_vram.mem_out_bus1_5\ : std_logic;
signal \this_vram.mem_out_bus0_5\ : std_logic;
signal \this_vram.mem_out_bus3_0\ : std_logic;
signal \this_vram.mem_out_bus2_0\ : std_logic;
signal \this_vram.mem_mem_0_0_RNILGFZ0Z11\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIPOJZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_N_2362\ : std_logic;
signal \this_vram.mem_N_2364_cascade_\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \this_vram.mem_out_bus3_3\ : std_logic;
signal \this_vram.mem_out_bus2_3\ : std_logic;
signal \this_vram.mem_mem_0_1_RNINGF11Z0Z_0\ : std_logic;
signal \this_vram.mem_mem_2_1_RNIROJ11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_out_bus4_3\ : std_logic;
signal \this_vram.mem_out_bus6_3\ : std_logic;
signal \this_vram.mem_mem_4_1_RNI14P11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_2336_cascade_\ : std_logic;
signal \this_vram.mem_N_2335\ : std_logic;
signal \this_vram.mem_out_bus3_2\ : std_logic;
signal \this_vram.mem_out_bus2_2\ : std_logic;
signal \this_vram.mem_mem_2_1_RNIROJZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_mem_0_1_RNINGFZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus3_5\ : std_logic;
signal \this_vram.mem_out_bus2_5\ : std_logic;
signal \this_vram.mem_mem_0_2_RNIPGF11Z0Z_0\ : std_logic;
signal \this_vram.mem_mem_2_2_RNITOJ11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_2371_cascade_\ : std_logic;
signal \this_vram.mem_out_bus2_4\ : std_logic;
signal \this_vram.mem_out_bus3_4\ : std_logic;
signal \this_vram.mem_mem_0_2_RNIPGFZ0Z11\ : std_logic;
signal \this_vram.mem_mem_2_2_RNITOJZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_N_2326_cascade_\ : std_logic;
signal \this_vram.mem_N_2373\ : std_logic;
signal \M_this_vram_read_data_5\ : std_logic;
signal \this_vram.mem_N_2328\ : std_logic;
signal \M_this_vram_read_data_4\ : std_logic;
signal \this_vram.mem_N_2337\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vram.mem_out_bus0_1\ : std_logic;
signal \this_vram.mem_out_bus1_1\ : std_logic;
signal \this_vram.mem_out_bus3_1\ : std_logic;
signal \this_vram.mem_out_bus2_1\ : std_logic;
signal \this_vram.mem_mem_0_0_RNILGF11Z0Z_0\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIPOJ11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_out_bus6_0\ : std_logic;
signal \this_vram.mem_out_bus4_0\ : std_logic;
signal \this_vram.mem_WE_27\ : std_logic;
signal \this_vram.mem_out_bus5_0\ : std_logic;
signal \this_vram.mem_out_bus7_0\ : std_logic;
signal \this_vram.mem_mem_5_0_RNI18RZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_mem_4_0_RNIV3PZ0Z11\ : std_logic;
signal \this_vram.mem_N_2363\ : std_logic;
signal \this_vram.mem_N_2344\ : std_logic;
signal \this_vram.mem_N_2346\ : std_logic;
signal \this_vram.mem_G_25_0_cascade_\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \this_vram.mem_WE_21\ : std_logic;
signal \this_vram.mem_N_2327\ : std_logic;
signal \this_vram.mem_N_2353\ : std_logic;
signal \this_vram.mem_N_2355_cascade_\ : std_logic;
signal \this_vram.mem_G_25_0\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \this_vram.mem_out_bus4_4\ : std_logic;
signal \this_vram.mem_out_bus6_4\ : std_logic;
signal \this_vram.mem_mem_4_2_RNI34PZ0Z11\ : std_logic;
signal \this_vram.mem_WE_18\ : std_logic;
signal \this_vram.mem_out_bus6_1\ : std_logic;
signal \this_vram.mem_out_bus4_1\ : std_logic;
signal \this_vram.mem_out_bus5_1\ : std_logic;
signal \this_vram.mem_out_bus7_1\ : std_logic;
signal \this_vram.mem_mem_4_0_RNIV3P11Z0Z_0\ : std_logic;
signal \this_vram.mem_mem_5_0_RNI18R11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_2354\ : std_logic;
signal \this_vram.mem_WE_24\ : std_logic;
signal \this_vram.mem_out_bus4_2\ : std_logic;
signal \this_vram.mem_out_bus6_2\ : std_logic;
signal \this_vram.mem_mem_4_1_RNI14PZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_N_2345\ : std_logic;
signal \this_vram.mem_WE_15\ : std_logic;
signal \this_vga_signals.m24_0_1_cascade_\ : std_logic;
signal \this_vga_signals.N_25_cascade_\ : std_logic;
signal \this_vga_signals.m24_0_1_0\ : std_logic;
signal \this_vga_signals.m27_0_o2_1\ : std_logic;
signal \this_vga_signals.m27_0_0_cascade_\ : std_logic;
signal \this_vga_signals.i9_mux_cascade_\ : std_logic;
signal \this_vga_signals.N_40\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \M_this_vga_signals_address_8\ : std_logic;
signal \this_vga_signals.address_1_cry_0\ : std_logic;
signal \M_this_vga_signals_address_9\ : std_logic;
signal \this_vga_signals.address_1_cry_1\ : std_logic;
signal \M_this_vga_signals_address_10\ : std_logic;
signal \this_vga_signals.address_1_cry_2\ : std_logic;
signal \this_vga_signals.address_1_cry_3\ : std_logic;
signal \this_vga_signals.address_1_cry_4\ : std_logic;
signal \this_vram.mem_radregZ0Z_13\ : std_logic;
signal \this_vga_signals.address_1_cry_5\ : std_logic;
signal \this_vga_signals.address_1_cry_6\ : std_logic;
signal \this_vram.mem_radregZ0Z_14\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vga_signals.address_1_0_cry_0\ : std_logic;
signal \this_vga_signals.address_1\ : std_logic;
signal \this_vga_signals.address_1_0_cry_1\ : std_logic;
signal \this_vga_signals.address_1_0_3\ : std_logic;
signal \this_vga_signals.address_1_0_cry_2\ : std_logic;
signal \this_vga_signals.address_1_0_4\ : std_logic;
signal \this_vga_signals.address_1_0_cry_3\ : std_logic;
signal \this_vga_signals.address_1_0_5\ : std_logic;
signal \this_vga_signals.address_1_0_cry_4\ : std_logic;
signal \this_vga_signals.address_1_0_6\ : std_logic;
signal \this_vga_signals.address_1_0_cry_5\ : std_logic;
signal \this_vga_signals.address_1_0_7\ : std_logic;
signal \this_vga_signals.address_1_0_cry_6\ : std_logic;
signal \this_vga_signals.address_1_0_8\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \this_vga_signals.address_1_0_8_THRU_CO\ : std_logic;
signal \this_vga_signals.m27_0_o2_0_3\ : std_logic;
signal \this_vga_signals.N_36\ : std_logic;
signal \this_vga_signals.m27_0_a2_1_5\ : std_logic;
signal \this_vga_signals.m27_0_a2_1_5_cascade_\ : std_logic;
signal \this_vga_signals.N_68_cascade_\ : std_logic;
signal \this_vga_signals.m27_0_a2_1_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_0_i_a2_0_0\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_vstate_qZ0Z_1\ : std_logic;
signal \this_vga_signals.m24_0_0\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_9\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_10\ : std_logic;
signal \this_vga_signals.M_hstate_q_ns_i_i_1_0\ : std_logic;
signal \this_vga_signals.N_76_cascade_\ : std_logic;
signal \this_vga_signals.N_29_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_0\ : std_logic;
signal \this_vga_signals.address_1_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_2\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_4\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_7\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_0_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_1_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_2_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_3_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_4_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_5_THRU_CO\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_6_THRU_CO\ : std_logic;
signal \this_vga_signals.N_68\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \N_112_g\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_10\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.N_37_cascade_\ : std_logic;
signal \this_vga_signals.M_hstate_q_ns_i_i_2_0\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_11\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.M_hstate_d_0_sqmuxa_0_a2_0_a2_0_cascade_\ : std_logic;
signal \this_vga_signals.N_169_4\ : std_logic;
signal \this_vga_signals.M_hstate_d_0_sqmuxa\ : std_logic;
signal \this_vga_signals.N_169\ : std_logic;
signal \this_vga_signals.N_42\ : std_logic;
signal \this_vga_signals.N_46\ : std_logic;
signal \this_vga_signals.N_83\ : std_logic;
signal \this_vga_signals.M_hstate_qZ0Z_1\ : std_logic;
signal \this_vga_signals.N_27\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal clk_c_g : std_logic;
signal \this_vram.mem_out_bus6_5\ : std_logic;
signal \this_vram.mem_out_bus4_5\ : std_logic;
signal \this_vram.mem_mem_4_2_RNI34P11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_2372\ : std_logic;
signal \this_vram.mem_WE_12\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \this_vram.mem_out_bus9_5\ : std_logic;
signal \this_vram.mem_out_bus8_5\ : std_logic;
signal \this_vram.mem_mem_8_2_RNI9H021Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus5_2\ : std_logic;
signal \this_vram.mem_out_bus7_2\ : std_logic;
signal \this_vram.mem_mem_5_1_RNI38RZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus5_3\ : std_logic;
signal \this_vram.mem_out_bus7_3\ : std_logic;
signal \this_vram.mem_mem_5_1_RNI38R11Z0Z_0\ : std_logic;
signal \this_vram.mem_WE_9\ : std_logic;
signal \this_vram.mem_out_bus7_4\ : std_logic;
signal \this_vram.mem_out_bus5_4\ : std_logic;
signal \this_vram.mem_mem_5_2_RNI58RZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus7_5\ : std_logic;
signal \this_vram.mem_radregZ0Z_12\ : std_logic;
signal \this_vram.mem_out_bus5_5\ : std_logic;
signal \this_vram.mem_mem_5_2_RNI58R11Z0Z_0\ : std_logic;
signal \this_vram.mem_WE_6\ : std_logic;
signal \this_vram.mem_out_bus9_0\ : std_logic;
signal \this_vram.mem_out_bus8_0\ : std_logic;
signal \this_vram.mem_mem_8_0_RNI5HZ0Z021\ : std_logic;
signal \this_vram.mem_out_bus8_1\ : std_logic;
signal \this_vram.mem_out_bus9_1\ : std_logic;
signal \this_vram.mem_mem_8_0_RNI5H021Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus8_2\ : std_logic;
signal \this_vram.mem_out_bus9_2\ : std_logic;
signal \this_vram.mem_mem_8_1_RNI7HZ0Z021\ : std_logic;
signal \this_vram.mem_N_27\ : std_logic;
signal \this_vram.mem_WE_0\ : std_logic;
signal write_address_c_13 : std_logic;
signal write_address_c_12 : std_logic;
signal \this_vram.mem_N_29\ : std_logic;
signal write_address_c_14 : std_logic;
signal write_address_c_11 : std_logic;
signal \this_vram.mem_N_29_cascade_\ : std_logic;
signal write_en_c : std_logic;
signal \this_vram.mem_WE_3\ : std_logic;
signal \this_vram.mem_out_bus9_3\ : std_logic;
signal \this_vram.mem_out_bus8_3\ : std_logic;
signal \this_vram.mem_mem_8_1_RNI7H021Z0Z_0\ : std_logic;
signal \this_vram.mem_radregZ0Z_11\ : std_logic;
signal \this_vram.mem_out_bus8_4\ : std_logic;
signal \this_vram.mem_out_bus9_4\ : std_logic;
signal \this_vram.mem_mem_8_2_RNI9HZ0Z021\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal write_address_wire : std_logic_vector(14 downto 0);
signal write_data_wire : std_logic_vector(5 downto 0);
signal write_en_wire : std_logic;
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_8_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_8_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_8_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_8_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_8_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_8_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_8_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_9_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_9_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_9_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_9_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_9_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_9_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_9_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    write_address_wire <= write_address;
    write_data_wire <= write_data;
    write_en_wire <= write_en;
    \this_vram.mem_out_bus0_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= \N__9071\&\N__9290\&\N__9500\&\N__9707\&\N__9968\&\N__10175\&\N__11210\&\N__11447\&\N__11678\&\N__12464\&\N__12725\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= \N__5789\&\N__7460\&\N__7253\&\N__7043\&\N__6833\&\N__6623\&\N__6410\&\N__6203\&\N__5993\&\N__5582\&\N__5378\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7758\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7610\&'0'&'0'&'0';
    \this_vram.mem_out_bus0_3\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_2\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_1_physical_RADDR_wire\ <= \N__9064\&\N__9283\&\N__9494\&\N__9701\&\N__9962\&\N__10169\&\N__11204\&\N__11441\&\N__11672\&\N__12458\&\N__12719\;
    \this_vram.mem_mem_0_1_physical_WADDR_wire\ <= \N__5783\&\N__7454\&\N__7247\&\N__7037\&\N__6827\&\N__6617\&\N__6404\&\N__6197\&\N__5987\&\N__5576\&\N__5372\;
    \this_vram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4954\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4832\&'0'&'0'&'0';
    \this_vram.mem_out_bus0_5\ <= \this_vram.mem_mem_0_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_4\ <= \this_vram.mem_mem_0_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_2_physical_RADDR_wire\ <= \N__9052\&\N__9271\&\N__9488\&\N__9695\&\N__9956\&\N__10163\&\N__11198\&\N__11435\&\N__11666\&\N__12451\&\N__12713\;
    \this_vram.mem_mem_0_2_physical_WADDR_wire\ <= \N__5777\&\N__7448\&\N__7240\&\N__7031\&\N__6821\&\N__6611\&\N__6398\&\N__6191\&\N__5977\&\N__5570\&\N__5362\;
    \this_vram.mem_mem_0_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5124\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5002\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_1\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_0\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_0_physical_RADDR_wire\ <= \N__9040\&\N__9259\&\N__9478\&\N__9685\&\N__9946\&\N__10153\&\N__11191\&\N__11428\&\N__11660\&\N__12439\&\N__12703\;
    \this_vram.mem_mem_1_0_physical_WADDR_wire\ <= \N__5767\&\N__7442\&\N__7228\&\N__7021\&\N__6815\&\N__6605\&\N__6391\&\N__6184\&\N__5965\&\N__5564\&\N__5350\;
    \this_vram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7765\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7580\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_3\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_2\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_1_physical_RADDR_wire\ <= \N__9028\&\N__9247\&\N__9466\&\N__9673\&\N__9934\&\N__10141\&\N__11179\&\N__11416\&\N__11650\&\N__12427\&\N__12691\;
    \this_vram.mem_mem_1_1_physical_WADDR_wire\ <= \N__5755\&\N__7432\&\N__7216\&\N__7009\&\N__6805\&\N__6595\&\N__6379\&\N__6172\&\N__5953\&\N__5557\&\N__5338\;
    \this_vram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4940\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4828\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_5\ <= \this_vram.mem_mem_1_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_4\ <= \this_vram.mem_mem_1_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_2_physical_RADDR_wire\ <= \N__9016\&\N__9235\&\N__9454\&\N__9661\&\N__9922\&\N__10129\&\N__11167\&\N__11404\&\N__11638\&\N__12415\&\N__12679\;
    \this_vram.mem_mem_1_2_physical_WADDR_wire\ <= \N__5743\&\N__7420\&\N__7204\&\N__6997\&\N__6793\&\N__6583\&\N__6367\&\N__6160\&\N__5941\&\N__5545\&\N__5326\;
    \this_vram.mem_mem_1_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5113\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5003\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_1\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_0\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_0_physical_RADDR_wire\ <= \N__9004\&\N__9223\&\N__9442\&\N__9649\&\N__9910\&\N__10117\&\N__11155\&\N__11392\&\N__11626\&\N__12403\&\N__12667\;
    \this_vram.mem_mem_2_0_physical_WADDR_wire\ <= \N__5731\&\N__7408\&\N__7192\&\N__6985\&\N__6781\&\N__6571\&\N__6355\&\N__6148\&\N__5929\&\N__5533\&\N__5314\;
    \this_vram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7738\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7590\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_3\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_2\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_1_physical_RADDR_wire\ <= \N__8992\&\N__9211\&\N__9430\&\N__9637\&\N__9898\&\N__10105\&\N__11143\&\N__11380\&\N__11614\&\N__12391\&\N__12655\;
    \this_vram.mem_mem_2_1_physical_WADDR_wire\ <= \N__5719\&\N__7396\&\N__7180\&\N__6973\&\N__6769\&\N__6559\&\N__6343\&\N__6136\&\N__5917\&\N__5521\&\N__5302\;
    \this_vram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4927\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4816\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_5\ <= \this_vram.mem_mem_2_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_4\ <= \this_vram.mem_mem_2_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_2_physical_RADDR_wire\ <= \N__8980\&\N__9199\&\N__9418\&\N__9625\&\N__9886\&\N__10093\&\N__11131\&\N__11368\&\N__11602\&\N__12379\&\N__12643\;
    \this_vram.mem_mem_2_2_physical_WADDR_wire\ <= \N__5707\&\N__7384\&\N__7168\&\N__6961\&\N__6757\&\N__6547\&\N__6331\&\N__6124\&\N__5905\&\N__5509\&\N__5290\;
    \this_vram.mem_mem_2_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5112\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5036\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_1\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_0\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_0_physical_RADDR_wire\ <= \N__8968\&\N__9187\&\N__9406\&\N__9613\&\N__9874\&\N__10081\&\N__11119\&\N__11356\&\N__11590\&\N__12367\&\N__12631\;
    \this_vram.mem_mem_3_0_physical_WADDR_wire\ <= \N__5695\&\N__7372\&\N__7156\&\N__6949\&\N__6745\&\N__6535\&\N__6319\&\N__6112\&\N__5893\&\N__5497\&\N__5278\;
    \this_vram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7748\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7565\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_3\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_2\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_1_physical_RADDR_wire\ <= \N__8956\&\N__9175\&\N__9394\&\N__9601\&\N__9862\&\N__10069\&\N__11107\&\N__11344\&\N__11578\&\N__12355\&\N__12619\;
    \this_vram.mem_mem_3_1_physical_WADDR_wire\ <= \N__5683\&\N__7360\&\N__7144\&\N__6937\&\N__6733\&\N__6523\&\N__6307\&\N__6100\&\N__5881\&\N__5485\&\N__5266\;
    \this_vram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4907\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4808\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_5\ <= \this_vram.mem_mem_3_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_4\ <= \this_vram.mem_mem_3_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_2_physical_RADDR_wire\ <= \N__8944\&\N__9163\&\N__9382\&\N__9589\&\N__9850\&\N__10057\&\N__11095\&\N__11332\&\N__11566\&\N__12343\&\N__12607\;
    \this_vram.mem_mem_3_2_physical_WADDR_wire\ <= \N__5671\&\N__7348\&\N__7132\&\N__6925\&\N__6721\&\N__6511\&\N__6295\&\N__6088\&\N__5869\&\N__5473\&\N__5254\;
    \this_vram.mem_mem_3_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5117\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5025\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_1\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_0\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_0_physical_RADDR_wire\ <= \N__8932\&\N__9151\&\N__9370\&\N__9577\&\N__9838\&\N__10045\&\N__11083\&\N__11320\&\N__11554\&\N__12331\&\N__12595\;
    \this_vram.mem_mem_4_0_physical_WADDR_wire\ <= \N__5659\&\N__7336\&\N__7120\&\N__6913\&\N__6709\&\N__6499\&\N__6283\&\N__6076\&\N__5857\&\N__5461\&\N__5242\;
    \this_vram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7713\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7533\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_3\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_2\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_1_physical_RADDR_wire\ <= \N__8920\&\N__9139\&\N__9358\&\N__9565\&\N__9826\&\N__10033\&\N__11071\&\N__11308\&\N__11542\&\N__12319\&\N__12583\;
    \this_vram.mem_mem_4_1_physical_WADDR_wire\ <= \N__5647\&\N__7324\&\N__7108\&\N__6901\&\N__6697\&\N__6487\&\N__6271\&\N__6064\&\N__5845\&\N__5449\&\N__5230\;
    \this_vram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4926\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4784\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_5\ <= \this_vram.mem_mem_4_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_4\ <= \this_vram.mem_mem_4_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_2_physical_RADDR_wire\ <= \N__8908\&\N__9127\&\N__9346\&\N__9553\&\N__9814\&\N__10021\&\N__11059\&\N__11296\&\N__11530\&\N__12307\&\N__12571\;
    \this_vram.mem_mem_4_2_physical_WADDR_wire\ <= \N__5635\&\N__7312\&\N__7096\&\N__6889\&\N__6685\&\N__6475\&\N__6259\&\N__6052\&\N__5833\&\N__5437\&\N__5218\;
    \this_vram.mem_mem_4_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5118\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5037\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_1\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_0\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_0_physical_RADDR_wire\ <= \N__8896\&\N__9115\&\N__9334\&\N__9541\&\N__9802\&\N__10009\&\N__11047\&\N__11284\&\N__11518\&\N__12295\&\N__12559\;
    \this_vram.mem_mem_5_0_physical_WADDR_wire\ <= \N__5623\&\N__7300\&\N__7084\&\N__6877\&\N__6673\&\N__6463\&\N__6247\&\N__6040\&\N__5821\&\N__5425\&\N__5206\;
    \this_vram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7712\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7509\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_3\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_2\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_1_physical_RADDR_wire\ <= \N__9067\&\N__9286\&\N__9487\&\N__9694\&\N__9955\&\N__10162\&\N__11194\&\N__11431\&\N__11659\&\N__12454\&\N__12712\;
    \this_vram.mem_mem_5_1_physical_WADDR_wire\ <= \N__5776\&\N__7441\&\N__7243\&\N__7030\&\N__6814\&\N__6604\&\N__6394\&\N__6187\&\N__5986\&\N__5560\&\N__5371\;
    \this_vram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4955\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4815\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_5\ <= \this_vram.mem_mem_5_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_4\ <= \this_vram.mem_mem_5_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_2_physical_RADDR_wire\ <= \N__9055\&\N__9274\&\N__9475\&\N__9682\&\N__9943\&\N__10150\&\N__11182\&\N__11419\&\N__11647\&\N__12442\&\N__12700\;
    \this_vram.mem_mem_5_2_physical_WADDR_wire\ <= \N__5764\&\N__7429\&\N__7231\&\N__7018\&\N__6802\&\N__6592\&\N__6382\&\N__6175\&\N__5974\&\N__5548\&\N__5359\;
    \this_vram.mem_mem_5_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5171\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5029\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_1\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_0\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_0_physical_RADDR_wire\ <= \N__9043\&\N__9262\&\N__9463\&\N__9670\&\N__9931\&\N__10138\&\N__11170\&\N__11407\&\N__11635\&\N__12430\&\N__12688\;
    \this_vram.mem_mem_6_0_physical_WADDR_wire\ <= \N__5752\&\N__7417\&\N__7219\&\N__7006\&\N__6790\&\N__6580\&\N__6370\&\N__6163\&\N__5962\&\N__5536\&\N__5347\;
    \this_vram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7772\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7628\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_3\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_2\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_1_physical_RADDR_wire\ <= \N__9031\&\N__9250\&\N__9451\&\N__9658\&\N__9919\&\N__10126\&\N__11158\&\N__11395\&\N__11623\&\N__12418\&\N__12676\;
    \this_vram.mem_mem_6_1_physical_WADDR_wire\ <= \N__5740\&\N__7405\&\N__7207\&\N__6994\&\N__6778\&\N__6568\&\N__6358\&\N__6151\&\N__5950\&\N__5524\&\N__5335\;
    \this_vram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4944\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4804\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_5\ <= \this_vram.mem_mem_6_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_4\ <= \this_vram.mem_mem_6_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_2_physical_RADDR_wire\ <= \N__9019\&\N__9238\&\N__9439\&\N__9646\&\N__9907\&\N__10114\&\N__11146\&\N__11383\&\N__11611\&\N__12406\&\N__12664\;
    \this_vram.mem_mem_6_2_physical_WADDR_wire\ <= \N__5728\&\N__7393\&\N__7195\&\N__6982\&\N__6766\&\N__6556\&\N__6346\&\N__6139\&\N__5938\&\N__5512\&\N__5323\;
    \this_vram.mem_mem_6_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5164\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5050\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_1\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_0\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_0_physical_RADDR_wire\ <= \N__9007\&\N__9226\&\N__9427\&\N__9634\&\N__9895\&\N__10102\&\N__11134\&\N__11371\&\N__11599\&\N__12394\&\N__12652\;
    \this_vram.mem_mem_7_0_physical_WADDR_wire\ <= \N__5716\&\N__7381\&\N__7183\&\N__6970\&\N__6754\&\N__6544\&\N__6334\&\N__6127\&\N__5926\&\N__5500\&\N__5311\;
    \this_vram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7771\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7624\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_3\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_2\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_1_physical_RADDR_wire\ <= \N__8995\&\N__9214\&\N__9415\&\N__9622\&\N__9883\&\N__10090\&\N__11122\&\N__11359\&\N__11587\&\N__12382\&\N__12640\;
    \this_vram.mem_mem_7_1_physical_WADDR_wire\ <= \N__5704\&\N__7369\&\N__7171\&\N__6958\&\N__6742\&\N__6532\&\N__6322\&\N__6115\&\N__5914\&\N__5488\&\N__5299\;
    \this_vram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4920\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4778\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_5\ <= \this_vram.mem_mem_7_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_4\ <= \this_vram.mem_mem_7_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_2_physical_RADDR_wire\ <= \N__8983\&\N__9202\&\N__9403\&\N__9610\&\N__9871\&\N__10078\&\N__11110\&\N__11347\&\N__11575\&\N__12370\&\N__12628\;
    \this_vram.mem_mem_7_2_physical_WADDR_wire\ <= \N__5692\&\N__7357\&\N__7159\&\N__6946\&\N__6730\&\N__6520\&\N__6310\&\N__6103\&\N__5902\&\N__5476\&\N__5287\;
    \this_vram.mem_mem_7_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5157\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5043\&'0'&'0'&'0';
    \this_vram.mem_out_bus8_1\ <= \this_vram.mem_mem_8_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus8_0\ <= \this_vram.mem_mem_8_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_8_0_physical_RADDR_wire\ <= \N__8971\&\N__9190\&\N__9391\&\N__9598\&\N__9859\&\N__10066\&\N__11098\&\N__11335\&\N__11563\&\N__12358\&\N__12616\;
    \this_vram.mem_mem_8_0_physical_WADDR_wire\ <= \N__5680\&\N__7345\&\N__7147\&\N__6934\&\N__6718\&\N__6508\&\N__6298\&\N__6091\&\N__5890\&\N__5464\&\N__5275\;
    \this_vram.mem_mem_8_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_8_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7766\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7614\&'0'&'0'&'0';
    \this_vram.mem_out_bus8_3\ <= \this_vram.mem_mem_8_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus8_2\ <= \this_vram.mem_mem_8_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_8_1_physical_RADDR_wire\ <= \N__8959\&\N__9178\&\N__9379\&\N__9586\&\N__9847\&\N__10054\&\N__11086\&\N__11323\&\N__11551\&\N__12346\&\N__12604\;
    \this_vram.mem_mem_8_1_physical_WADDR_wire\ <= \N__5668\&\N__7333\&\N__7135\&\N__6922\&\N__6706\&\N__6496\&\N__6286\&\N__6079\&\N__5878\&\N__5452\&\N__5263\;
    \this_vram.mem_mem_8_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_8_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4878\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4765\&'0'&'0'&'0';
    \this_vram.mem_out_bus8_5\ <= \this_vram.mem_mem_8_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus8_4\ <= \this_vram.mem_mem_8_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_8_2_physical_RADDR_wire\ <= \N__8947\&\N__9166\&\N__9367\&\N__9574\&\N__9835\&\N__10042\&\N__11074\&\N__11311\&\N__11539\&\N__12334\&\N__12592\;
    \this_vram.mem_mem_8_2_physical_WADDR_wire\ <= \N__5656\&\N__7321\&\N__7123\&\N__6910\&\N__6694\&\N__6484\&\N__6274\&\N__6067\&\N__5866\&\N__5440\&\N__5251\;
    \this_vram.mem_mem_8_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_8_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5144\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5065\&'0'&'0'&'0';
    \this_vram.mem_out_bus9_1\ <= \this_vram.mem_mem_9_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus9_0\ <= \this_vram.mem_mem_9_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_9_0_physical_RADDR_wire\ <= \N__8935\&\N__9154\&\N__9355\&\N__9562\&\N__9823\&\N__10030\&\N__11062\&\N__11299\&\N__11527\&\N__12322\&\N__12580\;
    \this_vram.mem_mem_9_0_physical_WADDR_wire\ <= \N__5644\&\N__7309\&\N__7111\&\N__6898\&\N__6682\&\N__6472\&\N__6262\&\N__6055\&\N__5854\&\N__5428\&\N__5239\;
    \this_vram.mem_mem_9_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_9_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__7770\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7600\&'0'&'0'&'0';
    \this_vram.mem_out_bus9_3\ <= \this_vram.mem_mem_9_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus9_2\ <= \this_vram.mem_mem_9_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_9_1_physical_RADDR_wire\ <= \N__8923\&\N__9142\&\N__9343\&\N__9550\&\N__9811\&\N__10018\&\N__11050\&\N__11287\&\N__11515\&\N__12310\&\N__12568\;
    \this_vram.mem_mem_9_1_physical_WADDR_wire\ <= \N__5632\&\N__7297\&\N__7099\&\N__6886\&\N__6670\&\N__6460\&\N__6250\&\N__6043\&\N__5842\&\N__5416\&\N__5227\;
    \this_vram.mem_mem_9_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_9_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4919\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4743\&'0'&'0'&'0';
    \this_vram.mem_out_bus9_5\ <= \this_vram.mem_mem_9_2_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus9_4\ <= \this_vram.mem_mem_9_2_physical_RDATA_wire\(3);
    \this_vram.mem_mem_9_2_physical_RADDR_wire\ <= \N__8911\&\N__9130\&\N__9331\&\N__9538\&\N__9799\&\N__10006\&\N__11038\&\N__11275\&\N__11503\&\N__12298\&\N__12556\;
    \this_vram.mem_mem_9_2_physical_WADDR_wire\ <= \N__5620\&\N__7285\&\N__7087\&\N__6874\&\N__6658\&\N__6448\&\N__6238\&\N__6031\&\N__5830\&\N__5404\&\N__5215\;
    \this_vram.mem_mem_9_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_9_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__5156\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5069\&'0'&'0'&'0';

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13655\,
            RE => \N__13208\,
            WCLKE => \N__8459\,
            WCLK => \N__13656\,
            WE => \N__13146\
        );

    \this_vram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13659\,
            RE => \N__13171\,
            WCLKE => \N__8458\,
            WCLK => \N__13660\,
            WE => \N__13131\
        );

    \this_vram.mem_mem_0_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13663\,
            RE => \N__13016\,
            WCLKE => \N__8451\,
            WCLK => \N__13664\,
            WE => \N__13110\
        );

    \this_vram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13667\,
            RE => \N__13194\,
            WCLKE => \N__8534\,
            WCLK => \N__13668\,
            WE => \N__13114\
        );

    \this_vram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13675\,
            RE => \N__13265\,
            WCLKE => \N__8533\,
            WCLK => \N__13674\,
            WE => \N__13172\
        );

    \this_vram.mem_mem_1_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13683\,
            RE => \N__13266\,
            WCLKE => \N__8526\,
            WCLK => \N__13684\,
            WE => \N__13173\
        );

    \this_vram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13690\,
            RE => \N__13237\,
            WCLKE => \N__8342\,
            WCLK => \N__13691\,
            WE => \N__13238\
        );

    \this_vram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13696\,
            RE => \N__13332\,
            WCLKE => \N__8338\,
            WCLK => \N__13697\,
            WE => \N__13239\
        );

    \this_vram.mem_mem_2_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13700\,
            RE => \N__13379\,
            WCLKE => \N__8337\,
            WCLK => \N__13701\,
            WE => \N__13300\
        );

    \this_vram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13704\,
            RE => \N__13380\,
            WCLKE => \N__8643\,
            WCLK => \N__13705\,
            WE => \N__13301\
        );

    \this_vram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13708\,
            RE => \N__13352\,
            WCLKE => \N__8644\,
            WCLK => \N__13709\,
            WE => \N__13353\
        );

    \this_vram.mem_mem_3_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13712\,
            RE => \N__13378\,
            WCLKE => \N__8648\,
            WCLK => \N__13713\,
            WE => \N__13354\
        );

    \this_vram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13716\,
            RE => \N__13384\,
            WCLKE => \N__8802\,
            WCLK => \N__13717\,
            WE => \N__13385\
        );

    \this_vram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13720\,
            RE => \N__13396\,
            WCLKE => \N__8803\,
            WCLK => \N__13721\,
            WE => \N__13386\
        );

    \this_vram.mem_mem_4_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13724\,
            RE => \N__13400\,
            WCLKE => \N__8807\,
            WCLK => \N__13725\,
            WE => \N__13401\
        );

    \this_vram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13726\,
            RE => \N__13403\,
            WCLKE => \N__13446\,
            WCLK => \N__13727\,
            WE => \N__13402\
        );

    \this_vram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13657\,
            RE => \N__13049\,
            WCLKE => \N__13451\,
            WCLK => \N__13658\,
            WE => \N__12997\
        );

    \this_vram.mem_mem_5_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13661\,
            RE => \N__12979\,
            WCLKE => \N__13447\,
            WCLK => \N__13662\,
            WE => \N__12993\
        );

    \this_vram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13665\,
            RE => \N__12897\,
            WCLKE => \N__14255\,
            WCLK => \N__13666\,
            WE => \N__12934\
        );

    \this_vram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13670\,
            RE => \N__12954\,
            WCLKE => \N__14254\,
            WCLK => \N__13671\,
            WE => \N__13030\
        );

    \this_vram.mem_mem_6_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13680\,
            RE => \N__12955\,
            WCLKE => \N__14247\,
            WCLK => \N__13679\,
            WE => \N__13087\
        );

    \this_vram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13686\,
            RE => \N__13149\,
            WCLKE => \N__13994\,
            WCLK => \N__13687\,
            WE => \N__13088\
        );

    \this_vram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13694\,
            RE => \N__13150\,
            WCLKE => \N__13993\,
            WCLK => \N__13695\,
            WE => \N__13147\
        );

    \this_vram.mem_mem_7_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13698\,
            RE => \N__13209\,
            WCLKE => \N__13992\,
            WCLK => \N__13699\,
            WE => \N__13148\
        );

    \this_vram.mem_mem_8_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_8_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_8_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_8_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_8_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_8_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13702\,
            RE => \N__13210\,
            WCLKE => \N__14543\,
            WCLK => \N__13703\,
            WE => \N__13276\
        );

    \this_vram.mem_mem_8_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_8_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_8_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_8_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_8_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_8_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13706\,
            RE => \N__13278\,
            WCLKE => \N__14535\,
            WCLK => \N__13707\,
            WE => \N__13277\
        );

    \this_vram.mem_mem_8_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_8_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_8_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_8_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_8_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_8_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13710\,
            RE => \N__13279\,
            WCLKE => \N__14542\,
            WCLK => \N__13711\,
            WE => \N__13339\
        );

    \this_vram.mem_mem_9_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_9_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_9_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_9_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_9_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_9_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13714\,
            RE => \N__13347\,
            WCLKE => \N__14919\,
            WCLK => \N__13715\,
            WE => \N__13340\
        );

    \this_vram.mem_mem_9_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_9_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_9_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_9_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_9_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_9_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13718\,
            RE => \N__13348\,
            WCLKE => \N__14926\,
            WCLK => \N__13719\,
            WE => \N__13381\
        );

    \this_vram.mem_mem_9_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_9_2_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_9_2_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_9_2_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_9_2_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_9_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13722\,
            RE => \N__13383\,
            WCLKE => \N__14927\,
            WCLK => \N__13723\,
            WE => \N__13382\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__15243\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15245\,
            DIN => \N__15244\,
            DOUT => \N__15243\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15245\,
            PADOUT => \N__15244\,
            PADIN => \N__15243\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15234\,
            DIN => \N__15233\,
            DOUT => \N__15232\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15234\,
            PADOUT => \N__15233\,
            PADIN => \N__15232\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7898\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15225\,
            DIN => \N__15224\,
            DOUT => \N__15223\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15225\,
            PADOUT => \N__15224\,
            PADIN => \N__15223\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7910\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15216\,
            DIN => \N__15215\,
            DOUT => \N__15214\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15216\,
            PADOUT => \N__15215\,
            PADIN => \N__15214\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7940\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__7892\
        );

    \rgb_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15207\,
            DIN => \N__15206\,
            DOUT => \N__15205\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15207\,
            PADOUT => \N__15206\,
            PADIN => \N__15205\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8699\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__7845\
        );

    \rgb_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15198\,
            DIN => \N__15197\,
            DOUT => \N__15196\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15198\,
            PADOUT => \N__15197\,
            PADIN => \N__15196\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8351\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__7846\
        );

    \rgb_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15189\,
            DIN => \N__15188\,
            DOUT => \N__15187\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15189\,
            PADOUT => \N__15188\,
            PADIN => \N__15187\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8216\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__7877\
        );

    \rgb_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15180\,
            DIN => \N__15179\,
            DOUT => \N__15178\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15180\,
            PADOUT => \N__15179\,
            PADIN => \N__15178\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8243\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__7888\
        );

    \rgb_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15171\,
            DIN => \N__15170\,
            DOUT => \N__15169\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15171\,
            PADOUT => \N__15170\,
            PADIN => \N__15169\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8270\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__7887\
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15162\,
            DIN => \N__15161\,
            DOUT => \N__15160\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15162\,
            PADOUT => \N__15161\,
            PADIN => \N__15160\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15153\,
            DIN => \N__15152\,
            DOUT => \N__15151\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15153\,
            PADOUT => \N__15152\,
            PADIN => \N__15151\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7823\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15144\,
            DIN => \N__15143\,
            DOUT => \N__15142\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15144\,
            PADOUT => \N__15143\,
            PADIN => \N__15142\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7829\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15135\,
            DIN => \N__15134\,
            DOUT => \N__15133\,
            PACKAGEPIN => write_address_wire(0)
        );

    \write_address_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15135\,
            PADOUT => \N__15134\,
            PADIN => \N__15133\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15126\,
            DIN => \N__15125\,
            DOUT => \N__15124\,
            PACKAGEPIN => write_address_wire(1)
        );

    \write_address_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15126\,
            PADOUT => \N__15125\,
            PADIN => \N__15124\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15117\,
            DIN => \N__15116\,
            DOUT => \N__15115\,
            PACKAGEPIN => write_address_wire(10)
        );

    \write_address_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15117\,
            PADOUT => \N__15116\,
            PADIN => \N__15115\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_10,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15108\,
            DIN => \N__15107\,
            DOUT => \N__15106\,
            PACKAGEPIN => write_address_wire(11)
        );

    \write_address_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15108\,
            PADOUT => \N__15107\,
            PADIN => \N__15106\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_11,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15099\,
            DIN => \N__15098\,
            DOUT => \N__15097\,
            PACKAGEPIN => write_address_wire(12)
        );

    \write_address_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15099\,
            PADOUT => \N__15098\,
            PADIN => \N__15097\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_12,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15090\,
            DIN => \N__15089\,
            DOUT => \N__15088\,
            PACKAGEPIN => write_address_wire(13)
        );

    \write_address_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15090\,
            PADOUT => \N__15089\,
            PADIN => \N__15088\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_13,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15081\,
            DIN => \N__15080\,
            DOUT => \N__15079\,
            PACKAGEPIN => write_address_wire(14)
        );

    \write_address_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15081\,
            PADOUT => \N__15080\,
            PADIN => \N__15079\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_14,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15072\,
            DIN => \N__15071\,
            DOUT => \N__15070\,
            PACKAGEPIN => write_address_wire(2)
        );

    \write_address_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15072\,
            PADOUT => \N__15071\,
            PADIN => \N__15070\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15063\,
            DIN => \N__15062\,
            DOUT => \N__15061\,
            PACKAGEPIN => write_address_wire(3)
        );

    \write_address_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15063\,
            PADOUT => \N__15062\,
            PADIN => \N__15061\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15054\,
            DIN => \N__15053\,
            DOUT => \N__15052\,
            PACKAGEPIN => write_address_wire(4)
        );

    \write_address_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15054\,
            PADOUT => \N__15053\,
            PADIN => \N__15052\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15045\,
            DIN => \N__15044\,
            DOUT => \N__15043\,
            PACKAGEPIN => write_address_wire(5)
        );

    \write_address_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15045\,
            PADOUT => \N__15044\,
            PADIN => \N__15043\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15036\,
            DIN => \N__15035\,
            DOUT => \N__15034\,
            PACKAGEPIN => write_address_wire(6)
        );

    \write_address_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15036\,
            PADOUT => \N__15035\,
            PADIN => \N__15034\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15027\,
            DIN => \N__15026\,
            DOUT => \N__15025\,
            PACKAGEPIN => write_address_wire(7)
        );

    \write_address_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15027\,
            PADOUT => \N__15026\,
            PADIN => \N__15025\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15018\,
            DIN => \N__15017\,
            DOUT => \N__15016\,
            PACKAGEPIN => write_address_wire(8)
        );

    \write_address_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15018\,
            PADOUT => \N__15017\,
            PADIN => \N__15016\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_8,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_address_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15009\,
            DIN => \N__15008\,
            DOUT => \N__15007\,
            PACKAGEPIN => write_address_wire(9)
        );

    \write_address_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15009\,
            PADOUT => \N__15008\,
            PADIN => \N__15007\,
            CLOCKENABLE => 'H',
            DIN0 => write_address_c_9,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15000\,
            DIN => \N__14999\,
            DOUT => \N__14998\,
            PACKAGEPIN => write_data_wire(0)
        );

    \write_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15000\,
            PADOUT => \N__14999\,
            PADIN => \N__14998\,
            CLOCKENABLE => 'H',
            DIN0 => write_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14991\,
            DIN => \N__14990\,
            DOUT => \N__14989\,
            PACKAGEPIN => write_data_wire(1)
        );

    \write_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14991\,
            PADOUT => \N__14990\,
            PADIN => \N__14989\,
            CLOCKENABLE => 'H',
            DIN0 => write_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14982\,
            DIN => \N__14981\,
            DOUT => \N__14980\,
            PACKAGEPIN => write_data_wire(2)
        );

    \write_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14982\,
            PADOUT => \N__14981\,
            PADIN => \N__14980\,
            CLOCKENABLE => 'H',
            DIN0 => write_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14973\,
            DIN => \N__14972\,
            DOUT => \N__14971\,
            PACKAGEPIN => write_data_wire(3)
        );

    \write_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14973\,
            PADOUT => \N__14972\,
            PADIN => \N__14971\,
            CLOCKENABLE => 'H',
            DIN0 => write_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14964\,
            DIN => \N__14963\,
            DOUT => \N__14962\,
            PACKAGEPIN => write_data_wire(4)
        );

    \write_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14964\,
            PADOUT => \N__14963\,
            PADIN => \N__14962\,
            CLOCKENABLE => 'H',
            DIN0 => write_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14955\,
            DIN => \N__14954\,
            DOUT => \N__14953\,
            PACKAGEPIN => write_data_wire(5)
        );

    \write_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14955\,
            PADOUT => \N__14954\,
            PADIN => \N__14953\,
            CLOCKENABLE => 'H',
            DIN0 => write_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \write_en_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14946\,
            DIN => \N__14945\,
            DOUT => \N__14944\,
            PACKAGEPIN => write_en_wire
        );

    \write_en_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14946\,
            PADOUT => \N__14945\,
            PADIN => \N__14944\,
            CLOCKENABLE => 'H',
            DIN0 => write_en_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__3638\ : CEMux
    port map (
            O => \N__14927\,
            I => \N__14923\
        );

    \I__3637\ : CEMux
    port map (
            O => \N__14926\,
            I => \N__14920\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14914\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__14920\,
            I => \N__14914\
        );

    \I__3634\ : CEMux
    port map (
            O => \N__14919\,
            I => \N__14911\
        );

    \I__3633\ : Span4Mux_v
    port map (
            O => \N__14914\,
            I => \N__14906\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__14911\,
            I => \N__14906\
        );

    \I__3631\ : Span4Mux_v
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__14903\,
            I => \this_vram.mem_WE_0\
        );

    \I__3629\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14896\
        );

    \I__3628\ : InMux
    port map (
            O => \N__14899\,
            I => \N__14892\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__14896\,
            I => \N__14889\
        );

    \I__3626\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14886\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__14892\,
            I => \N__14882\
        );

    \I__3624\ : Span4Mux_v
    port map (
            O => \N__14889\,
            I => \N__14877\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__14886\,
            I => \N__14877\
        );

    \I__3622\ : InMux
    port map (
            O => \N__14885\,
            I => \N__14874\
        );

    \I__3621\ : Span4Mux_v
    port map (
            O => \N__14882\,
            I => \N__14871\
        );

    \I__3620\ : Span4Mux_h
    port map (
            O => \N__14877\,
            I => \N__14865\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__14874\,
            I => \N__14865\
        );

    \I__3618\ : Span4Mux_h
    port map (
            O => \N__14871\,
            I => \N__14861\
        );

    \I__3617\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14858\
        );

    \I__3616\ : Span4Mux_v
    port map (
            O => \N__14865\,
            I => \N__14855\
        );

    \I__3615\ : InMux
    port map (
            O => \N__14864\,
            I => \N__14852\
        );

    \I__3614\ : Span4Mux_h
    port map (
            O => \N__14861\,
            I => \N__14847\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__14858\,
            I => \N__14847\
        );

    \I__3612\ : Sp12to4
    port map (
            O => \N__14855\,
            I => \N__14839\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__14852\,
            I => \N__14839\
        );

    \I__3610\ : Span4Mux_v
    port map (
            O => \N__14847\,
            I => \N__14836\
        );

    \I__3609\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14831\
        );

    \I__3608\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14831\
        );

    \I__3607\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14828\
        );

    \I__3606\ : Span12Mux_h
    port map (
            O => \N__14839\,
            I => \N__14825\
        );

    \I__3605\ : Span4Mux_h
    port map (
            O => \N__14836\,
            I => \N__14822\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N__14817\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__14828\,
            I => \N__14817\
        );

    \I__3602\ : Span12Mux_h
    port map (
            O => \N__14825\,
            I => \N__14814\
        );

    \I__3601\ : Sp12to4
    port map (
            O => \N__14822\,
            I => \N__14809\
        );

    \I__3600\ : Span12Mux_v
    port map (
            O => \N__14817\,
            I => \N__14809\
        );

    \I__3599\ : Odrv12
    port map (
            O => \N__14814\,
            I => write_address_c_13
        );

    \I__3598\ : Odrv12
    port map (
            O => \N__14809\,
            I => write_address_c_13
        );

    \I__3597\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14797\
        );

    \I__3596\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14794\
        );

    \I__3595\ : InMux
    port map (
            O => \N__14802\,
            I => \N__14790\
        );

    \I__3594\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14785\
        );

    \I__3593\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14785\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__14797\,
            I => \N__14781\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14778\
        );

    \I__3590\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14775\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__14790\,
            I => \N__14771\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__14785\,
            I => \N__14768\
        );

    \I__3587\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14764\
        );

    \I__3586\ : Span4Mux_v
    port map (
            O => \N__14781\,
            I => \N__14757\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__14778\,
            I => \N__14757\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__14775\,
            I => \N__14757\
        );

    \I__3583\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14754\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__14771\,
            I => \N__14751\
        );

    \I__3581\ : Span4Mux_h
    port map (
            O => \N__14768\,
            I => \N__14748\
        );

    \I__3580\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14745\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__14764\,
            I => \N__14738\
        );

    \I__3578\ : Sp12to4
    port map (
            O => \N__14757\,
            I => \N__14738\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__14754\,
            I => \N__14738\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__14751\,
            I => \N__14735\
        );

    \I__3575\ : Span4Mux_v
    port map (
            O => \N__14748\,
            I => \N__14730\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__14745\,
            I => \N__14730\
        );

    \I__3573\ : Span12Mux_v
    port map (
            O => \N__14738\,
            I => \N__14727\
        );

    \I__3572\ : Sp12to4
    port map (
            O => \N__14735\,
            I => \N__14724\
        );

    \I__3571\ : Span4Mux_v
    port map (
            O => \N__14730\,
            I => \N__14721\
        );

    \I__3570\ : Span12Mux_h
    port map (
            O => \N__14727\,
            I => \N__14718\
        );

    \I__3569\ : Span12Mux_h
    port map (
            O => \N__14724\,
            I => \N__14715\
        );

    \I__3568\ : Span4Mux_h
    port map (
            O => \N__14721\,
            I => \N__14712\
        );

    \I__3567\ : Odrv12
    port map (
            O => \N__14718\,
            I => write_address_c_12
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__14715\,
            I => write_address_c_12
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__14712\,
            I => write_address_c_12
        );

    \I__3564\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14702\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__14702\,
            I => \this_vram.mem_N_29\
        );

    \I__3562\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14690\
        );

    \I__3561\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14690\
        );

    \I__3560\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14690\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__14690\,
            I => \N__14687\
        );

    \I__3558\ : Span12Mux_v
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__3557\ : Odrv12
    port map (
            O => \N__14684\,
            I => write_address_c_14
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__14681\,
            I => \N__14677\
        );

    \I__3555\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14672\
        );

    \I__3554\ : InMux
    port map (
            O => \N__14677\,
            I => \N__14669\
        );

    \I__3553\ : InMux
    port map (
            O => \N__14676\,
            I => \N__14666\
        );

    \I__3552\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14663\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__14672\,
            I => \N__14660\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__14669\,
            I => \N__14656\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__14666\,
            I => \N__14651\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__14663\,
            I => \N__14651\
        );

    \I__3547\ : Span4Mux_v
    port map (
            O => \N__14660\,
            I => \N__14647\
        );

    \I__3546\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14644\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__14656\,
            I => \N__14639\
        );

    \I__3544\ : Span4Mux_v
    port map (
            O => \N__14651\,
            I => \N__14639\
        );

    \I__3543\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14636\
        );

    \I__3542\ : Span4Mux_v
    port map (
            O => \N__14647\,
            I => \N__14631\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__14644\,
            I => \N__14631\
        );

    \I__3540\ : Sp12to4
    port map (
            O => \N__14639\,
            I => \N__14626\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__14636\,
            I => \N__14623\
        );

    \I__3538\ : Span4Mux_v
    port map (
            O => \N__14631\,
            I => \N__14620\
        );

    \I__3537\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14615\
        );

    \I__3536\ : InMux
    port map (
            O => \N__14629\,
            I => \N__14615\
        );

    \I__3535\ : Span12Mux_h
    port map (
            O => \N__14626\,
            I => \N__14608\
        );

    \I__3534\ : Sp12to4
    port map (
            O => \N__14623\,
            I => \N__14608\
        );

    \I__3533\ : Span4Mux_v
    port map (
            O => \N__14620\,
            I => \N__14605\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__14615\,
            I => \N__14602\
        );

    \I__3531\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14597\
        );

    \I__3530\ : InMux
    port map (
            O => \N__14613\,
            I => \N__14597\
        );

    \I__3529\ : Span12Mux_v
    port map (
            O => \N__14608\,
            I => \N__14594\
        );

    \I__3528\ : Sp12to4
    port map (
            O => \N__14605\,
            I => \N__14591\
        );

    \I__3527\ : Sp12to4
    port map (
            O => \N__14602\,
            I => \N__14586\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__14597\,
            I => \N__14586\
        );

    \I__3525\ : Span12Mux_h
    port map (
            O => \N__14594\,
            I => \N__14583\
        );

    \I__3524\ : Span12Mux_h
    port map (
            O => \N__14591\,
            I => \N__14578\
        );

    \I__3523\ : Span12Mux_v
    port map (
            O => \N__14586\,
            I => \N__14578\
        );

    \I__3522\ : Odrv12
    port map (
            O => \N__14583\,
            I => write_address_c_11
        );

    \I__3521\ : Odrv12
    port map (
            O => \N__14578\,
            I => write_address_c_11
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__14573\,
            I => \this_vram.mem_N_29_cascade_\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__14570\,
            I => \N__14567\
        );

    \I__3518\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14562\
        );

    \I__3517\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14557\
        );

    \I__3516\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14557\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__14562\,
            I => \N__14552\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__14557\,
            I => \N__14552\
        );

    \I__3513\ : Span12Mux_v
    port map (
            O => \N__14552\,
            I => \N__14549\
        );

    \I__3512\ : Span12Mux_h
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__3511\ : Odrv12
    port map (
            O => \N__14546\,
            I => write_en_c
        );

    \I__3510\ : CEMux
    port map (
            O => \N__14543\,
            I => \N__14539\
        );

    \I__3509\ : CEMux
    port map (
            O => \N__14542\,
            I => \N__14536\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14532\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__14536\,
            I => \N__14529\
        );

    \I__3506\ : CEMux
    port map (
            O => \N__14535\,
            I => \N__14526\
        );

    \I__3505\ : Span4Mux_h
    port map (
            O => \N__14532\,
            I => \N__14521\
        );

    \I__3504\ : Span4Mux_h
    port map (
            O => \N__14529\,
            I => \N__14521\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__14526\,
            I => \N__14518\
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__14521\,
            I => \this_vram.mem_WE_3\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__14518\,
            I => \this_vram.mem_WE_3\
        );

    \I__3500\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14510\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__14510\,
            I => \N__14507\
        );

    \I__3498\ : Span4Mux_v
    port map (
            O => \N__14507\,
            I => \N__14504\
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__14504\,
            I => \this_vram.mem_out_bus9_3\
        );

    \I__3496\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14498\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__14495\,
            I => \this_vram.mem_out_bus8_3\
        );

    \I__3493\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14489\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__14489\,
            I => \N__14486\
        );

    \I__3491\ : Span12Mux_h
    port map (
            O => \N__14486\,
            I => \N__14483\
        );

    \I__3490\ : Odrv12
    port map (
            O => \N__14483\,
            I => \this_vram.mem_mem_8_1_RNI7H021Z0Z_0\
        );

    \I__3489\ : InMux
    port map (
            O => \N__14480\,
            I => \N__14471\
        );

    \I__3488\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14471\
        );

    \I__3487\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14468\
        );

    \I__3486\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14457\
        );

    \I__3485\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14457\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__14471\,
            I => \N__14449\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__14468\,
            I => \N__14446\
        );

    \I__3482\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14443\
        );

    \I__3481\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14440\
        );

    \I__3480\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14437\
        );

    \I__3479\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14432\
        );

    \I__3478\ : InMux
    port map (
            O => \N__14463\,
            I => \N__14426\
        );

    \I__3477\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14426\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__14457\,
            I => \N__14422\
        );

    \I__3475\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14419\
        );

    \I__3474\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14416\
        );

    \I__3473\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14413\
        );

    \I__3472\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14408\
        );

    \I__3471\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14408\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__14449\,
            I => \N__14395\
        );

    \I__3469\ : Span4Mux_v
    port map (
            O => \N__14446\,
            I => \N__14395\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__14443\,
            I => \N__14395\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__14440\,
            I => \N__14395\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14395\
        );

    \I__3465\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14392\
        );

    \I__3464\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14389\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__14432\,
            I => \N__14386\
        );

    \I__3462\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14383\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__14426\,
            I => \N__14380\
        );

    \I__3460\ : InMux
    port map (
            O => \N__14425\,
            I => \N__14377\
        );

    \I__3459\ : Span4Mux_v
    port map (
            O => \N__14422\,
            I => \N__14372\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__14419\,
            I => \N__14372\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__14416\,
            I => \N__14365\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__14413\,
            I => \N__14365\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__14408\,
            I => \N__14365\
        );

    \I__3454\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14362\
        );

    \I__3453\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14358\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__14395\,
            I => \N__14354\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__14392\,
            I => \N__14349\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__14389\,
            I => \N__14349\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__14386\,
            I => \N__14344\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__14383\,
            I => \N__14344\
        );

    \I__3447\ : Span4Mux_h
    port map (
            O => \N__14380\,
            I => \N__14339\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__14377\,
            I => \N__14339\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__14372\,
            I => \N__14334\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__14365\,
            I => \N__14334\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__14362\,
            I => \N__14331\
        );

    \I__3442\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14328\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__14358\,
            I => \N__14325\
        );

    \I__3440\ : InMux
    port map (
            O => \N__14357\,
            I => \N__14322\
        );

    \I__3439\ : Sp12to4
    port map (
            O => \N__14354\,
            I => \N__14319\
        );

    \I__3438\ : Span12Mux_h
    port map (
            O => \N__14349\,
            I => \N__14316\
        );

    \I__3437\ : Span4Mux_v
    port map (
            O => \N__14344\,
            I => \N__14311\
        );

    \I__3436\ : Span4Mux_v
    port map (
            O => \N__14339\,
            I => \N__14311\
        );

    \I__3435\ : Span4Mux_h
    port map (
            O => \N__14334\,
            I => \N__14306\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__14331\,
            I => \N__14306\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__14328\,
            I => \N__14299\
        );

    \I__3432\ : Span12Mux_v
    port map (
            O => \N__14325\,
            I => \N__14299\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__14322\,
            I => \N__14299\
        );

    \I__3430\ : Odrv12
    port map (
            O => \N__14319\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3429\ : Odrv12
    port map (
            O => \N__14316\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__14311\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__14306\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3426\ : Odrv12
    port map (
            O => \N__14299\,
            I => \this_vram.mem_radregZ0Z_11\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__14288\,
            I => \N__14285\
        );

    \I__3424\ : InMux
    port map (
            O => \N__14285\,
            I => \N__14282\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__14282\,
            I => \this_vram.mem_out_bus8_4\
        );

    \I__3422\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14276\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__14276\,
            I => \N__14273\
        );

    \I__3420\ : Sp12to4
    port map (
            O => \N__14273\,
            I => \N__14270\
        );

    \I__3419\ : Odrv12
    port map (
            O => \N__14270\,
            I => \this_vram.mem_out_bus9_4\
        );

    \I__3418\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14264\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__14264\,
            I => \N__14261\
        );

    \I__3416\ : Span12Mux_h
    port map (
            O => \N__14261\,
            I => \N__14258\
        );

    \I__3415\ : Odrv12
    port map (
            O => \N__14258\,
            I => \this_vram.mem_mem_8_2_RNI9HZ0Z021\
        );

    \I__3414\ : CEMux
    port map (
            O => \N__14255\,
            I => \N__14251\
        );

    \I__3413\ : CEMux
    port map (
            O => \N__14254\,
            I => \N__14248\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14242\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__14248\,
            I => \N__14242\
        );

    \I__3410\ : CEMux
    port map (
            O => \N__14247\,
            I => \N__14239\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__14242\,
            I => \N__14234\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__14239\,
            I => \N__14234\
        );

    \I__3407\ : Span4Mux_v
    port map (
            O => \N__14234\,
            I => \N__14231\
        );

    \I__3406\ : Span4Mux_h
    port map (
            O => \N__14231\,
            I => \N__14228\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__14228\,
            I => \this_vram.mem_WE_9\
        );

    \I__3404\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__14222\,
            I => \N__14219\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__14219\,
            I => \this_vram.mem_out_bus7_4\
        );

    \I__3401\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14213\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__3399\ : Span4Mux_v
    port map (
            O => \N__14210\,
            I => \N__14207\
        );

    \I__3398\ : Span4Mux_v
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__14204\,
            I => \this_vram.mem_out_bus5_4\
        );

    \I__3396\ : InMux
    port map (
            O => \N__14201\,
            I => \N__14198\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__14198\,
            I => \N__14195\
        );

    \I__3394\ : Span4Mux_v
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__3393\ : Sp12to4
    port map (
            O => \N__14192\,
            I => \N__14189\
        );

    \I__3392\ : Span12Mux_h
    port map (
            O => \N__14189\,
            I => \N__14186\
        );

    \I__3391\ : Odrv12
    port map (
            O => \N__14186\,
            I => \this_vram.mem_mem_5_2_RNI58RZ0Z11\
        );

    \I__3390\ : InMux
    port map (
            O => \N__14183\,
            I => \N__14180\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__14180\,
            I => \this_vram.mem_out_bus7_5\
        );

    \I__3388\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14165\
        );

    \I__3387\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14162\
        );

    \I__3386\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14158\
        );

    \I__3385\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14153\
        );

    \I__3384\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14150\
        );

    \I__3383\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14145\
        );

    \I__3382\ : InMux
    port map (
            O => \N__14171\,
            I => \N__14145\
        );

    \I__3381\ : InMux
    port map (
            O => \N__14170\,
            I => \N__14142\
        );

    \I__3380\ : InMux
    port map (
            O => \N__14169\,
            I => \N__14134\
        );

    \I__3379\ : InMux
    port map (
            O => \N__14168\,
            I => \N__14134\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__14165\,
            I => \N__14129\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__14162\,
            I => \N__14129\
        );

    \I__3376\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14126\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__14158\,
            I => \N__14123\
        );

    \I__3374\ : InMux
    port map (
            O => \N__14157\,
            I => \N__14120\
        );

    \I__3373\ : InMux
    port map (
            O => \N__14156\,
            I => \N__14117\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__14153\,
            I => \N__14110\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__14150\,
            I => \N__14110\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__14145\,
            I => \N__14110\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__14142\,
            I => \N__14107\
        );

    \I__3368\ : InMux
    port map (
            O => \N__14141\,
            I => \N__14104\
        );

    \I__3367\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14101\
        );

    \I__3366\ : InMux
    port map (
            O => \N__14139\,
            I => \N__14098\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__14134\,
            I => \N__14092\
        );

    \I__3364\ : Span4Mux_v
    port map (
            O => \N__14129\,
            I => \N__14087\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__14126\,
            I => \N__14087\
        );

    \I__3362\ : Span4Mux_h
    port map (
            O => \N__14123\,
            I => \N__14082\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__14120\,
            I => \N__14082\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__14117\,
            I => \N__14079\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__14110\,
            I => \N__14076\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__14107\,
            I => \N__14071\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__14104\,
            I => \N__14071\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__14101\,
            I => \N__14066\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14066\
        );

    \I__3354\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14063\
        );

    \I__3353\ : InMux
    port map (
            O => \N__14096\,
            I => \N__14058\
        );

    \I__3352\ : InMux
    port map (
            O => \N__14095\,
            I => \N__14058\
        );

    \I__3351\ : Span12Mux_v
    port map (
            O => \N__14092\,
            I => \N__14055\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__14087\,
            I => \N__14050\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__14082\,
            I => \N__14050\
        );

    \I__3348\ : Span4Mux_v
    port map (
            O => \N__14079\,
            I => \N__14047\
        );

    \I__3347\ : Span4Mux_h
    port map (
            O => \N__14076\,
            I => \N__14042\
        );

    \I__3346\ : Span4Mux_v
    port map (
            O => \N__14071\,
            I => \N__14042\
        );

    \I__3345\ : Span12Mux_h
    port map (
            O => \N__14066\,
            I => \N__14035\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__14063\,
            I => \N__14035\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__14058\,
            I => \N__14035\
        );

    \I__3342\ : Odrv12
    port map (
            O => \N__14055\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__3341\ : Odrv4
    port map (
            O => \N__14050\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__14047\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__14042\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__3338\ : Odrv12
    port map (
            O => \N__14035\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__3337\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__14021\,
            I => \N__14018\
        );

    \I__3335\ : Sp12to4
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__3334\ : Span12Mux_v
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__3333\ : Odrv12
    port map (
            O => \N__14012\,
            I => \this_vram.mem_out_bus5_5\
        );

    \I__3332\ : InMux
    port map (
            O => \N__14009\,
            I => \N__14006\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__14003\,
            I => \N__14000\
        );

    \I__3329\ : Span4Mux_h
    port map (
            O => \N__14000\,
            I => \N__13997\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__13997\,
            I => \this_vram.mem_mem_5_2_RNI58R11Z0Z_0\
        );

    \I__3327\ : CEMux
    port map (
            O => \N__13994\,
            I => \N__13989\
        );

    \I__3326\ : CEMux
    port map (
            O => \N__13993\,
            I => \N__13986\
        );

    \I__3325\ : CEMux
    port map (
            O => \N__13992\,
            I => \N__13983\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__13989\,
            I => \N__13978\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__13986\,
            I => \N__13978\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__13983\,
            I => \N__13975\
        );

    \I__3321\ : Span4Mux_v
    port map (
            O => \N__13978\,
            I => \N__13972\
        );

    \I__3320\ : Span4Mux_h
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__13972\,
            I => \this_vram.mem_WE_6\
        );

    \I__3318\ : Odrv4
    port map (
            O => \N__13969\,
            I => \this_vram.mem_WE_6\
        );

    \I__3317\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__3315\ : Span4Mux_v
    port map (
            O => \N__13958\,
            I => \N__13955\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__13955\,
            I => \this_vram.mem_out_bus9_0\
        );

    \I__3313\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13949\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__13949\,
            I => \this_vram.mem_out_bus8_0\
        );

    \I__3311\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__3309\ : Span12Mux_v
    port map (
            O => \N__13940\,
            I => \N__13937\
        );

    \I__3308\ : Span12Mux_h
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__3307\ : Odrv12
    port map (
            O => \N__13934\,
            I => \this_vram.mem_mem_8_0_RNI5HZ0Z021\
        );

    \I__3306\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__13928\,
            I => \this_vram.mem_out_bus8_1\
        );

    \I__3304\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13922\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__3302\ : Span4Mux_v
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__13916\,
            I => \this_vram.mem_out_bus9_1\
        );

    \I__3300\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13910\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__3298\ : Sp12to4
    port map (
            O => \N__13907\,
            I => \N__13904\
        );

    \I__3297\ : Span12Mux_h
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__3296\ : Odrv12
    port map (
            O => \N__13901\,
            I => \this_vram.mem_mem_8_0_RNI5H021Z0Z_0\
        );

    \I__3295\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__13895\,
            I => \this_vram.mem_out_bus8_2\
        );

    \I__3293\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__3291\ : Span4Mux_v
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__13883\,
            I => \this_vram.mem_out_bus9_2\
        );

    \I__3289\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__3287\ : Span12Mux_v
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__3286\ : Span12Mux_h
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__3285\ : Odrv12
    port map (
            O => \N__13868\,
            I => \this_vram.mem_mem_8_1_RNI7HZ0Z021\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__13865\,
            I => \N__13861\
        );

    \I__3283\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13855\
        );

    \I__3282\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13852\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__13860\,
            I => \N__13849\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__13859\,
            I => \N__13846\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__13858\,
            I => \N__13843\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__13855\,
            I => \N__13838\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__13852\,
            I => \N__13838\
        );

    \I__3276\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13835\
        );

    \I__3275\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13832\
        );

    \I__3274\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13829\
        );

    \I__3273\ : Span4Mux_v
    port map (
            O => \N__13838\,
            I => \N__13821\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__13835\,
            I => \N__13821\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__13832\,
            I => \N__13821\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__13829\,
            I => \N__13818\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__13828\,
            I => \N__13815\
        );

    \I__3268\ : Span4Mux_v
    port map (
            O => \N__13821\,
            I => \N__13812\
        );

    \I__3267\ : Span4Mux_v
    port map (
            O => \N__13818\,
            I => \N__13809\
        );

    \I__3266\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13806\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__13812\,
            I => \N__13801\
        );

    \I__3264\ : Span4Mux_h
    port map (
            O => \N__13809\,
            I => \N__13798\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__13806\,
            I => \N__13795\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__13805\,
            I => \N__13792\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__13804\,
            I => \N__13789\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__13801\,
            I => \N__13786\
        );

    \I__3259\ : Span4Mux_h
    port map (
            O => \N__13798\,
            I => \N__13781\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__13795\,
            I => \N__13781\
        );

    \I__3257\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13776\
        );

    \I__3256\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13776\
        );

    \I__3255\ : Span4Mux_h
    port map (
            O => \N__13786\,
            I => \N__13773\
        );

    \I__3254\ : Span4Mux_h
    port map (
            O => \N__13781\,
            I => \N__13770\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__13776\,
            I => \N__13767\
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__13773\,
            I => \this_vram.mem_N_27\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__13770\,
            I => \this_vram.mem_N_27\
        );

    \I__3250\ : Odrv12
    port map (
            O => \N__13767\,
            I => \this_vram.mem_N_27\
        );

    \I__3249\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13748\
        );

    \I__3248\ : InMux
    port map (
            O => \N__13759\,
            I => \N__13748\
        );

    \I__3247\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13748\
        );

    \I__3246\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13748\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__13748\,
            I => \N__13745\
        );

    \I__3244\ : Span4Mux_v
    port map (
            O => \N__13745\,
            I => \N__13742\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__13742\,
            I => \N__13739\
        );

    \I__3242\ : Sp12to4
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__3241\ : Odrv12
    port map (
            O => \N__13736\,
            I => rst_n_c
        );

    \I__3240\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13730\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__13730\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__3238\ : ClkMux
    port map (
            O => \N__13727\,
            I => \N__13508\
        );

    \I__3237\ : ClkMux
    port map (
            O => \N__13726\,
            I => \N__13508\
        );

    \I__3236\ : ClkMux
    port map (
            O => \N__13725\,
            I => \N__13508\
        );

    \I__3235\ : ClkMux
    port map (
            O => \N__13724\,
            I => \N__13508\
        );

    \I__3234\ : ClkMux
    port map (
            O => \N__13723\,
            I => \N__13508\
        );

    \I__3233\ : ClkMux
    port map (
            O => \N__13722\,
            I => \N__13508\
        );

    \I__3232\ : ClkMux
    port map (
            O => \N__13721\,
            I => \N__13508\
        );

    \I__3231\ : ClkMux
    port map (
            O => \N__13720\,
            I => \N__13508\
        );

    \I__3230\ : ClkMux
    port map (
            O => \N__13719\,
            I => \N__13508\
        );

    \I__3229\ : ClkMux
    port map (
            O => \N__13718\,
            I => \N__13508\
        );

    \I__3228\ : ClkMux
    port map (
            O => \N__13717\,
            I => \N__13508\
        );

    \I__3227\ : ClkMux
    port map (
            O => \N__13716\,
            I => \N__13508\
        );

    \I__3226\ : ClkMux
    port map (
            O => \N__13715\,
            I => \N__13508\
        );

    \I__3225\ : ClkMux
    port map (
            O => \N__13714\,
            I => \N__13508\
        );

    \I__3224\ : ClkMux
    port map (
            O => \N__13713\,
            I => \N__13508\
        );

    \I__3223\ : ClkMux
    port map (
            O => \N__13712\,
            I => \N__13508\
        );

    \I__3222\ : ClkMux
    port map (
            O => \N__13711\,
            I => \N__13508\
        );

    \I__3221\ : ClkMux
    port map (
            O => \N__13710\,
            I => \N__13508\
        );

    \I__3220\ : ClkMux
    port map (
            O => \N__13709\,
            I => \N__13508\
        );

    \I__3219\ : ClkMux
    port map (
            O => \N__13708\,
            I => \N__13508\
        );

    \I__3218\ : ClkMux
    port map (
            O => \N__13707\,
            I => \N__13508\
        );

    \I__3217\ : ClkMux
    port map (
            O => \N__13706\,
            I => \N__13508\
        );

    \I__3216\ : ClkMux
    port map (
            O => \N__13705\,
            I => \N__13508\
        );

    \I__3215\ : ClkMux
    port map (
            O => \N__13704\,
            I => \N__13508\
        );

    \I__3214\ : ClkMux
    port map (
            O => \N__13703\,
            I => \N__13508\
        );

    \I__3213\ : ClkMux
    port map (
            O => \N__13702\,
            I => \N__13508\
        );

    \I__3212\ : ClkMux
    port map (
            O => \N__13701\,
            I => \N__13508\
        );

    \I__3211\ : ClkMux
    port map (
            O => \N__13700\,
            I => \N__13508\
        );

    \I__3210\ : ClkMux
    port map (
            O => \N__13699\,
            I => \N__13508\
        );

    \I__3209\ : ClkMux
    port map (
            O => \N__13698\,
            I => \N__13508\
        );

    \I__3208\ : ClkMux
    port map (
            O => \N__13697\,
            I => \N__13508\
        );

    \I__3207\ : ClkMux
    port map (
            O => \N__13696\,
            I => \N__13508\
        );

    \I__3206\ : ClkMux
    port map (
            O => \N__13695\,
            I => \N__13508\
        );

    \I__3205\ : ClkMux
    port map (
            O => \N__13694\,
            I => \N__13508\
        );

    \I__3204\ : ClkMux
    port map (
            O => \N__13693\,
            I => \N__13508\
        );

    \I__3203\ : ClkMux
    port map (
            O => \N__13692\,
            I => \N__13508\
        );

    \I__3202\ : ClkMux
    port map (
            O => \N__13691\,
            I => \N__13508\
        );

    \I__3201\ : ClkMux
    port map (
            O => \N__13690\,
            I => \N__13508\
        );

    \I__3200\ : ClkMux
    port map (
            O => \N__13689\,
            I => \N__13508\
        );

    \I__3199\ : ClkMux
    port map (
            O => \N__13688\,
            I => \N__13508\
        );

    \I__3198\ : ClkMux
    port map (
            O => \N__13687\,
            I => \N__13508\
        );

    \I__3197\ : ClkMux
    port map (
            O => \N__13686\,
            I => \N__13508\
        );

    \I__3196\ : ClkMux
    port map (
            O => \N__13685\,
            I => \N__13508\
        );

    \I__3195\ : ClkMux
    port map (
            O => \N__13684\,
            I => \N__13508\
        );

    \I__3194\ : ClkMux
    port map (
            O => \N__13683\,
            I => \N__13508\
        );

    \I__3193\ : ClkMux
    port map (
            O => \N__13682\,
            I => \N__13508\
        );

    \I__3192\ : ClkMux
    port map (
            O => \N__13681\,
            I => \N__13508\
        );

    \I__3191\ : ClkMux
    port map (
            O => \N__13680\,
            I => \N__13508\
        );

    \I__3190\ : ClkMux
    port map (
            O => \N__13679\,
            I => \N__13508\
        );

    \I__3189\ : ClkMux
    port map (
            O => \N__13678\,
            I => \N__13508\
        );

    \I__3188\ : ClkMux
    port map (
            O => \N__13677\,
            I => \N__13508\
        );

    \I__3187\ : ClkMux
    port map (
            O => \N__13676\,
            I => \N__13508\
        );

    \I__3186\ : ClkMux
    port map (
            O => \N__13675\,
            I => \N__13508\
        );

    \I__3185\ : ClkMux
    port map (
            O => \N__13674\,
            I => \N__13508\
        );

    \I__3184\ : ClkMux
    port map (
            O => \N__13673\,
            I => \N__13508\
        );

    \I__3183\ : ClkMux
    port map (
            O => \N__13672\,
            I => \N__13508\
        );

    \I__3182\ : ClkMux
    port map (
            O => \N__13671\,
            I => \N__13508\
        );

    \I__3181\ : ClkMux
    port map (
            O => \N__13670\,
            I => \N__13508\
        );

    \I__3180\ : ClkMux
    port map (
            O => \N__13669\,
            I => \N__13508\
        );

    \I__3179\ : ClkMux
    port map (
            O => \N__13668\,
            I => \N__13508\
        );

    \I__3178\ : ClkMux
    port map (
            O => \N__13667\,
            I => \N__13508\
        );

    \I__3177\ : ClkMux
    port map (
            O => \N__13666\,
            I => \N__13508\
        );

    \I__3176\ : ClkMux
    port map (
            O => \N__13665\,
            I => \N__13508\
        );

    \I__3175\ : ClkMux
    port map (
            O => \N__13664\,
            I => \N__13508\
        );

    \I__3174\ : ClkMux
    port map (
            O => \N__13663\,
            I => \N__13508\
        );

    \I__3173\ : ClkMux
    port map (
            O => \N__13662\,
            I => \N__13508\
        );

    \I__3172\ : ClkMux
    port map (
            O => \N__13661\,
            I => \N__13508\
        );

    \I__3171\ : ClkMux
    port map (
            O => \N__13660\,
            I => \N__13508\
        );

    \I__3170\ : ClkMux
    port map (
            O => \N__13659\,
            I => \N__13508\
        );

    \I__3169\ : ClkMux
    port map (
            O => \N__13658\,
            I => \N__13508\
        );

    \I__3168\ : ClkMux
    port map (
            O => \N__13657\,
            I => \N__13508\
        );

    \I__3167\ : ClkMux
    port map (
            O => \N__13656\,
            I => \N__13508\
        );

    \I__3166\ : ClkMux
    port map (
            O => \N__13655\,
            I => \N__13508\
        );

    \I__3165\ : GlobalMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__3164\ : gio2CtrlBuf
    port map (
            O => \N__13505\,
            I => clk_c_g
        );

    \I__3163\ : InMux
    port map (
            O => \N__13502\,
            I => \N__13499\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__13499\,
            I => \N__13496\
        );

    \I__3161\ : Span12Mux_v
    port map (
            O => \N__13496\,
            I => \N__13493\
        );

    \I__3160\ : Odrv12
    port map (
            O => \N__13493\,
            I => \this_vram.mem_out_bus6_5\
        );

    \I__3159\ : InMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__3157\ : Span4Mux_v
    port map (
            O => \N__13484\,
            I => \N__13481\
        );

    \I__3156\ : Span4Mux_v
    port map (
            O => \N__13481\,
            I => \N__13478\
        );

    \I__3155\ : Sp12to4
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__3154\ : Span12Mux_h
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__3153\ : Odrv12
    port map (
            O => \N__13472\,
            I => \this_vram.mem_out_bus4_5\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__13469\,
            I => \this_vram.mem_mem_4_2_RNI34P11Z0Z_0_cascade_\
        );

    \I__3151\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__13463\,
            I => \N__13460\
        );

    \I__3149\ : Span4Mux_v
    port map (
            O => \N__13460\,
            I => \N__13457\
        );

    \I__3148\ : Sp12to4
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__3147\ : Odrv12
    port map (
            O => \N__13454\,
            I => \this_vram.mem_N_2372\
        );

    \I__3146\ : CEMux
    port map (
            O => \N__13451\,
            I => \N__13448\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__13448\,
            I => \N__13443\
        );

    \I__3144\ : CEMux
    port map (
            O => \N__13447\,
            I => \N__13440\
        );

    \I__3143\ : CEMux
    port map (
            O => \N__13446\,
            I => \N__13437\
        );

    \I__3142\ : Span4Mux_s1_v
    port map (
            O => \N__13443\,
            I => \N__13432\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__13440\,
            I => \N__13432\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__13437\,
            I => \N__13429\
        );

    \I__3139\ : Span4Mux_v
    port map (
            O => \N__13432\,
            I => \N__13426\
        );

    \I__3138\ : Span4Mux_s3_v
    port map (
            O => \N__13429\,
            I => \N__13423\
        );

    \I__3137\ : Sp12to4
    port map (
            O => \N__13426\,
            I => \N__13420\
        );

    \I__3136\ : Sp12to4
    port map (
            O => \N__13423\,
            I => \N__13417\
        );

    \I__3135\ : Span12Mux_h
    port map (
            O => \N__13420\,
            I => \N__13414\
        );

    \I__3134\ : Span12Mux_v
    port map (
            O => \N__13417\,
            I => \N__13411\
        );

    \I__3133\ : Span12Mux_v
    port map (
            O => \N__13414\,
            I => \N__13408\
        );

    \I__3132\ : Odrv12
    port map (
            O => \N__13411\,
            I => \this_vram.mem_WE_12\
        );

    \I__3131\ : Odrv12
    port map (
            O => \N__13408\,
            I => \this_vram.mem_WE_12\
        );

    \I__3130\ : SRMux
    port map (
            O => \N__13403\,
            I => \N__13397\
        );

    \I__3129\ : SRMux
    port map (
            O => \N__13402\,
            I => \N__13393\
        );

    \I__3128\ : SRMux
    port map (
            O => \N__13401\,
            I => \N__13390\
        );

    \I__3127\ : SRMux
    port map (
            O => \N__13400\,
            I => \N__13387\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__13397\,
            I => \N__13375\
        );

    \I__3125\ : SRMux
    port map (
            O => \N__13396\,
            I => \N__13372\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__13393\,
            I => \N__13367\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__13390\,
            I => \N__13367\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__13387\,
            I => \N__13364\
        );

    \I__3121\ : SRMux
    port map (
            O => \N__13386\,
            I => \N__13361\
        );

    \I__3120\ : SRMux
    port map (
            O => \N__13385\,
            I => \N__13358\
        );

    \I__3119\ : SRMux
    port map (
            O => \N__13384\,
            I => \N__13355\
        );

    \I__3118\ : SRMux
    port map (
            O => \N__13383\,
            I => \N__13349\
        );

    \I__3117\ : SRMux
    port map (
            O => \N__13382\,
            I => \N__13344\
        );

    \I__3116\ : SRMux
    port map (
            O => \N__13381\,
            I => \N__13341\
        );

    \I__3115\ : SRMux
    port map (
            O => \N__13380\,
            I => \N__13336\
        );

    \I__3114\ : SRMux
    port map (
            O => \N__13379\,
            I => \N__13333\
        );

    \I__3113\ : SRMux
    port map (
            O => \N__13378\,
            I => \N__13329\
        );

    \I__3112\ : Span4Mux_s3_v
    port map (
            O => \N__13375\,
            I => \N__13326\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__13372\,
            I => \N__13323\
        );

    \I__3110\ : Span4Mux_s3_v
    port map (
            O => \N__13367\,
            I => \N__13314\
        );

    \I__3109\ : Span4Mux_h
    port map (
            O => \N__13364\,
            I => \N__13314\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__13361\,
            I => \N__13314\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__13358\,
            I => \N__13314\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__13355\,
            I => \N__13311\
        );

    \I__3105\ : SRMux
    port map (
            O => \N__13354\,
            I => \N__13308\
        );

    \I__3104\ : SRMux
    port map (
            O => \N__13353\,
            I => \N__13305\
        );

    \I__3103\ : SRMux
    port map (
            O => \N__13352\,
            I => \N__13302\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__13349\,
            I => \N__13297\
        );

    \I__3101\ : SRMux
    port map (
            O => \N__13348\,
            I => \N__13294\
        );

    \I__3100\ : SRMux
    port map (
            O => \N__13347\,
            I => \N__13291\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__13344\,
            I => \N__13286\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__13341\,
            I => \N__13286\
        );

    \I__3097\ : SRMux
    port map (
            O => \N__13340\,
            I => \N__13283\
        );

    \I__3096\ : SRMux
    port map (
            O => \N__13339\,
            I => \N__13280\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__13336\,
            I => \N__13273\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__13333\,
            I => \N__13270\
        );

    \I__3093\ : SRMux
    port map (
            O => \N__13332\,
            I => \N__13267\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__13329\,
            I => \N__13262\
        );

    \I__3091\ : Span4Mux_v
    port map (
            O => \N__13326\,
            I => \N__13249\
        );

    \I__3090\ : Span4Mux_v
    port map (
            O => \N__13323\,
            I => \N__13249\
        );

    \I__3089\ : Span4Mux_v
    port map (
            O => \N__13314\,
            I => \N__13249\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__13311\,
            I => \N__13249\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__13308\,
            I => \N__13249\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__13305\,
            I => \N__13249\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__13302\,
            I => \N__13246\
        );

    \I__3084\ : SRMux
    port map (
            O => \N__13301\,
            I => \N__13243\
        );

    \I__3083\ : SRMux
    port map (
            O => \N__13300\,
            I => \N__13240\
        );

    \I__3082\ : Span4Mux_v
    port map (
            O => \N__13297\,
            I => \N__13230\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__13294\,
            I => \N__13230\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__13291\,
            I => \N__13230\
        );

    \I__3079\ : Span4Mux_v
    port map (
            O => \N__13286\,
            I => \N__13223\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__13283\,
            I => \N__13223\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__13280\,
            I => \N__13223\
        );

    \I__3076\ : SRMux
    port map (
            O => \N__13279\,
            I => \N__13220\
        );

    \I__3075\ : SRMux
    port map (
            O => \N__13278\,
            I => \N__13217\
        );

    \I__3074\ : SRMux
    port map (
            O => \N__13277\,
            I => \N__13214\
        );

    \I__3073\ : SRMux
    port map (
            O => \N__13276\,
            I => \N__13211\
        );

    \I__3072\ : Span4Mux_v
    port map (
            O => \N__13273\,
            I => \N__13201\
        );

    \I__3071\ : Span4Mux_h
    port map (
            O => \N__13270\,
            I => \N__13201\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__13267\,
            I => \N__13201\
        );

    \I__3069\ : SRMux
    port map (
            O => \N__13266\,
            I => \N__13198\
        );

    \I__3068\ : SRMux
    port map (
            O => \N__13265\,
            I => \N__13195\
        );

    \I__3067\ : Span4Mux_v
    port map (
            O => \N__13262\,
            I => \N__13183\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__13249\,
            I => \N__13183\
        );

    \I__3065\ : Span4Mux_h
    port map (
            O => \N__13246\,
            I => \N__13183\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__13243\,
            I => \N__13183\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__13240\,
            I => \N__13183\
        );

    \I__3062\ : SRMux
    port map (
            O => \N__13239\,
            I => \N__13180\
        );

    \I__3061\ : SRMux
    port map (
            O => \N__13238\,
            I => \N__13177\
        );

    \I__3060\ : SRMux
    port map (
            O => \N__13237\,
            I => \N__13174\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__13230\,
            I => \N__13162\
        );

    \I__3058\ : Span4Mux_v
    port map (
            O => \N__13223\,
            I => \N__13162\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__13220\,
            I => \N__13162\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__13217\,
            I => \N__13162\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__13214\,
            I => \N__13157\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__13211\,
            I => \N__13157\
        );

    \I__3053\ : SRMux
    port map (
            O => \N__13210\,
            I => \N__13154\
        );

    \I__3052\ : SRMux
    port map (
            O => \N__13209\,
            I => \N__13151\
        );

    \I__3051\ : SRMux
    port map (
            O => \N__13208\,
            I => \N__13143\
        );

    \I__3050\ : Span4Mux_v
    port map (
            O => \N__13201\,
            I => \N__13138\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__13198\,
            I => \N__13138\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__13195\,
            I => \N__13135\
        );

    \I__3047\ : SRMux
    port map (
            O => \N__13194\,
            I => \N__13132\
        );

    \I__3046\ : Span4Mux_v
    port map (
            O => \N__13183\,
            I => \N__13124\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__13180\,
            I => \N__13124\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__13177\,
            I => \N__13124\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__13174\,
            I => \N__13121\
        );

    \I__3042\ : SRMux
    port map (
            O => \N__13173\,
            I => \N__13118\
        );

    \I__3041\ : SRMux
    port map (
            O => \N__13172\,
            I => \N__13115\
        );

    \I__3040\ : SRMux
    port map (
            O => \N__13171\,
            I => \N__13111\
        );

    \I__3039\ : Span4Mux_v
    port map (
            O => \N__13162\,
            I => \N__13101\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__13157\,
            I => \N__13101\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__13154\,
            I => \N__13101\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__13151\,
            I => \N__13101\
        );

    \I__3035\ : SRMux
    port map (
            O => \N__13150\,
            I => \N__13098\
        );

    \I__3034\ : SRMux
    port map (
            O => \N__13149\,
            I => \N__13095\
        );

    \I__3033\ : SRMux
    port map (
            O => \N__13148\,
            I => \N__13092\
        );

    \I__3032\ : SRMux
    port map (
            O => \N__13147\,
            I => \N__13089\
        );

    \I__3031\ : SRMux
    port map (
            O => \N__13146\,
            I => \N__13081\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__13143\,
            I => \N__13078\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__13138\,
            I => \N__13071\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__13135\,
            I => \N__13071\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__13132\,
            I => \N__13071\
        );

    \I__3026\ : SRMux
    port map (
            O => \N__13131\,
            I => \N__13068\
        );

    \I__3025\ : Span4Mux_v
    port map (
            O => \N__13124\,
            I => \N__13059\
        );

    \I__3024\ : Span4Mux_h
    port map (
            O => \N__13121\,
            I => \N__13059\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__13118\,
            I => \N__13059\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__13115\,
            I => \N__13059\
        );

    \I__3021\ : SRMux
    port map (
            O => \N__13114\,
            I => \N__13056\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13053\
        );

    \I__3019\ : SRMux
    port map (
            O => \N__13110\,
            I => \N__13050\
        );

    \I__3018\ : Span4Mux_v
    port map (
            O => \N__13101\,
            I => \N__13042\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__13098\,
            I => \N__13042\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__13095\,
            I => \N__13042\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__13092\,
            I => \N__13037\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__13089\,
            I => \N__13037\
        );

    \I__3013\ : SRMux
    port map (
            O => \N__13088\,
            I => \N__13034\
        );

    \I__3012\ : SRMux
    port map (
            O => \N__13087\,
            I => \N__13031\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__13086\,
            I => \N__13026\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__13085\,
            I => \N__13022\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__13084\,
            I => \N__13018\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__13081\,
            I => \N__13007\
        );

    \I__3007\ : Span4Mux_h
    port map (
            O => \N__13078\,
            I => \N__13007\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__13071\,
            I => \N__13007\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__13068\,
            I => \N__13007\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__13059\,
            I => \N__12998\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__13056\,
            I => \N__12998\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__13053\,
            I => \N__12998\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__13050\,
            I => \N__12998\
        );

    \I__3000\ : SRMux
    port map (
            O => \N__13049\,
            I => \N__12994\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__13042\,
            I => \N__12990\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__13037\,
            I => \N__12983\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__13034\,
            I => \N__12983\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__13031\,
            I => \N__12983\
        );

    \I__2995\ : SRMux
    port map (
            O => \N__13030\,
            I => \N__12980\
        );

    \I__2994\ : InMux
    port map (
            O => \N__13029\,
            I => \N__12964\
        );

    \I__2993\ : InMux
    port map (
            O => \N__13026\,
            I => \N__12964\
        );

    \I__2992\ : InMux
    port map (
            O => \N__13025\,
            I => \N__12964\
        );

    \I__2991\ : InMux
    port map (
            O => \N__13022\,
            I => \N__12964\
        );

    \I__2990\ : InMux
    port map (
            O => \N__13021\,
            I => \N__12964\
        );

    \I__2989\ : InMux
    port map (
            O => \N__13018\,
            I => \N__12964\
        );

    \I__2988\ : InMux
    port map (
            O => \N__13017\,
            I => \N__12964\
        );

    \I__2987\ : SRMux
    port map (
            O => \N__13016\,
            I => \N__12961\
        );

    \I__2986\ : Span4Mux_v
    port map (
            O => \N__13007\,
            I => \N__12956\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__12998\,
            I => \N__12956\
        );

    \I__2984\ : SRMux
    port map (
            O => \N__12997\,
            I => \N__12951\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__12994\,
            I => \N__12948\
        );

    \I__2982\ : SRMux
    port map (
            O => \N__12993\,
            I => \N__12945\
        );

    \I__2981\ : Span4Mux_h
    port map (
            O => \N__12990\,
            I => \N__12938\
        );

    \I__2980\ : Span4Mux_v
    port map (
            O => \N__12983\,
            I => \N__12938\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__12980\,
            I => \N__12938\
        );

    \I__2978\ : SRMux
    port map (
            O => \N__12979\,
            I => \N__12935\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__12964\,
            I => \N__12931\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__12961\,
            I => \N__12928\
        );

    \I__2975\ : Span4Mux_h
    port map (
            O => \N__12956\,
            I => \N__12925\
        );

    \I__2974\ : SRMux
    port map (
            O => \N__12955\,
            I => \N__12922\
        );

    \I__2973\ : SRMux
    port map (
            O => \N__12954\,
            I => \N__12919\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__12951\,
            I => \N__12912\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__12948\,
            I => \N__12912\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__12945\,
            I => \N__12912\
        );

    \I__2969\ : Span4Mux_v
    port map (
            O => \N__12938\,
            I => \N__12907\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__12935\,
            I => \N__12907\
        );

    \I__2967\ : SRMux
    port map (
            O => \N__12934\,
            I => \N__12904\
        );

    \I__2966\ : Span4Mux_v
    port map (
            O => \N__12931\,
            I => \N__12901\
        );

    \I__2965\ : Span4Mux_h
    port map (
            O => \N__12928\,
            I => \N__12898\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__12925\,
            I => \N__12894\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__12922\,
            I => \N__12885\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__12919\,
            I => \N__12885\
        );

    \I__2961\ : Span4Mux_v
    port map (
            O => \N__12912\,
            I => \N__12885\
        );

    \I__2960\ : Span4Mux_v
    port map (
            O => \N__12907\,
            I => \N__12885\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__12904\,
            I => \N__12882\
        );

    \I__2958\ : Sp12to4
    port map (
            O => \N__12901\,
            I => \N__12879\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__12898\,
            I => \N__12876\
        );

    \I__2956\ : SRMux
    port map (
            O => \N__12897\,
            I => \N__12873\
        );

    \I__2955\ : Span4Mux_h
    port map (
            O => \N__12894\,
            I => \N__12868\
        );

    \I__2954\ : Span4Mux_v
    port map (
            O => \N__12885\,
            I => \N__12868\
        );

    \I__2953\ : Span4Mux_h
    port map (
            O => \N__12882\,
            I => \N__12865\
        );

    \I__2952\ : Span12Mux_v
    port map (
            O => \N__12879\,
            I => \N__12858\
        );

    \I__2951\ : Sp12to4
    port map (
            O => \N__12876\,
            I => \N__12858\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__12873\,
            I => \N__12858\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__12868\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2948\ : Odrv4
    port map (
            O => \N__12865\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2947\ : Odrv12
    port map (
            O => \N__12858\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2946\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__12848\,
            I => \N__12845\
        );

    \I__2944\ : Span4Mux_v
    port map (
            O => \N__12845\,
            I => \N__12842\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__12842\,
            I => \N__12839\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__12839\,
            I => \this_vram.mem_out_bus9_5\
        );

    \I__2941\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12830\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__12830\,
            I => \this_vram.mem_out_bus8_5\
        );

    \I__2938\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12824\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__12824\,
            I => \N__12821\
        );

    \I__2936\ : Span4Mux_v
    port map (
            O => \N__12821\,
            I => \N__12818\
        );

    \I__2935\ : Sp12to4
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__2934\ : Span12Mux_h
    port map (
            O => \N__12815\,
            I => \N__12812\
        );

    \I__2933\ : Odrv12
    port map (
            O => \N__12812\,
            I => \this_vram.mem_mem_8_2_RNI9H021Z0Z_0\
        );

    \I__2932\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__12806\,
            I => \N__12803\
        );

    \I__2930\ : Sp12to4
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__2929\ : Span12Mux_v
    port map (
            O => \N__12800\,
            I => \N__12797\
        );

    \I__2928\ : Odrv12
    port map (
            O => \N__12797\,
            I => \this_vram.mem_out_bus5_2\
        );

    \I__2927\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12791\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__12791\,
            I => \this_vram.mem_out_bus7_2\
        );

    \I__2925\ : InMux
    port map (
            O => \N__12788\,
            I => \N__12785\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__12785\,
            I => \N__12782\
        );

    \I__2923\ : Span4Mux_v
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__2922\ : Sp12to4
    port map (
            O => \N__12779\,
            I => \N__12776\
        );

    \I__2921\ : Span12Mux_h
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__2920\ : Odrv12
    port map (
            O => \N__12773\,
            I => \this_vram.mem_mem_5_1_RNI38RZ0Z11\
        );

    \I__2919\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__12767\,
            I => \N__12764\
        );

    \I__2917\ : Sp12to4
    port map (
            O => \N__12764\,
            I => \N__12761\
        );

    \I__2916\ : Span12Mux_v
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__2915\ : Odrv12
    port map (
            O => \N__12758\,
            I => \this_vram.mem_out_bus5_3\
        );

    \I__2914\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__12752\,
            I => \this_vram.mem_out_bus7_3\
        );

    \I__2912\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__12746\,
            I => \N__12743\
        );

    \I__2910\ : Span12Mux_s11_h
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__2909\ : Span12Mux_h
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__2908\ : Odrv12
    port map (
            O => \N__12737\,
            I => \this_vram.mem_mem_5_1_RNI38R11Z0Z_0\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__12734\,
            I => \this_vga_signals.N_37_cascade_\
        );

    \I__2906\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__12728\,
            I => \this_vga_signals.M_hstate_q_ns_i_i_2_0\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__12725\,
            I => \N__12722\
        );

    \I__2903\ : CascadeBuf
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__12719\,
            I => \N__12716\
        );

    \I__2901\ : CascadeBuf
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__12713\,
            I => \N__12709\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__12712\,
            I => \N__12706\
        );

    \I__2898\ : CascadeBuf
    port map (
            O => \N__12709\,
            I => \N__12703\
        );

    \I__2897\ : CascadeBuf
    port map (
            O => \N__12706\,
            I => \N__12700\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__12703\,
            I => \N__12697\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__12700\,
            I => \N__12694\
        );

    \I__2894\ : CascadeBuf
    port map (
            O => \N__12697\,
            I => \N__12691\
        );

    \I__2893\ : CascadeBuf
    port map (
            O => \N__12694\,
            I => \N__12688\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__12691\,
            I => \N__12685\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__12688\,
            I => \N__12682\
        );

    \I__2890\ : CascadeBuf
    port map (
            O => \N__12685\,
            I => \N__12679\
        );

    \I__2889\ : CascadeBuf
    port map (
            O => \N__12682\,
            I => \N__12676\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__12679\,
            I => \N__12673\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__12676\,
            I => \N__12670\
        );

    \I__2886\ : CascadeBuf
    port map (
            O => \N__12673\,
            I => \N__12667\
        );

    \I__2885\ : CascadeBuf
    port map (
            O => \N__12670\,
            I => \N__12664\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__12667\,
            I => \N__12661\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__12664\,
            I => \N__12658\
        );

    \I__2882\ : CascadeBuf
    port map (
            O => \N__12661\,
            I => \N__12655\
        );

    \I__2881\ : CascadeBuf
    port map (
            O => \N__12658\,
            I => \N__12652\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__12655\,
            I => \N__12649\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__12652\,
            I => \N__12646\
        );

    \I__2878\ : CascadeBuf
    port map (
            O => \N__12649\,
            I => \N__12643\
        );

    \I__2877\ : CascadeBuf
    port map (
            O => \N__12646\,
            I => \N__12640\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__12643\,
            I => \N__12637\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__12640\,
            I => \N__12634\
        );

    \I__2874\ : CascadeBuf
    port map (
            O => \N__12637\,
            I => \N__12631\
        );

    \I__2873\ : CascadeBuf
    port map (
            O => \N__12634\,
            I => \N__12628\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__12631\,
            I => \N__12625\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__12628\,
            I => \N__12622\
        );

    \I__2870\ : CascadeBuf
    port map (
            O => \N__12625\,
            I => \N__12619\
        );

    \I__2869\ : CascadeBuf
    port map (
            O => \N__12622\,
            I => \N__12616\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__12619\,
            I => \N__12613\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__12616\,
            I => \N__12610\
        );

    \I__2866\ : CascadeBuf
    port map (
            O => \N__12613\,
            I => \N__12607\
        );

    \I__2865\ : CascadeBuf
    port map (
            O => \N__12610\,
            I => \N__12604\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__12607\,
            I => \N__12601\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__12604\,
            I => \N__12598\
        );

    \I__2862\ : CascadeBuf
    port map (
            O => \N__12601\,
            I => \N__12595\
        );

    \I__2861\ : CascadeBuf
    port map (
            O => \N__12598\,
            I => \N__12592\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__12595\,
            I => \N__12589\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__12592\,
            I => \N__12586\
        );

    \I__2858\ : CascadeBuf
    port map (
            O => \N__12589\,
            I => \N__12583\
        );

    \I__2857\ : CascadeBuf
    port map (
            O => \N__12586\,
            I => \N__12580\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__12583\,
            I => \N__12577\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__12580\,
            I => \N__12574\
        );

    \I__2854\ : CascadeBuf
    port map (
            O => \N__12577\,
            I => \N__12571\
        );

    \I__2853\ : CascadeBuf
    port map (
            O => \N__12574\,
            I => \N__12568\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__12571\,
            I => \N__12565\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__12568\,
            I => \N__12562\
        );

    \I__2850\ : CascadeBuf
    port map (
            O => \N__12565\,
            I => \N__12559\
        );

    \I__2849\ : CascadeBuf
    port map (
            O => \N__12562\,
            I => \N__12556\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__12559\,
            I => \N__12553\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__12556\,
            I => \N__12550\
        );

    \I__2846\ : InMux
    port map (
            O => \N__12553\,
            I => \N__12547\
        );

    \I__2845\ : InMux
    port map (
            O => \N__12550\,
            I => \N__12544\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__12547\,
            I => \N__12541\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__12544\,
            I => \N__12536\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__12541\,
            I => \N__12533\
        );

    \I__2841\ : InMux
    port map (
            O => \N__12540\,
            I => \N__12530\
        );

    \I__2840\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12527\
        );

    \I__2839\ : Sp12to4
    port map (
            O => \N__12536\,
            I => \N__12524\
        );

    \I__2838\ : Span4Mux_h
    port map (
            O => \N__12533\,
            I => \N__12521\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__12530\,
            I => \N__12515\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__12527\,
            I => \N__12515\
        );

    \I__2835\ : Span12Mux_s6_v
    port map (
            O => \N__12524\,
            I => \N__12512\
        );

    \I__2834\ : Sp12to4
    port map (
            O => \N__12521\,
            I => \N__12509\
        );

    \I__2833\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12506\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__12515\,
            I => \N__12503\
        );

    \I__2831\ : Span12Mux_h
    port map (
            O => \N__12512\,
            I => \N__12498\
        );

    \I__2830\ : Span12Mux_s6_v
    port map (
            O => \N__12509\,
            I => \N__12498\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__12506\,
            I => \M_this_vga_signals_address_0\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__12503\,
            I => \M_this_vga_signals_address_0\
        );

    \I__2827\ : Odrv12
    port map (
            O => \N__12498\,
            I => \M_this_vga_signals_address_0\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__12491\,
            I => \N__12486\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__12490\,
            I => \N__12482\
        );

    \I__2824\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12479\
        );

    \I__2823\ : InMux
    port map (
            O => \N__12486\,
            I => \N__12474\
        );

    \I__2822\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12474\
        );

    \I__2821\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12471\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__12479\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__12474\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__12471\,
            I => \this_vga_signals.M_hcounter_qZ0Z_11\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__12464\,
            I => \N__12461\
        );

    \I__2816\ : CascadeBuf
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__12458\,
            I => \N__12455\
        );

    \I__2814\ : CascadeBuf
    port map (
            O => \N__12455\,
            I => \N__12451\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__12454\,
            I => \N__12448\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__12451\,
            I => \N__12445\
        );

    \I__2811\ : CascadeBuf
    port map (
            O => \N__12448\,
            I => \N__12442\
        );

    \I__2810\ : CascadeBuf
    port map (
            O => \N__12445\,
            I => \N__12439\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__12442\,
            I => \N__12436\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__12439\,
            I => \N__12433\
        );

    \I__2807\ : CascadeBuf
    port map (
            O => \N__12436\,
            I => \N__12430\
        );

    \I__2806\ : CascadeBuf
    port map (
            O => \N__12433\,
            I => \N__12427\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__12430\,
            I => \N__12424\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__12427\,
            I => \N__12421\
        );

    \I__2803\ : CascadeBuf
    port map (
            O => \N__12424\,
            I => \N__12418\
        );

    \I__2802\ : CascadeBuf
    port map (
            O => \N__12421\,
            I => \N__12415\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__12418\,
            I => \N__12412\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__12415\,
            I => \N__12409\
        );

    \I__2799\ : CascadeBuf
    port map (
            O => \N__12412\,
            I => \N__12406\
        );

    \I__2798\ : CascadeBuf
    port map (
            O => \N__12409\,
            I => \N__12403\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__12406\,
            I => \N__12400\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__12403\,
            I => \N__12397\
        );

    \I__2795\ : CascadeBuf
    port map (
            O => \N__12400\,
            I => \N__12394\
        );

    \I__2794\ : CascadeBuf
    port map (
            O => \N__12397\,
            I => \N__12391\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__12394\,
            I => \N__12388\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__12391\,
            I => \N__12385\
        );

    \I__2791\ : CascadeBuf
    port map (
            O => \N__12388\,
            I => \N__12382\
        );

    \I__2790\ : CascadeBuf
    port map (
            O => \N__12385\,
            I => \N__12379\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__12382\,
            I => \N__12376\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__12379\,
            I => \N__12373\
        );

    \I__2787\ : CascadeBuf
    port map (
            O => \N__12376\,
            I => \N__12370\
        );

    \I__2786\ : CascadeBuf
    port map (
            O => \N__12373\,
            I => \N__12367\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__12370\,
            I => \N__12364\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__12367\,
            I => \N__12361\
        );

    \I__2783\ : CascadeBuf
    port map (
            O => \N__12364\,
            I => \N__12358\
        );

    \I__2782\ : CascadeBuf
    port map (
            O => \N__12361\,
            I => \N__12355\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__12358\,
            I => \N__12352\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__12355\,
            I => \N__12349\
        );

    \I__2779\ : CascadeBuf
    port map (
            O => \N__12352\,
            I => \N__12346\
        );

    \I__2778\ : CascadeBuf
    port map (
            O => \N__12349\,
            I => \N__12343\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__12346\,
            I => \N__12340\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__12343\,
            I => \N__12337\
        );

    \I__2775\ : CascadeBuf
    port map (
            O => \N__12340\,
            I => \N__12334\
        );

    \I__2774\ : CascadeBuf
    port map (
            O => \N__12337\,
            I => \N__12331\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__12334\,
            I => \N__12328\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__12331\,
            I => \N__12325\
        );

    \I__2771\ : CascadeBuf
    port map (
            O => \N__12328\,
            I => \N__12322\
        );

    \I__2770\ : CascadeBuf
    port map (
            O => \N__12325\,
            I => \N__12319\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__12322\,
            I => \N__12316\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__12319\,
            I => \N__12313\
        );

    \I__2767\ : CascadeBuf
    port map (
            O => \N__12316\,
            I => \N__12310\
        );

    \I__2766\ : CascadeBuf
    port map (
            O => \N__12313\,
            I => \N__12307\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__12310\,
            I => \N__12304\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__12307\,
            I => \N__12301\
        );

    \I__2763\ : CascadeBuf
    port map (
            O => \N__12304\,
            I => \N__12298\
        );

    \I__2762\ : CascadeBuf
    port map (
            O => \N__12301\,
            I => \N__12295\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__12298\,
            I => \N__12292\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__12295\,
            I => \N__12289\
        );

    \I__2759\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12285\
        );

    \I__2758\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12282\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__12288\,
            I => \N__12279\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__12285\,
            I => \N__12275\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__12282\,
            I => \N__12272\
        );

    \I__2754\ : InMux
    port map (
            O => \N__12279\,
            I => \N__12266\
        );

    \I__2753\ : InMux
    port map (
            O => \N__12278\,
            I => \N__12266\
        );

    \I__2752\ : Span12Mux_h
    port map (
            O => \N__12275\,
            I => \N__12263\
        );

    \I__2751\ : Span12Mux_h
    port map (
            O => \N__12272\,
            I => \N__12260\
        );

    \I__2750\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12257\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__12266\,
            I => \N__12254\
        );

    \I__2748\ : Span12Mux_v
    port map (
            O => \N__12263\,
            I => \N__12251\
        );

    \I__2747\ : Span12Mux_v
    port map (
            O => \N__12260\,
            I => \N__12248\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__12257\,
            I => \M_this_vga_signals_address_1\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__12254\,
            I => \M_this_vga_signals_address_1\
        );

    \I__2744\ : Odrv12
    port map (
            O => \N__12251\,
            I => \M_this_vga_signals_address_1\
        );

    \I__2743\ : Odrv12
    port map (
            O => \N__12248\,
            I => \M_this_vga_signals_address_1\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__12239\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa_0_a2_0_a2_0_cascade_\
        );

    \I__2741\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12230\
        );

    \I__2740\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12230\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__12230\,
            I => \this_vga_signals.N_169_4\
        );

    \I__2738\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12220\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \N__12217\
        );

    \I__2736\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12214\
        );

    \I__2735\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12211\
        );

    \I__2734\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12208\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__12220\,
            I => \N__12205\
        );

    \I__2732\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12202\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__12214\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__12211\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__12208\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__12205\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__12202\,
            I => \this_vga_signals.M_hstate_d_0_sqmuxa\
        );

    \I__2726\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12188\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__12188\,
            I => \N__12184\
        );

    \I__2724\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12181\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__12184\,
            I => \this_vga_signals.N_169\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__12181\,
            I => \this_vga_signals.N_169\
        );

    \I__2721\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12172\
        );

    \I__2720\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12169\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__12172\,
            I => \this_vga_signals.N_42\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__12169\,
            I => \this_vga_signals.N_42\
        );

    \I__2717\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12158\
        );

    \I__2716\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12158\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__12158\,
            I => \this_vga_signals.N_46\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__12155\,
            I => \N__12152\
        );

    \I__2713\ : InMux
    port map (
            O => \N__12152\,
            I => \N__12143\
        );

    \I__2712\ : InMux
    port map (
            O => \N__12151\,
            I => \N__12143\
        );

    \I__2711\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12143\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__12143\,
            I => \this_vga_signals.N_83\
        );

    \I__2709\ : InMux
    port map (
            O => \N__12140\,
            I => \N__12136\
        );

    \I__2708\ : InMux
    port map (
            O => \N__12139\,
            I => \N__12133\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__12136\,
            I => \N__12130\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__12133\,
            I => \N__12127\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__12130\,
            I => \N__12121\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__12127\,
            I => \N__12121\
        );

    \I__2703\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12118\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__12121\,
            I => \N__12115\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__12118\,
            I => \N__12112\
        );

    \I__2700\ : Sp12to4
    port map (
            O => \N__12115\,
            I => \N__12102\
        );

    \I__2699\ : Span12Mux_s5_h
    port map (
            O => \N__12112\,
            I => \N__12102\
        );

    \I__2698\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12099\
        );

    \I__2697\ : InMux
    port map (
            O => \N__12110\,
            I => \N__12090\
        );

    \I__2696\ : InMux
    port map (
            O => \N__12109\,
            I => \N__12090\
        );

    \I__2695\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12090\
        );

    \I__2694\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12090\
        );

    \I__2693\ : Odrv12
    port map (
            O => \N__12102\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__12099\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__12090\,
            I => \this_vga_signals.M_hstate_qZ0Z_1\
        );

    \I__2690\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12080\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__12080\,
            I => \this_vga_signals.N_27\
        );

    \I__2688\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12071\
        );

    \I__2687\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12071\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__12071\,
            I => \N__12067\
        );

    \I__2685\ : IoInMux
    port map (
            O => \N__12070\,
            I => \N__12062\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__12067\,
            I => \N__12059\
        );

    \I__2683\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12056\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__12065\,
            I => \N__12053\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__12062\,
            I => \N__12050\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__12059\,
            I => \N__12047\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__12056\,
            I => \N__12044\
        );

    \I__2678\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12041\
        );

    \I__2677\ : Span12Mux_s11_v
    port map (
            O => \N__12050\,
            I => \N__12038\
        );

    \I__2676\ : Odrv4
    port map (
            O => \N__12047\,
            I => \M_this_reset_cond_out_0\
        );

    \I__2675\ : Odrv12
    port map (
            O => \N__12044\,
            I => \M_this_reset_cond_out_0\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12041\,
            I => \M_this_reset_cond_out_0\
        );

    \I__2673\ : Odrv12
    port map (
            O => \N__12038\,
            I => \M_this_reset_cond_out_0\
        );

    \I__2672\ : InMux
    port map (
            O => \N__12029\,
            I => \N__12026\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__12026\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__2670\ : InMux
    port map (
            O => \N__12023\,
            I => \N__12020\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__12020\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__2668\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12012\
        );

    \I__2667\ : InMux
    port map (
            O => \N__12016\,
            I => \N__12006\
        );

    \I__2666\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12006\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__12012\,
            I => \N__12003\
        );

    \I__2664\ : InMux
    port map (
            O => \N__12011\,
            I => \N__12000\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__12006\,
            I => \N__11997\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__12003\,
            I => \this_vga_signals.N_68\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__12000\,
            I => \this_vga_signals.N_68\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__11997\,
            I => \this_vga_signals.N_68\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11990\,
            I => \bfn_14_20_0_\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11981\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11978\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__11985\,
            I => \N__11975\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11972\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__11981\,
            I => \N__11968\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11978\,
            I => \N__11965\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11962\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__11972\,
            I => \N__11959\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11956\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__11968\,
            I => \N__11951\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__11965\,
            I => \N__11951\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__11962\,
            I => \N__11948\
        );

    \I__2646\ : Span4Mux_h
    port map (
            O => \N__11959\,
            I => \N__11945\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__11956\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__11951\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__11948\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__11945\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__11936\,
            I => \N__11930\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__11935\,
            I => \N__11926\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \N__11923\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11918\
        );

    \I__2637\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11918\
        );

    \I__2636\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11915\
        );

    \I__2635\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11912\
        );

    \I__2634\ : InMux
    port map (
            O => \N__11923\,
            I => \N__11909\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__11918\,
            I => \N__11901\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__11915\,
            I => \N__11898\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__11912\,
            I => \N__11895\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__11909\,
            I => \N__11892\
        );

    \I__2629\ : SRMux
    port map (
            O => \N__11908\,
            I => \N__11873\
        );

    \I__2628\ : SRMux
    port map (
            O => \N__11907\,
            I => \N__11873\
        );

    \I__2627\ : SRMux
    port map (
            O => \N__11906\,
            I => \N__11873\
        );

    \I__2626\ : SRMux
    port map (
            O => \N__11905\,
            I => \N__11873\
        );

    \I__2625\ : SRMux
    port map (
            O => \N__11904\,
            I => \N__11873\
        );

    \I__2624\ : Glb2LocalMux
    port map (
            O => \N__11901\,
            I => \N__11873\
        );

    \I__2623\ : Glb2LocalMux
    port map (
            O => \N__11898\,
            I => \N__11873\
        );

    \I__2622\ : Glb2LocalMux
    port map (
            O => \N__11895\,
            I => \N__11873\
        );

    \I__2621\ : Glb2LocalMux
    port map (
            O => \N__11892\,
            I => \N__11873\
        );

    \I__2620\ : GlobalMux
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__2619\ : gio2CtrlBuf
    port map (
            O => \N__11870\,
            I => \N_112_g\
        );

    \I__2618\ : InMux
    port map (
            O => \N__11867\,
            I => \N__11859\
        );

    \I__2617\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11859\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11856\
        );

    \I__2615\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11853\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__11859\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__11856\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__11853\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11842\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11839\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11842\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__11839\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__11834\,
            I => \N__11829\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__11833\,
            I => \N__11826\
        );

    \I__2605\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11823\
        );

    \I__2604\ : InMux
    port map (
            O => \N__11829\,
            I => \N__11820\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11817\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11823\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__11820\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__11817\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2599\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11806\
        );

    \I__2598\ : InMux
    port map (
            O => \N__11809\,
            I => \N__11803\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__11806\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__11803\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__2595\ : InMux
    port map (
            O => \N__11798\,
            I => \N__11794\
        );

    \I__2594\ : InMux
    port map (
            O => \N__11797\,
            I => \N__11791\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__11794\,
            I => \N__11788\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__11791\,
            I => \N__11785\
        );

    \I__2591\ : Span4Mux_v
    port map (
            O => \N__11788\,
            I => \N__11779\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__11785\,
            I => \N__11779\
        );

    \I__2589\ : InMux
    port map (
            O => \N__11784\,
            I => \N__11776\
        );

    \I__2588\ : Sp12to4
    port map (
            O => \N__11779\,
            I => \N__11771\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__11776\,
            I => \N__11771\
        );

    \I__2586\ : Span12Mux_s10_h
    port map (
            O => \N__11771\,
            I => \N__11764\
        );

    \I__2585\ : InMux
    port map (
            O => \N__11770\,
            I => \N__11757\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11757\
        );

    \I__2583\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11757\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11754\
        );

    \I__2581\ : Odrv12
    port map (
            O => \N__11764\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__11757\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__11754\,
            I => \this_vga_signals.M_hstate_qZ0Z_0\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__11747\,
            I => \N__11741\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__11746\,
            I => \N__11737\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11734\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11731\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11728\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11723\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11737\,
            I => \N__11723\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__11734\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__11731\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11728\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__11723\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__11714\,
            I => \N__11708\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__11713\,
            I => \N__11705\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \N__11701\
        );

    \I__2564\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11698\
        );

    \I__2563\ : InMux
    port map (
            O => \N__11708\,
            I => \N__11695\
        );

    \I__2562\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11690\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11690\
        );

    \I__2560\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11687\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__11698\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__11695\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__11690\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__11687\,
            I => \this_vga_signals.M_hcounter_qZ0Z_10\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__11678\,
            I => \N__11675\
        );

    \I__2554\ : CascadeBuf
    port map (
            O => \N__11675\,
            I => \N__11672\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__11672\,
            I => \N__11669\
        );

    \I__2552\ : CascadeBuf
    port map (
            O => \N__11669\,
            I => \N__11666\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__11666\,
            I => \N__11663\
        );

    \I__2550\ : CascadeBuf
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__11660\,
            I => \N__11656\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__11659\,
            I => \N__11653\
        );

    \I__2547\ : CascadeBuf
    port map (
            O => \N__11656\,
            I => \N__11650\
        );

    \I__2546\ : CascadeBuf
    port map (
            O => \N__11653\,
            I => \N__11647\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__11650\,
            I => \N__11644\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__11647\,
            I => \N__11641\
        );

    \I__2543\ : CascadeBuf
    port map (
            O => \N__11644\,
            I => \N__11638\
        );

    \I__2542\ : CascadeBuf
    port map (
            O => \N__11641\,
            I => \N__11635\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__11638\,
            I => \N__11632\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__11635\,
            I => \N__11629\
        );

    \I__2539\ : CascadeBuf
    port map (
            O => \N__11632\,
            I => \N__11626\
        );

    \I__2538\ : CascadeBuf
    port map (
            O => \N__11629\,
            I => \N__11623\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__11626\,
            I => \N__11620\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__11623\,
            I => \N__11617\
        );

    \I__2535\ : CascadeBuf
    port map (
            O => \N__11620\,
            I => \N__11614\
        );

    \I__2534\ : CascadeBuf
    port map (
            O => \N__11617\,
            I => \N__11611\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__11614\,
            I => \N__11608\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__11611\,
            I => \N__11605\
        );

    \I__2531\ : CascadeBuf
    port map (
            O => \N__11608\,
            I => \N__11602\
        );

    \I__2530\ : CascadeBuf
    port map (
            O => \N__11605\,
            I => \N__11599\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__11602\,
            I => \N__11596\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__11599\,
            I => \N__11593\
        );

    \I__2527\ : CascadeBuf
    port map (
            O => \N__11596\,
            I => \N__11590\
        );

    \I__2526\ : CascadeBuf
    port map (
            O => \N__11593\,
            I => \N__11587\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__11590\,
            I => \N__11584\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__11587\,
            I => \N__11581\
        );

    \I__2523\ : CascadeBuf
    port map (
            O => \N__11584\,
            I => \N__11578\
        );

    \I__2522\ : CascadeBuf
    port map (
            O => \N__11581\,
            I => \N__11575\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__11578\,
            I => \N__11572\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__11575\,
            I => \N__11569\
        );

    \I__2519\ : CascadeBuf
    port map (
            O => \N__11572\,
            I => \N__11566\
        );

    \I__2518\ : CascadeBuf
    port map (
            O => \N__11569\,
            I => \N__11563\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__11566\,
            I => \N__11560\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__11563\,
            I => \N__11557\
        );

    \I__2515\ : CascadeBuf
    port map (
            O => \N__11560\,
            I => \N__11554\
        );

    \I__2514\ : CascadeBuf
    port map (
            O => \N__11557\,
            I => \N__11551\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__11554\,
            I => \N__11548\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__11551\,
            I => \N__11545\
        );

    \I__2511\ : CascadeBuf
    port map (
            O => \N__11548\,
            I => \N__11542\
        );

    \I__2510\ : CascadeBuf
    port map (
            O => \N__11545\,
            I => \N__11539\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__11542\,
            I => \N__11536\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \N__11533\
        );

    \I__2507\ : CascadeBuf
    port map (
            O => \N__11536\,
            I => \N__11530\
        );

    \I__2506\ : CascadeBuf
    port map (
            O => \N__11533\,
            I => \N__11527\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__11530\,
            I => \N__11524\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__11527\,
            I => \N__11521\
        );

    \I__2503\ : CascadeBuf
    port map (
            O => \N__11524\,
            I => \N__11518\
        );

    \I__2502\ : CascadeBuf
    port map (
            O => \N__11521\,
            I => \N__11515\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__11518\,
            I => \N__11512\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__11515\,
            I => \N__11509\
        );

    \I__2499\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11506\
        );

    \I__2498\ : CascadeBuf
    port map (
            O => \N__11509\,
            I => \N__11503\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__11506\,
            I => \N__11500\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__11503\,
            I => \N__11497\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__11500\,
            I => \N__11494\
        );

    \I__2494\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11490\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__11494\,
            I => \N__11487\
        );

    \I__2492\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11482\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__11490\,
            I => \N__11478\
        );

    \I__2490\ : Sp12to4
    port map (
            O => \N__11487\,
            I => \N__11475\
        );

    \I__2489\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11470\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11470\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__11482\,
            I => \N__11467\
        );

    \I__2486\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11464\
        );

    \I__2485\ : Span12Mux_v
    port map (
            O => \N__11478\,
            I => \N__11461\
        );

    \I__2484\ : Span12Mux_v
    port map (
            O => \N__11475\,
            I => \N__11458\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__11470\,
            I => \M_this_vga_signals_address_2\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__11467\,
            I => \M_this_vga_signals_address_2\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11464\,
            I => \M_this_vga_signals_address_2\
        );

    \I__2480\ : Odrv12
    port map (
            O => \N__11461\,
            I => \M_this_vga_signals_address_2\
        );

    \I__2479\ : Odrv12
    port map (
            O => \N__11458\,
            I => \M_this_vga_signals_address_2\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__11447\,
            I => \N__11444\
        );

    \I__2477\ : CascadeBuf
    port map (
            O => \N__11444\,
            I => \N__11441\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__11441\,
            I => \N__11438\
        );

    \I__2475\ : CascadeBuf
    port map (
            O => \N__11438\,
            I => \N__11435\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__11435\,
            I => \N__11432\
        );

    \I__2473\ : CascadeBuf
    port map (
            O => \N__11432\,
            I => \N__11428\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11425\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__11428\,
            I => \N__11422\
        );

    \I__2470\ : CascadeBuf
    port map (
            O => \N__11425\,
            I => \N__11419\
        );

    \I__2469\ : CascadeBuf
    port map (
            O => \N__11422\,
            I => \N__11416\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__11419\,
            I => \N__11413\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__11416\,
            I => \N__11410\
        );

    \I__2466\ : CascadeBuf
    port map (
            O => \N__11413\,
            I => \N__11407\
        );

    \I__2465\ : CascadeBuf
    port map (
            O => \N__11410\,
            I => \N__11404\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__11407\,
            I => \N__11401\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__11404\,
            I => \N__11398\
        );

    \I__2462\ : CascadeBuf
    port map (
            O => \N__11401\,
            I => \N__11395\
        );

    \I__2461\ : CascadeBuf
    port map (
            O => \N__11398\,
            I => \N__11392\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__11395\,
            I => \N__11389\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__11392\,
            I => \N__11386\
        );

    \I__2458\ : CascadeBuf
    port map (
            O => \N__11389\,
            I => \N__11383\
        );

    \I__2457\ : CascadeBuf
    port map (
            O => \N__11386\,
            I => \N__11380\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__11383\,
            I => \N__11377\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__11380\,
            I => \N__11374\
        );

    \I__2454\ : CascadeBuf
    port map (
            O => \N__11377\,
            I => \N__11371\
        );

    \I__2453\ : CascadeBuf
    port map (
            O => \N__11374\,
            I => \N__11368\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__11371\,
            I => \N__11365\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__11368\,
            I => \N__11362\
        );

    \I__2450\ : CascadeBuf
    port map (
            O => \N__11365\,
            I => \N__11359\
        );

    \I__2449\ : CascadeBuf
    port map (
            O => \N__11362\,
            I => \N__11356\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__11359\,
            I => \N__11353\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__11356\,
            I => \N__11350\
        );

    \I__2446\ : CascadeBuf
    port map (
            O => \N__11353\,
            I => \N__11347\
        );

    \I__2445\ : CascadeBuf
    port map (
            O => \N__11350\,
            I => \N__11344\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__11347\,
            I => \N__11341\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__11344\,
            I => \N__11338\
        );

    \I__2442\ : CascadeBuf
    port map (
            O => \N__11341\,
            I => \N__11335\
        );

    \I__2441\ : CascadeBuf
    port map (
            O => \N__11338\,
            I => \N__11332\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__11335\,
            I => \N__11329\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__11332\,
            I => \N__11326\
        );

    \I__2438\ : CascadeBuf
    port map (
            O => \N__11329\,
            I => \N__11323\
        );

    \I__2437\ : CascadeBuf
    port map (
            O => \N__11326\,
            I => \N__11320\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11317\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__11320\,
            I => \N__11314\
        );

    \I__2434\ : CascadeBuf
    port map (
            O => \N__11317\,
            I => \N__11311\
        );

    \I__2433\ : CascadeBuf
    port map (
            O => \N__11314\,
            I => \N__11308\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__11311\,
            I => \N__11305\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__11308\,
            I => \N__11302\
        );

    \I__2430\ : CascadeBuf
    port map (
            O => \N__11305\,
            I => \N__11299\
        );

    \I__2429\ : CascadeBuf
    port map (
            O => \N__11302\,
            I => \N__11296\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__11299\,
            I => \N__11293\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__2426\ : CascadeBuf
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__2425\ : CascadeBuf
    port map (
            O => \N__11290\,
            I => \N__11284\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__11287\,
            I => \N__11281\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__11284\,
            I => \N__11278\
        );

    \I__2422\ : CascadeBuf
    port map (
            O => \N__11281\,
            I => \N__11275\
        );

    \I__2421\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11272\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__11275\,
            I => \N__11269\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__11272\,
            I => \N__11266\
        );

    \I__2418\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11263\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__11266\,
            I => \N__11260\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__11263\,
            I => \N__11256\
        );

    \I__2415\ : Span4Mux_h
    port map (
            O => \N__11260\,
            I => \N__11252\
        );

    \I__2414\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11247\
        );

    \I__2413\ : Span12Mux_s8_h
    port map (
            O => \N__11256\,
            I => \N__11244\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11241\
        );

    \I__2411\ : Sp12to4
    port map (
            O => \N__11252\,
            I => \N__11238\
        );

    \I__2410\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11235\
        );

    \I__2409\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11232\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__11247\,
            I => \N__11229\
        );

    \I__2407\ : Span12Mux_v
    port map (
            O => \N__11244\,
            I => \N__11226\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__11241\,
            I => \N__11221\
        );

    \I__2405\ : Span12Mux_s11_v
    port map (
            O => \N__11238\,
            I => \N__11221\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__11235\,
            I => \M_this_vga_signals_address_3\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__11232\,
            I => \M_this_vga_signals_address_3\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__11229\,
            I => \M_this_vga_signals_address_3\
        );

    \I__2401\ : Odrv12
    port map (
            O => \N__11226\,
            I => \M_this_vga_signals_address_3\
        );

    \I__2400\ : Odrv12
    port map (
            O => \N__11221\,
            I => \M_this_vga_signals_address_3\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__2398\ : CascadeBuf
    port map (
            O => \N__11207\,
            I => \N__11204\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__2396\ : CascadeBuf
    port map (
            O => \N__11201\,
            I => \N__11198\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__2394\ : CascadeBuf
    port map (
            O => \N__11195\,
            I => \N__11191\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__11194\,
            I => \N__11188\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__11191\,
            I => \N__11185\
        );

    \I__2391\ : CascadeBuf
    port map (
            O => \N__11188\,
            I => \N__11182\
        );

    \I__2390\ : CascadeBuf
    port map (
            O => \N__11185\,
            I => \N__11179\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__11182\,
            I => \N__11176\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__11179\,
            I => \N__11173\
        );

    \I__2387\ : CascadeBuf
    port map (
            O => \N__11176\,
            I => \N__11170\
        );

    \I__2386\ : CascadeBuf
    port map (
            O => \N__11173\,
            I => \N__11167\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__11170\,
            I => \N__11164\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__11167\,
            I => \N__11161\
        );

    \I__2383\ : CascadeBuf
    port map (
            O => \N__11164\,
            I => \N__11158\
        );

    \I__2382\ : CascadeBuf
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__11158\,
            I => \N__11152\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__11155\,
            I => \N__11149\
        );

    \I__2379\ : CascadeBuf
    port map (
            O => \N__11152\,
            I => \N__11146\
        );

    \I__2378\ : CascadeBuf
    port map (
            O => \N__11149\,
            I => \N__11143\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__11146\,
            I => \N__11140\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__11143\,
            I => \N__11137\
        );

    \I__2375\ : CascadeBuf
    port map (
            O => \N__11140\,
            I => \N__11134\
        );

    \I__2374\ : CascadeBuf
    port map (
            O => \N__11137\,
            I => \N__11131\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__11134\,
            I => \N__11128\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__11131\,
            I => \N__11125\
        );

    \I__2371\ : CascadeBuf
    port map (
            O => \N__11128\,
            I => \N__11122\
        );

    \I__2370\ : CascadeBuf
    port map (
            O => \N__11125\,
            I => \N__11119\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__11122\,
            I => \N__11116\
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__11119\,
            I => \N__11113\
        );

    \I__2367\ : CascadeBuf
    port map (
            O => \N__11116\,
            I => \N__11110\
        );

    \I__2366\ : CascadeBuf
    port map (
            O => \N__11113\,
            I => \N__11107\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__11110\,
            I => \N__11104\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__11107\,
            I => \N__11101\
        );

    \I__2363\ : CascadeBuf
    port map (
            O => \N__11104\,
            I => \N__11098\
        );

    \I__2362\ : CascadeBuf
    port map (
            O => \N__11101\,
            I => \N__11095\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__11098\,
            I => \N__11092\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__11095\,
            I => \N__11089\
        );

    \I__2359\ : CascadeBuf
    port map (
            O => \N__11092\,
            I => \N__11086\
        );

    \I__2358\ : CascadeBuf
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__11086\,
            I => \N__11080\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__11083\,
            I => \N__11077\
        );

    \I__2355\ : CascadeBuf
    port map (
            O => \N__11080\,
            I => \N__11074\
        );

    \I__2354\ : CascadeBuf
    port map (
            O => \N__11077\,
            I => \N__11071\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__11074\,
            I => \N__11068\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__11071\,
            I => \N__11065\
        );

    \I__2351\ : CascadeBuf
    port map (
            O => \N__11068\,
            I => \N__11062\
        );

    \I__2350\ : CascadeBuf
    port map (
            O => \N__11065\,
            I => \N__11059\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__11062\,
            I => \N__11056\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__11059\,
            I => \N__11053\
        );

    \I__2347\ : CascadeBuf
    port map (
            O => \N__11056\,
            I => \N__11050\
        );

    \I__2346\ : CascadeBuf
    port map (
            O => \N__11053\,
            I => \N__11047\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__11050\,
            I => \N__11044\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__11047\,
            I => \N__11041\
        );

    \I__2343\ : CascadeBuf
    port map (
            O => \N__11044\,
            I => \N__11038\
        );

    \I__2342\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11035\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__11038\,
            I => \N__11032\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__11035\,
            I => \N__11029\
        );

    \I__2339\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11026\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__11029\,
            I => \N__11023\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__11026\,
            I => \N__11019\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__11023\,
            I => \N__11015\
        );

    \I__2335\ : InMux
    port map (
            O => \N__11022\,
            I => \N__11011\
        );

    \I__2334\ : Span12Mux_s9_h
    port map (
            O => \N__11019\,
            I => \N__11007\
        );

    \I__2333\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11004\
        );

    \I__2332\ : Sp12to4
    port map (
            O => \N__11015\,
            I => \N__11001\
        );

    \I__2331\ : InMux
    port map (
            O => \N__11014\,
            I => \N__10998\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__11011\,
            I => \N__10995\
        );

    \I__2329\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10992\
        );

    \I__2328\ : Span12Mux_v
    port map (
            O => \N__11007\,
            I => \N__10989\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__11004\,
            I => \N__10984\
        );

    \I__2326\ : Span12Mux_s10_v
    port map (
            O => \N__11001\,
            I => \N__10984\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10998\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__10995\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10992\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2322\ : Odrv12
    port map (
            O => \N__10989\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2321\ : Odrv12
    port map (
            O => \N__10984\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__10973\,
            I => \N__10970\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__2317\ : Span4Mux_h
    port map (
            O => \N__10964\,
            I => \N__10957\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10954\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10949\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10949\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10946\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__10957\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__10954\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__10949\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10946\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10937\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_6\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__10934\,
            I => \N__10930\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10927\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10930\,
            I => \N__10924\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__10927\,
            I => \N__10919\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10924\,
            I => \N__10915\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10912\
        );

    \I__2301\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10909\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__10919\,
            I => \N__10906\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10903\
        );

    \I__2298\ : Span4Mux_v
    port map (
            O => \N__10915\,
            I => \N__10898\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10912\,
            I => \N__10898\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__10909\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__10906\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__10903\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__10898\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10889\,
            I => \bfn_14_19_0_\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__10883\,
            I => \N__10880\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__10880\,
            I => \this_vga_signals.M_hstate_q_ns_i_i_1_0\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__10877\,
            I => \this_vga_signals.N_76_cascade_\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__10874\,
            I => \this_vga_signals.N_29_cascade_\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10866\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10863\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__10869\,
            I => \N__10859\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__10866\,
            I => \N__10854\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10863\,
            I => \N__10854\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10849\
        );

    \I__2280\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10849\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__10854\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10849\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__10844\,
            I => \N__10839\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__10843\,
            I => \N__10835\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10831\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10828\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10823\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10835\,
            I => \N__10823\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10820\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10831\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10828\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10823\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__10820\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__10805\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_CO\
        );

    \I__2263\ : InMux
    port map (
            O => \N__10802\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_0\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10794\
        );

    \I__2261\ : InMux
    port map (
            O => \N__10798\,
            I => \N__10789\
        );

    \I__2260\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10784\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10794\,
            I => \N__10781\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10778\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10775\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10789\,
            I => \N__10772\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10788\,
            I => \N__10769\
        );

    \I__2254\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10766\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__10784\,
            I => \this_vga_signals.address_1_0\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__10781\,
            I => \this_vga_signals.address_1_0\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__10778\,
            I => \this_vga_signals.address_1_0\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__10775\,
            I => \this_vga_signals.address_1_0\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__10772\,
            I => \this_vga_signals.address_1_0\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__10769\,
            I => \this_vga_signals.address_1_0\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__10766\,
            I => \this_vga_signals.address_1_0\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__10745\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_CO\
        );

    \I__2243\ : InMux
    port map (
            O => \N__10742\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_1\
        );

    \I__2242\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10734\
        );

    \I__2241\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10731\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10724\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__10734\,
            I => \N__10719\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__10731\,
            I => \N__10719\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10714\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10714\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10728\,
            I => \N__10711\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10708\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10724\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__10719\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10714\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__10711\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10708\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__10688\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_CO\
        );

    \I__2224\ : InMux
    port map (
            O => \N__10685\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_2\
        );

    \I__2223\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10677\
        );

    \I__2222\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10672\
        );

    \I__2221\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10672\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10667\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__10672\,
            I => \N__10663\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10671\,
            I => \N__10660\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10657\
        );

    \I__2216\ : Span4Mux_v
    port map (
            O => \N__10667\,
            I => \N__10654\
        );

    \I__2215\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10651\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__10663\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__10660\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__10657\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__10654\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__10651\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__2209\ : InMux
    port map (
            O => \N__10640\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_3\
        );

    \I__2208\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10633\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__10636\,
            I => \N__10627\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__10633\,
            I => \N__10624\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10621\
        );

    \I__2204\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10616\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10616\
        );

    \I__2202\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10613\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__10624\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__10621\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10616\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__10613\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__2197\ : InMux
    port map (
            O => \N__10604\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_4\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__2195\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10595\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__10592\,
            I => \N__10585\
        );

    \I__2192\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10582\
        );

    \I__2191\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10577\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10577\
        );

    \I__2189\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10574\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__10585\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__10582\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__10577\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__10574\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__2184\ : InMux
    port map (
            O => \N__10565\,
            I => \this_vga_signals.un1_M_vcounter_q_6_cry_5\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10562\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__2182\ : InMux
    port map (
            O => \N__10559\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__2181\ : InMux
    port map (
            O => \N__10556\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__2180\ : InMux
    port map (
            O => \N__10553\,
            I => \bfn_14_16_0_\
        );

    \I__2179\ : InMux
    port map (
            O => \N__10550\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_9\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10547\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_10\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \this_vga_signals.N_68_cascade_\
        );

    \I__2176\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10536\
        );

    \I__2175\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10531\
        );

    \I__2174\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10531\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__10536\,
            I => \this_vga_signals.m27_0_a2_1_4\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__10531\,
            I => \this_vga_signals.m27_0_a2_1_4\
        );

    \I__2171\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10523\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__10523\,
            I => \this_vga_signals.M_vcounter_q_0_i_a2_0_0\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__10520\,
            I => \N__10516\
        );

    \I__2168\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10510\
        );

    \I__2167\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10510\
        );

    \I__2166\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10507\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__10510\,
            I => \N__10502\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10502\
        );

    \I__2163\ : Span12Mux_s5_h
    port map (
            O => \N__10502\,
            I => \N__10493\
        );

    \I__2162\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10484\
        );

    \I__2161\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10484\
        );

    \I__2160\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10484\
        );

    \I__2159\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10484\
        );

    \I__2158\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10479\
        );

    \I__2157\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10479\
        );

    \I__2156\ : Odrv12
    port map (
            O => \N__10493\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__10484\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__10479\,
            I => \this_vga_signals.M_vstate_qZ0Z_0\
        );

    \I__2153\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10466\
        );

    \I__2152\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10466\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__10466\,
            I => \N__10458\
        );

    \I__2150\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10455\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__10464\,
            I => \N__10450\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__10463\,
            I => \N__10447\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__10462\,
            I => \N__10444\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__10461\,
            I => \N__10440\
        );

    \I__2145\ : Sp12to4
    port map (
            O => \N__10458\,
            I => \N__10435\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10455\,
            I => \N__10435\
        );

    \I__2143\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10428\
        );

    \I__2142\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10428\
        );

    \I__2141\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10428\
        );

    \I__2140\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10423\
        );

    \I__2139\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10423\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10418\
        );

    \I__2137\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10418\
        );

    \I__2136\ : Odrv12
    port map (
            O => \N__10435\,
            I => \this_vga_signals.M_vstate_qZ0Z_1\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__10428\,
            I => \this_vga_signals.M_vstate_qZ0Z_1\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__10423\,
            I => \this_vga_signals.M_vstate_qZ0Z_1\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__10418\,
            I => \this_vga_signals.M_vstate_qZ0Z_1\
        );

    \I__2132\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__10406\,
            I => \this_vga_signals.m24_0_0\
        );

    \I__2130\ : InMux
    port map (
            O => \N__10403\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__2129\ : InMux
    port map (
            O => \N__10400\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__2128\ : InMux
    port map (
            O => \N__10397\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__2127\ : InMux
    port map (
            O => \N__10394\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__2126\ : InMux
    port map (
            O => \N__10391\,
            I => \this_vga_signals.address_1_0_cry_2\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__2124\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__10379\,
            I => \this_vga_signals.address_1_0_4\
        );

    \I__2121\ : InMux
    port map (
            O => \N__10376\,
            I => \this_vga_signals.address_1_0_cry_3\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \N__10370\
        );

    \I__2119\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__10364\,
            I => \this_vga_signals.address_1_0_5\
        );

    \I__2116\ : InMux
    port map (
            O => \N__10361\,
            I => \this_vga_signals.address_1_0_cry_4\
        );

    \I__2115\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__10352\,
            I => \this_vga_signals.address_1_0_6\
        );

    \I__2112\ : InMux
    port map (
            O => \N__10349\,
            I => \this_vga_signals.address_1_0_cry_5\
        );

    \I__2111\ : InMux
    port map (
            O => \N__10346\,
            I => \N__10343\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__10340\,
            I => \this_vga_signals.address_1_0_7\
        );

    \I__2108\ : InMux
    port map (
            O => \N__10337\,
            I => \this_vga_signals.address_1_0_cry_6\
        );

    \I__2107\ : InMux
    port map (
            O => \N__10334\,
            I => \bfn_13_18_0_\
        );

    \I__2106\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__10325\,
            I => \this_vga_signals.address_1_0_8_THRU_CO\
        );

    \I__2103\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__10319\,
            I => \this_vga_signals.m27_0_o2_0_3\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10313\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__10313\,
            I => \this_vga_signals.N_36\
        );

    \I__2099\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10304\
        );

    \I__2098\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10304\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__10304\,
            I => \this_vga_signals.m27_0_a2_1_5\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__10301\,
            I => \this_vga_signals.m27_0_a2_1_5_cascade_\
        );

    \I__2095\ : InMux
    port map (
            O => \N__10298\,
            I => \this_vga_signals.address_1_cry_4\
        );

    \I__2094\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10290\
        );

    \I__2093\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10287\
        );

    \I__2092\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10284\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__10290\,
            I => \N__10274\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__10287\,
            I => \N__10274\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__10284\,
            I => \N__10274\
        );

    \I__2088\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10270\
        );

    \I__2087\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10267\
        );

    \I__2086\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10264\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__10274\,
            I => \N__10261\
        );

    \I__2084\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10258\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__10270\,
            I => \N__10251\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__10267\,
            I => \N__10251\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10251\
        );

    \I__2080\ : Sp12to4
    port map (
            O => \N__10261\,
            I => \N__10246\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10258\,
            I => \N__10246\
        );

    \I__2078\ : Span4Mux_v
    port map (
            O => \N__10251\,
            I => \N__10243\
        );

    \I__2077\ : Odrv12
    port map (
            O => \N__10246\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__10243\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__2075\ : InMux
    port map (
            O => \N__10238\,
            I => \this_vga_signals.address_1_cry_5\
        );

    \I__2074\ : InMux
    port map (
            O => \N__10235\,
            I => \this_vga_signals.address_1_cry_6\
        );

    \I__2073\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10225\
        );

    \I__2072\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__2071\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10222\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10217\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N__10217\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__10217\,
            I => \N__10211\
        );

    \I__2067\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10208\
        );

    \I__2066\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10203\
        );

    \I__2065\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10203\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__10211\,
            I => \N__10199\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__10208\,
            I => \N__10194\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10194\
        );

    \I__2061\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10191\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__10199\,
            I => \N__10188\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__10194\,
            I => \N__10185\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__10191\,
            I => \N__10182\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__10188\,
            I => \this_vram.mem_radregZ0Z_14\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__10185\,
            I => \this_vram.mem_radregZ0Z_14\
        );

    \I__2055\ : Odrv12
    port map (
            O => \N__10182\,
            I => \this_vram.mem_radregZ0Z_14\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__2053\ : CascadeBuf
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__2051\ : CascadeBuf
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__10163\,
            I => \N__10159\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__10162\,
            I => \N__10156\
        );

    \I__2048\ : CascadeBuf
    port map (
            O => \N__10159\,
            I => \N__10153\
        );

    \I__2047\ : CascadeBuf
    port map (
            O => \N__10156\,
            I => \N__10150\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__10153\,
            I => \N__10147\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__10150\,
            I => \N__10144\
        );

    \I__2044\ : CascadeBuf
    port map (
            O => \N__10147\,
            I => \N__10141\
        );

    \I__2043\ : CascadeBuf
    port map (
            O => \N__10144\,
            I => \N__10138\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__10141\,
            I => \N__10135\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__10138\,
            I => \N__10132\
        );

    \I__2040\ : CascadeBuf
    port map (
            O => \N__10135\,
            I => \N__10129\
        );

    \I__2039\ : CascadeBuf
    port map (
            O => \N__10132\,
            I => \N__10126\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__10129\,
            I => \N__10123\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__10126\,
            I => \N__10120\
        );

    \I__2036\ : CascadeBuf
    port map (
            O => \N__10123\,
            I => \N__10117\
        );

    \I__2035\ : CascadeBuf
    port map (
            O => \N__10120\,
            I => \N__10114\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__10117\,
            I => \N__10111\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__10114\,
            I => \N__10108\
        );

    \I__2032\ : CascadeBuf
    port map (
            O => \N__10111\,
            I => \N__10105\
        );

    \I__2031\ : CascadeBuf
    port map (
            O => \N__10108\,
            I => \N__10102\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__10105\,
            I => \N__10099\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__10102\,
            I => \N__10096\
        );

    \I__2028\ : CascadeBuf
    port map (
            O => \N__10099\,
            I => \N__10093\
        );

    \I__2027\ : CascadeBuf
    port map (
            O => \N__10096\,
            I => \N__10090\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__10093\,
            I => \N__10087\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__10090\,
            I => \N__10084\
        );

    \I__2024\ : CascadeBuf
    port map (
            O => \N__10087\,
            I => \N__10081\
        );

    \I__2023\ : CascadeBuf
    port map (
            O => \N__10084\,
            I => \N__10078\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__10081\,
            I => \N__10075\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__10078\,
            I => \N__10072\
        );

    \I__2020\ : CascadeBuf
    port map (
            O => \N__10075\,
            I => \N__10069\
        );

    \I__2019\ : CascadeBuf
    port map (
            O => \N__10072\,
            I => \N__10066\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__10069\,
            I => \N__10063\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__10066\,
            I => \N__10060\
        );

    \I__2016\ : CascadeBuf
    port map (
            O => \N__10063\,
            I => \N__10057\
        );

    \I__2015\ : CascadeBuf
    port map (
            O => \N__10060\,
            I => \N__10054\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__10057\,
            I => \N__10051\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__10054\,
            I => \N__10048\
        );

    \I__2012\ : CascadeBuf
    port map (
            O => \N__10051\,
            I => \N__10045\
        );

    \I__2011\ : CascadeBuf
    port map (
            O => \N__10048\,
            I => \N__10042\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__10045\,
            I => \N__10039\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__10042\,
            I => \N__10036\
        );

    \I__2008\ : CascadeBuf
    port map (
            O => \N__10039\,
            I => \N__10033\
        );

    \I__2007\ : CascadeBuf
    port map (
            O => \N__10036\,
            I => \N__10030\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__10033\,
            I => \N__10027\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__10030\,
            I => \N__10024\
        );

    \I__2004\ : CascadeBuf
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__2003\ : CascadeBuf
    port map (
            O => \N__10024\,
            I => \N__10018\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__10021\,
            I => \N__10015\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__10018\,
            I => \N__10012\
        );

    \I__2000\ : CascadeBuf
    port map (
            O => \N__10015\,
            I => \N__10009\
        );

    \I__1999\ : CascadeBuf
    port map (
            O => \N__10012\,
            I => \N__10006\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__10009\,
            I => \N__10003\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__10006\,
            I => \N__10000\
        );

    \I__1996\ : InMux
    port map (
            O => \N__10003\,
            I => \N__9997\
        );

    \I__1995\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9994\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__9997\,
            I => \N__9991\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9994\,
            I => \N__9988\
        );

    \I__1992\ : Sp12to4
    port map (
            O => \N__9991\,
            I => \N__9985\
        );

    \I__1991\ : Span12Mux_v
    port map (
            O => \N__9988\,
            I => \N__9982\
        );

    \I__1990\ : Span12Mux_s3_v
    port map (
            O => \N__9985\,
            I => \N__9979\
        );

    \I__1989\ : Span12Mux_h
    port map (
            O => \N__9982\,
            I => \N__9976\
        );

    \I__1988\ : Span12Mux_v
    port map (
            O => \N__9979\,
            I => \N__9973\
        );

    \I__1987\ : Odrv12
    port map (
            O => \N__9976\,
            I => \M_this_vga_signals_address_5\
        );

    \I__1986\ : Odrv12
    port map (
            O => \N__9973\,
            I => \M_this_vga_signals_address_5\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__1984\ : CascadeBuf
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__9962\,
            I => \N__9959\
        );

    \I__1982\ : CascadeBuf
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__9956\,
            I => \N__9952\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__9955\,
            I => \N__9949\
        );

    \I__1979\ : CascadeBuf
    port map (
            O => \N__9952\,
            I => \N__9946\
        );

    \I__1978\ : CascadeBuf
    port map (
            O => \N__9949\,
            I => \N__9943\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__9946\,
            I => \N__9940\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__9943\,
            I => \N__9937\
        );

    \I__1975\ : CascadeBuf
    port map (
            O => \N__9940\,
            I => \N__9934\
        );

    \I__1974\ : CascadeBuf
    port map (
            O => \N__9937\,
            I => \N__9931\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__9934\,
            I => \N__9928\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__9931\,
            I => \N__9925\
        );

    \I__1971\ : CascadeBuf
    port map (
            O => \N__9928\,
            I => \N__9922\
        );

    \I__1970\ : CascadeBuf
    port map (
            O => \N__9925\,
            I => \N__9919\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__9922\,
            I => \N__9916\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__9919\,
            I => \N__9913\
        );

    \I__1967\ : CascadeBuf
    port map (
            O => \N__9916\,
            I => \N__9910\
        );

    \I__1966\ : CascadeBuf
    port map (
            O => \N__9913\,
            I => \N__9907\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__9910\,
            I => \N__9904\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__9907\,
            I => \N__9901\
        );

    \I__1963\ : CascadeBuf
    port map (
            O => \N__9904\,
            I => \N__9898\
        );

    \I__1962\ : CascadeBuf
    port map (
            O => \N__9901\,
            I => \N__9895\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__9898\,
            I => \N__9892\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__9895\,
            I => \N__9889\
        );

    \I__1959\ : CascadeBuf
    port map (
            O => \N__9892\,
            I => \N__9886\
        );

    \I__1958\ : CascadeBuf
    port map (
            O => \N__9889\,
            I => \N__9883\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__9886\,
            I => \N__9880\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__9883\,
            I => \N__9877\
        );

    \I__1955\ : CascadeBuf
    port map (
            O => \N__9880\,
            I => \N__9874\
        );

    \I__1954\ : CascadeBuf
    port map (
            O => \N__9877\,
            I => \N__9871\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__9874\,
            I => \N__9868\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__9871\,
            I => \N__9865\
        );

    \I__1951\ : CascadeBuf
    port map (
            O => \N__9868\,
            I => \N__9862\
        );

    \I__1950\ : CascadeBuf
    port map (
            O => \N__9865\,
            I => \N__9859\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__9862\,
            I => \N__9856\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__9859\,
            I => \N__9853\
        );

    \I__1947\ : CascadeBuf
    port map (
            O => \N__9856\,
            I => \N__9850\
        );

    \I__1946\ : CascadeBuf
    port map (
            O => \N__9853\,
            I => \N__9847\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__9850\,
            I => \N__9844\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__9847\,
            I => \N__9841\
        );

    \I__1943\ : CascadeBuf
    port map (
            O => \N__9844\,
            I => \N__9838\
        );

    \I__1942\ : CascadeBuf
    port map (
            O => \N__9841\,
            I => \N__9835\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__9838\,
            I => \N__9832\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__9835\,
            I => \N__9829\
        );

    \I__1939\ : CascadeBuf
    port map (
            O => \N__9832\,
            I => \N__9826\
        );

    \I__1938\ : CascadeBuf
    port map (
            O => \N__9829\,
            I => \N__9823\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__9826\,
            I => \N__9820\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__9823\,
            I => \N__9817\
        );

    \I__1935\ : CascadeBuf
    port map (
            O => \N__9820\,
            I => \N__9814\
        );

    \I__1934\ : CascadeBuf
    port map (
            O => \N__9817\,
            I => \N__9811\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__9814\,
            I => \N__9808\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__1931\ : CascadeBuf
    port map (
            O => \N__9808\,
            I => \N__9802\
        );

    \I__1930\ : CascadeBuf
    port map (
            O => \N__9805\,
            I => \N__9799\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__9802\,
            I => \N__9796\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__9799\,
            I => \N__9793\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9790\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9787\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9790\,
            I => \N__9784\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9787\,
            I => \N__9781\
        );

    \I__1923\ : Span4Mux_s2_v
    port map (
            O => \N__9784\,
            I => \N__9778\
        );

    \I__1922\ : Span12Mux_v
    port map (
            O => \N__9781\,
            I => \N__9775\
        );

    \I__1921\ : Sp12to4
    port map (
            O => \N__9778\,
            I => \N__9772\
        );

    \I__1920\ : Span12Mux_h
    port map (
            O => \N__9775\,
            I => \N__9769\
        );

    \I__1919\ : Span12Mux_v
    port map (
            O => \N__9772\,
            I => \N__9766\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__9769\,
            I => \M_this_vga_signals_address_6\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__9766\,
            I => \M_this_vga_signals_address_6\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9761\,
            I => \this_vga_signals.address_1_0_cry_0\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__9758\,
            I => \N__9755\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__9749\,
            I => \this_vga_signals.address_1\
        );

    \I__1911\ : InMux
    port map (
            O => \N__9746\,
            I => \this_vga_signals.address_1_0_cry_1\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__9743\,
            I => \N__9740\
        );

    \I__1909\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9737\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__9737\,
            I => \N__9734\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__9734\,
            I => \this_vga_signals.address_1_0_3\
        );

    \I__1906\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9725\
        );

    \I__1905\ : InMux
    port map (
            O => \N__9730\,
            I => \N__9725\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9725\,
            I => \this_vga_signals.m27_0_o2_1\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__9722\,
            I => \this_vga_signals.m27_0_0_cascade_\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__9719\,
            I => \this_vga_signals.i9_mux_cascade_\
        );

    \I__1901\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9710\
        );

    \I__1900\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9710\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__9710\,
            I => \this_vga_signals.N_40\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__1897\ : CascadeBuf
    port map (
            O => \N__9704\,
            I => \N__9701\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__9701\,
            I => \N__9698\
        );

    \I__1895\ : CascadeBuf
    port map (
            O => \N__9698\,
            I => \N__9695\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__9695\,
            I => \N__9691\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__9694\,
            I => \N__9688\
        );

    \I__1892\ : CascadeBuf
    port map (
            O => \N__9691\,
            I => \N__9685\
        );

    \I__1891\ : CascadeBuf
    port map (
            O => \N__9688\,
            I => \N__9682\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__9685\,
            I => \N__9679\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__9682\,
            I => \N__9676\
        );

    \I__1888\ : CascadeBuf
    port map (
            O => \N__9679\,
            I => \N__9673\
        );

    \I__1887\ : CascadeBuf
    port map (
            O => \N__9676\,
            I => \N__9670\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__9673\,
            I => \N__9667\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__9670\,
            I => \N__9664\
        );

    \I__1884\ : CascadeBuf
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__1883\ : CascadeBuf
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__9661\,
            I => \N__9655\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__9658\,
            I => \N__9652\
        );

    \I__1880\ : CascadeBuf
    port map (
            O => \N__9655\,
            I => \N__9649\
        );

    \I__1879\ : CascadeBuf
    port map (
            O => \N__9652\,
            I => \N__9646\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__9649\,
            I => \N__9643\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__9646\,
            I => \N__9640\
        );

    \I__1876\ : CascadeBuf
    port map (
            O => \N__9643\,
            I => \N__9637\
        );

    \I__1875\ : CascadeBuf
    port map (
            O => \N__9640\,
            I => \N__9634\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__9637\,
            I => \N__9631\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__9634\,
            I => \N__9628\
        );

    \I__1872\ : CascadeBuf
    port map (
            O => \N__9631\,
            I => \N__9625\
        );

    \I__1871\ : CascadeBuf
    port map (
            O => \N__9628\,
            I => \N__9622\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__9625\,
            I => \N__9619\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__9622\,
            I => \N__9616\
        );

    \I__1868\ : CascadeBuf
    port map (
            O => \N__9619\,
            I => \N__9613\
        );

    \I__1867\ : CascadeBuf
    port map (
            O => \N__9616\,
            I => \N__9610\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__9613\,
            I => \N__9607\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__9610\,
            I => \N__9604\
        );

    \I__1864\ : CascadeBuf
    port map (
            O => \N__9607\,
            I => \N__9601\
        );

    \I__1863\ : CascadeBuf
    port map (
            O => \N__9604\,
            I => \N__9598\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__9601\,
            I => \N__9595\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__9598\,
            I => \N__9592\
        );

    \I__1860\ : CascadeBuf
    port map (
            O => \N__9595\,
            I => \N__9589\
        );

    \I__1859\ : CascadeBuf
    port map (
            O => \N__9592\,
            I => \N__9586\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__9589\,
            I => \N__9583\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__9586\,
            I => \N__9580\
        );

    \I__1856\ : CascadeBuf
    port map (
            O => \N__9583\,
            I => \N__9577\
        );

    \I__1855\ : CascadeBuf
    port map (
            O => \N__9580\,
            I => \N__9574\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__9577\,
            I => \N__9571\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__9574\,
            I => \N__9568\
        );

    \I__1852\ : CascadeBuf
    port map (
            O => \N__9571\,
            I => \N__9565\
        );

    \I__1851\ : CascadeBuf
    port map (
            O => \N__9568\,
            I => \N__9562\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__9565\,
            I => \N__9559\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__9562\,
            I => \N__9556\
        );

    \I__1848\ : CascadeBuf
    port map (
            O => \N__9559\,
            I => \N__9553\
        );

    \I__1847\ : CascadeBuf
    port map (
            O => \N__9556\,
            I => \N__9550\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__9553\,
            I => \N__9547\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__9550\,
            I => \N__9544\
        );

    \I__1844\ : CascadeBuf
    port map (
            O => \N__9547\,
            I => \N__9541\
        );

    \I__1843\ : CascadeBuf
    port map (
            O => \N__9544\,
            I => \N__9538\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__9541\,
            I => \N__9535\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__9538\,
            I => \N__9532\
        );

    \I__1840\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9529\
        );

    \I__1839\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9526\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__9529\,
            I => \N__9523\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__9526\,
            I => \N__9520\
        );

    \I__1836\ : Sp12to4
    port map (
            O => \N__9523\,
            I => \N__9517\
        );

    \I__1835\ : Span12Mux_s9_v
    port map (
            O => \N__9520\,
            I => \N__9514\
        );

    \I__1834\ : Span12Mux_s5_v
    port map (
            O => \N__9517\,
            I => \N__9511\
        );

    \I__1833\ : Span12Mux_h
    port map (
            O => \N__9514\,
            I => \N__9508\
        );

    \I__1832\ : Span12Mux_v
    port map (
            O => \N__9511\,
            I => \N__9505\
        );

    \I__1831\ : Odrv12
    port map (
            O => \N__9508\,
            I => \M_this_vga_signals_address_7\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__9505\,
            I => \M_this_vga_signals_address_7\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__1828\ : CascadeBuf
    port map (
            O => \N__9497\,
            I => \N__9494\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__1826\ : CascadeBuf
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__9488\,
            I => \N__9484\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__9487\,
            I => \N__9481\
        );

    \I__1823\ : CascadeBuf
    port map (
            O => \N__9484\,
            I => \N__9478\
        );

    \I__1822\ : CascadeBuf
    port map (
            O => \N__9481\,
            I => \N__9475\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__9478\,
            I => \N__9472\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__9475\,
            I => \N__9469\
        );

    \I__1819\ : CascadeBuf
    port map (
            O => \N__9472\,
            I => \N__9466\
        );

    \I__1818\ : CascadeBuf
    port map (
            O => \N__9469\,
            I => \N__9463\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__9466\,
            I => \N__9460\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__9463\,
            I => \N__9457\
        );

    \I__1815\ : CascadeBuf
    port map (
            O => \N__9460\,
            I => \N__9454\
        );

    \I__1814\ : CascadeBuf
    port map (
            O => \N__9457\,
            I => \N__9451\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__9454\,
            I => \N__9448\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__9451\,
            I => \N__9445\
        );

    \I__1811\ : CascadeBuf
    port map (
            O => \N__9448\,
            I => \N__9442\
        );

    \I__1810\ : CascadeBuf
    port map (
            O => \N__9445\,
            I => \N__9439\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__9442\,
            I => \N__9436\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__9439\,
            I => \N__9433\
        );

    \I__1807\ : CascadeBuf
    port map (
            O => \N__9436\,
            I => \N__9430\
        );

    \I__1806\ : CascadeBuf
    port map (
            O => \N__9433\,
            I => \N__9427\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__9430\,
            I => \N__9424\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__9427\,
            I => \N__9421\
        );

    \I__1803\ : CascadeBuf
    port map (
            O => \N__9424\,
            I => \N__9418\
        );

    \I__1802\ : CascadeBuf
    port map (
            O => \N__9421\,
            I => \N__9415\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__9418\,
            I => \N__9412\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__9415\,
            I => \N__9409\
        );

    \I__1799\ : CascadeBuf
    port map (
            O => \N__9412\,
            I => \N__9406\
        );

    \I__1798\ : CascadeBuf
    port map (
            O => \N__9409\,
            I => \N__9403\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__9406\,
            I => \N__9400\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__9403\,
            I => \N__9397\
        );

    \I__1795\ : CascadeBuf
    port map (
            O => \N__9400\,
            I => \N__9394\
        );

    \I__1794\ : CascadeBuf
    port map (
            O => \N__9397\,
            I => \N__9391\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__9394\,
            I => \N__9388\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__9391\,
            I => \N__9385\
        );

    \I__1791\ : CascadeBuf
    port map (
            O => \N__9388\,
            I => \N__9382\
        );

    \I__1790\ : CascadeBuf
    port map (
            O => \N__9385\,
            I => \N__9379\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__9382\,
            I => \N__9376\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__9379\,
            I => \N__9373\
        );

    \I__1787\ : CascadeBuf
    port map (
            O => \N__9376\,
            I => \N__9370\
        );

    \I__1786\ : CascadeBuf
    port map (
            O => \N__9373\,
            I => \N__9367\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__9370\,
            I => \N__9364\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__9367\,
            I => \N__9361\
        );

    \I__1783\ : CascadeBuf
    port map (
            O => \N__9364\,
            I => \N__9358\
        );

    \I__1782\ : CascadeBuf
    port map (
            O => \N__9361\,
            I => \N__9355\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__9358\,
            I => \N__9352\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__9355\,
            I => \N__9349\
        );

    \I__1779\ : CascadeBuf
    port map (
            O => \N__9352\,
            I => \N__9346\
        );

    \I__1778\ : CascadeBuf
    port map (
            O => \N__9349\,
            I => \N__9343\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__9346\,
            I => \N__9340\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__9343\,
            I => \N__9337\
        );

    \I__1775\ : CascadeBuf
    port map (
            O => \N__9340\,
            I => \N__9334\
        );

    \I__1774\ : CascadeBuf
    port map (
            O => \N__9337\,
            I => \N__9331\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__9334\,
            I => \N__9328\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__9331\,
            I => \N__9325\
        );

    \I__1771\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9322\
        );

    \I__1770\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9319\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N__9316\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N__9313\
        );

    \I__1767\ : Sp12to4
    port map (
            O => \N__9316\,
            I => \N__9310\
        );

    \I__1766\ : Span12Mux_s8_v
    port map (
            O => \N__9313\,
            I => \N__9307\
        );

    \I__1765\ : Span12Mux_s5_v
    port map (
            O => \N__9310\,
            I => \N__9304\
        );

    \I__1764\ : Span12Mux_h
    port map (
            O => \N__9307\,
            I => \N__9301\
        );

    \I__1763\ : Span12Mux_v
    port map (
            O => \N__9304\,
            I => \N__9298\
        );

    \I__1762\ : Odrv12
    port map (
            O => \N__9301\,
            I => \M_this_vga_signals_address_8\
        );

    \I__1761\ : Odrv12
    port map (
            O => \N__9298\,
            I => \M_this_vga_signals_address_8\
        );

    \I__1760\ : InMux
    port map (
            O => \N__9293\,
            I => \this_vga_signals.address_1_cry_0\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__1758\ : CascadeBuf
    port map (
            O => \N__9287\,
            I => \N__9283\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__9286\,
            I => \N__9280\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__9283\,
            I => \N__9277\
        );

    \I__1755\ : CascadeBuf
    port map (
            O => \N__9280\,
            I => \N__9274\
        );

    \I__1754\ : CascadeBuf
    port map (
            O => \N__9277\,
            I => \N__9271\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__9274\,
            I => \N__9268\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__9271\,
            I => \N__9265\
        );

    \I__1751\ : CascadeBuf
    port map (
            O => \N__9268\,
            I => \N__9262\
        );

    \I__1750\ : CascadeBuf
    port map (
            O => \N__9265\,
            I => \N__9259\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__9262\,
            I => \N__9256\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__9259\,
            I => \N__9253\
        );

    \I__1747\ : CascadeBuf
    port map (
            O => \N__9256\,
            I => \N__9250\
        );

    \I__1746\ : CascadeBuf
    port map (
            O => \N__9253\,
            I => \N__9247\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__9250\,
            I => \N__9244\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__9247\,
            I => \N__9241\
        );

    \I__1743\ : CascadeBuf
    port map (
            O => \N__9244\,
            I => \N__9238\
        );

    \I__1742\ : CascadeBuf
    port map (
            O => \N__9241\,
            I => \N__9235\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__9238\,
            I => \N__9232\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__1739\ : CascadeBuf
    port map (
            O => \N__9232\,
            I => \N__9226\
        );

    \I__1738\ : CascadeBuf
    port map (
            O => \N__9229\,
            I => \N__9223\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N__9220\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__9223\,
            I => \N__9217\
        );

    \I__1735\ : CascadeBuf
    port map (
            O => \N__9220\,
            I => \N__9214\
        );

    \I__1734\ : CascadeBuf
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__9214\,
            I => \N__9208\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__9211\,
            I => \N__9205\
        );

    \I__1731\ : CascadeBuf
    port map (
            O => \N__9208\,
            I => \N__9202\
        );

    \I__1730\ : CascadeBuf
    port map (
            O => \N__9205\,
            I => \N__9199\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__9202\,
            I => \N__9196\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__9199\,
            I => \N__9193\
        );

    \I__1727\ : CascadeBuf
    port map (
            O => \N__9196\,
            I => \N__9190\
        );

    \I__1726\ : CascadeBuf
    port map (
            O => \N__9193\,
            I => \N__9187\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__9187\,
            I => \N__9181\
        );

    \I__1723\ : CascadeBuf
    port map (
            O => \N__9184\,
            I => \N__9178\
        );

    \I__1722\ : CascadeBuf
    port map (
            O => \N__9181\,
            I => \N__9175\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__9178\,
            I => \N__9172\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__9175\,
            I => \N__9169\
        );

    \I__1719\ : CascadeBuf
    port map (
            O => \N__9172\,
            I => \N__9166\
        );

    \I__1718\ : CascadeBuf
    port map (
            O => \N__9169\,
            I => \N__9163\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__9166\,
            I => \N__9160\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__1715\ : CascadeBuf
    port map (
            O => \N__9160\,
            I => \N__9154\
        );

    \I__1714\ : CascadeBuf
    port map (
            O => \N__9157\,
            I => \N__9151\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__9154\,
            I => \N__9148\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__9151\,
            I => \N__9145\
        );

    \I__1711\ : CascadeBuf
    port map (
            O => \N__9148\,
            I => \N__9142\
        );

    \I__1710\ : CascadeBuf
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__9139\,
            I => \N__9133\
        );

    \I__1707\ : CascadeBuf
    port map (
            O => \N__9136\,
            I => \N__9130\
        );

    \I__1706\ : CascadeBuf
    port map (
            O => \N__9133\,
            I => \N__9127\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__9130\,
            I => \N__9124\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__9127\,
            I => \N__9121\
        );

    \I__1703\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9118\
        );

    \I__1702\ : CascadeBuf
    port map (
            O => \N__9121\,
            I => \N__9115\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__9118\,
            I => \N__9112\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__9115\,
            I => \N__9109\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__9112\,
            I => \N__9106\
        );

    \I__1698\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9103\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__9106\,
            I => \N__9100\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__9103\,
            I => \N__9097\
        );

    \I__1695\ : Span4Mux_h
    port map (
            O => \N__9100\,
            I => \N__9094\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__9097\,
            I => \N__9091\
        );

    \I__1693\ : Span4Mux_h
    port map (
            O => \N__9094\,
            I => \N__9088\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__9091\,
            I => \N__9085\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__9088\,
            I => \N__9080\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__9085\,
            I => \N__9080\
        );

    \I__1689\ : Sp12to4
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__9077\,
            I => \M_this_vga_signals_address_9\
        );

    \I__1687\ : InMux
    port map (
            O => \N__9074\,
            I => \this_vga_signals.address_1_cry_1\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__1685\ : CascadeBuf
    port map (
            O => \N__9068\,
            I => \N__9064\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__9067\,
            I => \N__9061\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__9064\,
            I => \N__9058\
        );

    \I__1682\ : CascadeBuf
    port map (
            O => \N__9061\,
            I => \N__9055\
        );

    \I__1681\ : CascadeBuf
    port map (
            O => \N__9058\,
            I => \N__9052\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__9055\,
            I => \N__9049\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__9052\,
            I => \N__9046\
        );

    \I__1678\ : CascadeBuf
    port map (
            O => \N__9049\,
            I => \N__9043\
        );

    \I__1677\ : CascadeBuf
    port map (
            O => \N__9046\,
            I => \N__9040\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__9043\,
            I => \N__9037\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__9040\,
            I => \N__9034\
        );

    \I__1674\ : CascadeBuf
    port map (
            O => \N__9037\,
            I => \N__9031\
        );

    \I__1673\ : CascadeBuf
    port map (
            O => \N__9034\,
            I => \N__9028\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__9031\,
            I => \N__9025\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__9028\,
            I => \N__9022\
        );

    \I__1670\ : CascadeBuf
    port map (
            O => \N__9025\,
            I => \N__9019\
        );

    \I__1669\ : CascadeBuf
    port map (
            O => \N__9022\,
            I => \N__9016\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__9019\,
            I => \N__9013\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__9016\,
            I => \N__9010\
        );

    \I__1666\ : CascadeBuf
    port map (
            O => \N__9013\,
            I => \N__9007\
        );

    \I__1665\ : CascadeBuf
    port map (
            O => \N__9010\,
            I => \N__9004\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__9007\,
            I => \N__9001\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__9004\,
            I => \N__8998\
        );

    \I__1662\ : CascadeBuf
    port map (
            O => \N__9001\,
            I => \N__8995\
        );

    \I__1661\ : CascadeBuf
    port map (
            O => \N__8998\,
            I => \N__8992\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__8995\,
            I => \N__8989\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__8992\,
            I => \N__8986\
        );

    \I__1658\ : CascadeBuf
    port map (
            O => \N__8989\,
            I => \N__8983\
        );

    \I__1657\ : CascadeBuf
    port map (
            O => \N__8986\,
            I => \N__8980\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__8983\,
            I => \N__8977\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__8980\,
            I => \N__8974\
        );

    \I__1654\ : CascadeBuf
    port map (
            O => \N__8977\,
            I => \N__8971\
        );

    \I__1653\ : CascadeBuf
    port map (
            O => \N__8974\,
            I => \N__8968\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__8971\,
            I => \N__8965\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__8968\,
            I => \N__8962\
        );

    \I__1650\ : CascadeBuf
    port map (
            O => \N__8965\,
            I => \N__8959\
        );

    \I__1649\ : CascadeBuf
    port map (
            O => \N__8962\,
            I => \N__8956\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__8959\,
            I => \N__8953\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__8956\,
            I => \N__8950\
        );

    \I__1646\ : CascadeBuf
    port map (
            O => \N__8953\,
            I => \N__8947\
        );

    \I__1645\ : CascadeBuf
    port map (
            O => \N__8950\,
            I => \N__8944\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__8947\,
            I => \N__8941\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__8944\,
            I => \N__8938\
        );

    \I__1642\ : CascadeBuf
    port map (
            O => \N__8941\,
            I => \N__8935\
        );

    \I__1641\ : CascadeBuf
    port map (
            O => \N__8938\,
            I => \N__8932\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__8932\,
            I => \N__8926\
        );

    \I__1638\ : CascadeBuf
    port map (
            O => \N__8929\,
            I => \N__8923\
        );

    \I__1637\ : CascadeBuf
    port map (
            O => \N__8926\,
            I => \N__8920\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__8923\,
            I => \N__8917\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__8920\,
            I => \N__8914\
        );

    \I__1634\ : CascadeBuf
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__1633\ : CascadeBuf
    port map (
            O => \N__8914\,
            I => \N__8908\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__8911\,
            I => \N__8905\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__8908\,
            I => \N__8902\
        );

    \I__1630\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8899\
        );

    \I__1629\ : CascadeBuf
    port map (
            O => \N__8902\,
            I => \N__8896\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__8899\,
            I => \N__8893\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__8896\,
            I => \N__8890\
        );

    \I__1626\ : Span4Mux_v
    port map (
            O => \N__8893\,
            I => \N__8887\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8884\
        );

    \I__1624\ : Span4Mux_h
    port map (
            O => \N__8887\,
            I => \N__8881\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8884\,
            I => \N__8878\
        );

    \I__1622\ : Span4Mux_h
    port map (
            O => \N__8881\,
            I => \N__8875\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__8878\,
            I => \N__8872\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__8875\,
            I => \N__8869\
        );

    \I__1619\ : Span4Mux_h
    port map (
            O => \N__8872\,
            I => \N__8866\
        );

    \I__1618\ : Sp12to4
    port map (
            O => \N__8869\,
            I => \N__8861\
        );

    \I__1617\ : Sp12to4
    port map (
            O => \N__8866\,
            I => \N__8861\
        );

    \I__1616\ : Odrv12
    port map (
            O => \N__8861\,
            I => \M_this_vga_signals_address_10\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8858\,
            I => \this_vga_signals.address_1_cry_2\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8855\,
            I => \this_vga_signals.address_1_cry_3\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__1611\ : Span12Mux_s11_h
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1610\ : Span12Mux_v
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1609\ : Odrv12
    port map (
            O => \N__8840\,
            I => \this_vram.mem_out_bus4_2\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1606\ : Span4Mux_h
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1605\ : Sp12to4
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__1604\ : Span12Mux_v
    port map (
            O => \N__8825\,
            I => \N__8822\
        );

    \I__1603\ : Span12Mux_h
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__8819\,
            I => \this_vram.mem_out_bus6_2\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \this_vram.mem_mem_4_1_RNI14PZ0Z11_cascade_\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8810\,
            I => \this_vram.mem_N_2345\
        );

    \I__1598\ : CEMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__8804\,
            I => \N__8799\
        );

    \I__1596\ : CEMux
    port map (
            O => \N__8803\,
            I => \N__8796\
        );

    \I__1595\ : CEMux
    port map (
            O => \N__8802\,
            I => \N__8793\
        );

    \I__1594\ : Span4Mux_s3_v
    port map (
            O => \N__8799\,
            I => \N__8786\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__8796\,
            I => \N__8786\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__8793\,
            I => \N__8786\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__8780\,
            I => \this_vram.mem_WE_15\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__8777\,
            I => \this_vga_signals.m24_0_1_cascade_\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__8774\,
            I => \this_vga_signals.N_25_cascade_\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__8768\,
            I => \this_vga_signals.m24_0_1_0\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8762\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__8759\,
            I => \this_vram.mem_N_2327\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8753\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__8753\,
            I => \N__8750\
        );

    \I__1579\ : Span12Mux_v
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__1578\ : Odrv12
    port map (
            O => \N__8747\,
            I => \this_vram.mem_N_2353\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__8744\,
            I => \this_vram.mem_N_2355_cascade_\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__8741\,
            I => \N__8737\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__8740\,
            I => \N__8734\
        );

    \I__1574\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8727\
        );

    \I__1573\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8727\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8724\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8721\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8727\,
            I => \N__8716\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__8724\,
            I => \N__8716\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__8721\,
            I => \N__8713\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__8716\,
            I => \N__8707\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__8713\,
            I => \N__8707\
        );

    \I__1565\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8704\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__8707\,
            I => \this_vram.mem_G_25_0\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__8704\,
            I => \this_vram.mem_G_25_0\
        );

    \I__1562\ : IoInMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__8693\,
            I => \M_this_vram_read_data_1\
        );

    \I__1559\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8687\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1555\ : Odrv4
    port map (
            O => \N__8678\,
            I => \this_vram.mem_out_bus4_4\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1551\ : Sp12to4
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1550\ : Span12Mux_h
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__1549\ : Span12Mux_v
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__1548\ : Odrv12
    port map (
            O => \N__8657\,
            I => \this_vram.mem_out_bus6_4\
        );

    \I__1547\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__8651\,
            I => \this_vram.mem_mem_4_2_RNI34PZ0Z11\
        );

    \I__1545\ : CEMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__8645\,
            I => \N__8640\
        );

    \I__1543\ : CEMux
    port map (
            O => \N__8644\,
            I => \N__8637\
        );

    \I__1542\ : CEMux
    port map (
            O => \N__8643\,
            I => \N__8634\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__8640\,
            I => \N__8627\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8637\,
            I => \N__8627\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__8634\,
            I => \N__8627\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__8624\,
            I => \this_vram.mem_WE_18\
        );

    \I__1536\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__8618\,
            I => \N__8615\
        );

    \I__1534\ : Span4Mux_v
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1533\ : Sp12to4
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1532\ : Span12Mux_h
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1531\ : Span12Mux_v
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__8603\,
            I => \this_vram.mem_out_bus6_1\
        );

    \I__1529\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__8597\,
            I => \N__8594\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__8591\,
            I => \this_vram.mem_out_bus4_1\
        );

    \I__1525\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1521\ : Odrv4
    port map (
            O => \N__8576\,
            I => \this_vram.mem_out_bus5_1\
        );

    \I__1520\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__1518\ : Span4Mux_v
    port map (
            O => \N__8567\,
            I => \N__8564\
        );

    \I__1517\ : Sp12to4
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__1516\ : Span12Mux_h
    port map (
            O => \N__8561\,
            I => \N__8558\
        );

    \I__1515\ : Span12Mux_v
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1514\ : Odrv12
    port map (
            O => \N__8555\,
            I => \this_vram.mem_out_bus7_1\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8549\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__8549\,
            I => \this_vram.mem_mem_4_0_RNIV3P11Z0Z_0\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__8546\,
            I => \this_vram.mem_mem_5_0_RNI18R11Z0Z_0_cascade_\
        );

    \I__1510\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1508\ : Odrv12
    port map (
            O => \N__8537\,
            I => \this_vram.mem_N_2354\
        );

    \I__1507\ : CEMux
    port map (
            O => \N__8534\,
            I => \N__8530\
        );

    \I__1506\ : CEMux
    port map (
            O => \N__8533\,
            I => \N__8527\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__8530\,
            I => \N__8521\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__8527\,
            I => \N__8521\
        );

    \I__1503\ : CEMux
    port map (
            O => \N__8526\,
            I => \N__8518\
        );

    \I__1502\ : Span4Mux_v
    port map (
            O => \N__8521\,
            I => \N__8513\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8513\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__8510\,
            I => \this_vram.mem_WE_24\
        );

    \I__1498\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__8504\,
            I => \N__8501\
        );

    \I__1496\ : Odrv12
    port map (
            O => \N__8501\,
            I => \this_vram.mem_mem_0_0_RNILGF11Z0Z_0\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__8498\,
            I => \this_vram.mem_mem_2_0_RNIPOJ11Z0Z_0_cascade_\
        );

    \I__1494\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1492\ : Span4Mux_v
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1491\ : Sp12to4
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__1490\ : Span12Mux_h
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1489\ : Span12Mux_v
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__8477\,
            I => \this_vram.mem_out_bus6_0\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__1485\ : Span4Mux_v
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__8462\,
            I => \this_vram.mem_out_bus4_0\
        );

    \I__1482\ : CEMux
    port map (
            O => \N__8459\,
            I => \N__8455\
        );

    \I__1481\ : CEMux
    port map (
            O => \N__8458\,
            I => \N__8452\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__8455\,
            I => \N__8446\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__8452\,
            I => \N__8446\
        );

    \I__1478\ : CEMux
    port map (
            O => \N__8451\,
            I => \N__8443\
        );

    \I__1477\ : Span4Mux_v
    port map (
            O => \N__8446\,
            I => \N__8438\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__8443\,
            I => \N__8438\
        );

    \I__1475\ : Span4Mux_v
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__8432\,
            I => \this_vram.mem_WE_27\
        );

    \I__1472\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__8417\,
            I => \N__8414\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__8411\,
            I => \this_vram.mem_out_bus5_0\
        );

    \I__1465\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__8402\,
            I => \N__8399\
        );

    \I__1462\ : Sp12to4
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__1461\ : Span12Mux_h
    port map (
            O => \N__8396\,
            I => \N__8393\
        );

    \I__1460\ : Odrv12
    port map (
            O => \N__8393\,
            I => \this_vram.mem_out_bus7_0\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__8390\,
            I => \this_vram.mem_mem_5_0_RNI18RZ0Z11_cascade_\
        );

    \I__1458\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__8384\,
            I => \this_vram.mem_mem_4_0_RNIV3PZ0Z11\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8378\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__8375\,
            I => \N__8372\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__8372\,
            I => \this_vram.mem_N_2363\
        );

    \I__1452\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__8366\,
            I => \N__8363\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__8363\,
            I => \this_vram.mem_N_2344\
        );

    \I__1449\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8357\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__8357\,
            I => \this_vram.mem_N_2346\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__8354\,
            I => \this_vram.mem_G_25_0_cascade_\
        );

    \I__1446\ : IoInMux
    port map (
            O => \N__8351\,
            I => \N__8348\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__8348\,
            I => \N__8345\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__8345\,
            I => \M_this_vram_read_data_2\
        );

    \I__1443\ : CEMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8334\
        );

    \I__1441\ : CEMux
    port map (
            O => \N__8338\,
            I => \N__8331\
        );

    \I__1440\ : CEMux
    port map (
            O => \N__8337\,
            I => \N__8328\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__8334\,
            I => \N__8321\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__8331\,
            I => \N__8321\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__8328\,
            I => \N__8321\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__8321\,
            I => \this_vram.mem_WE_21\
        );

    \I__1435\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8315\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__8315\,
            I => \this_vram.mem_out_bus2_4\
        );

    \I__1433\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8309\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__8309\,
            I => \N__8306\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__8306\,
            I => \N__8303\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__8303\,
            I => \this_vram.mem_out_bus3_4\
        );

    \I__1429\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__1427\ : Span4Mux_v
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__8291\,
            I => \this_vram.mem_mem_0_2_RNIPGFZ0Z11\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__8288\,
            I => \this_vram.mem_mem_2_2_RNITOJZ0Z11_cascade_\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__8285\,
            I => \this_vram.mem_N_2326_cascade_\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__8282\,
            I => \N__8279\
        );

    \I__1422\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8276\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__8273\,
            I => \this_vram.mem_N_2373\
        );

    \I__1419\ : IoInMux
    port map (
            O => \N__8270\,
            I => \N__8267\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__8267\,
            I => \N__8264\
        );

    \I__1417\ : Span4Mux_s1_h
    port map (
            O => \N__8264\,
            I => \N__8261\
        );

    \I__1416\ : Sp12to4
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__1415\ : Span12Mux_v
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__8255\,
            I => \M_this_vram_read_data_5\
        );

    \I__1413\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8249\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__8249\,
            I => \N__8246\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__8246\,
            I => \this_vram.mem_N_2328\
        );

    \I__1410\ : IoInMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__1408\ : IoSpan4Mux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1407\ : Sp12to4
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__1406\ : Span12Mux_s6_h
    port map (
            O => \N__8231\,
            I => \N__8228\
        );

    \I__1405\ : Odrv12
    port map (
            O => \N__8228\,
            I => \M_this_vram_read_data_4\
        );

    \I__1404\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8222\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__1402\ : Odrv12
    port map (
            O => \N__8219\,
            I => \this_vram.mem_N_2337\
        );

    \I__1401\ : IoInMux
    port map (
            O => \N__8216\,
            I => \N__8213\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8210\
        );

    \I__1399\ : Span4Mux_s3_h
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__1398\ : Span4Mux_v
    port map (
            O => \N__8207\,
            I => \N__8204\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__8204\,
            I => \M_this_vram_read_data_3\
        );

    \I__1396\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8198\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1394\ : Span4Mux_v
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__8192\,
            I => \this_vram.mem_out_bus0_1\
        );

    \I__1392\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__8186\,
            I => \this_vram.mem_out_bus1_1\
        );

    \I__1390\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__8180\,
            I => \N__8177\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__8177\,
            I => \N__8174\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__8174\,
            I => \this_vram.mem_out_bus3_1\
        );

    \I__1386\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__8168\,
            I => \this_vram.mem_out_bus2_1\
        );

    \I__1384\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8162\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__8162\,
            I => \N__8159\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__8159\,
            I => \this_vram.mem_mem_0_1_RNINGF11Z0Z_0\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__8156\,
            I => \this_vram.mem_mem_2_1_RNIROJ11Z0Z_0_cascade_\
        );

    \I__1380\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8150\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__1378\ : Sp12to4
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__1377\ : Span12Mux_v
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__1376\ : Odrv12
    port map (
            O => \N__8141\,
            I => \this_vram.mem_out_bus4_3\
        );

    \I__1375\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8135\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__8135\,
            I => \N__8132\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__8132\,
            I => \N__8129\
        );

    \I__1372\ : Sp12to4
    port map (
            O => \N__8129\,
            I => \N__8126\
        );

    \I__1371\ : Span12Mux_h
    port map (
            O => \N__8126\,
            I => \N__8123\
        );

    \I__1370\ : Span12Mux_v
    port map (
            O => \N__8123\,
            I => \N__8120\
        );

    \I__1369\ : Odrv12
    port map (
            O => \N__8120\,
            I => \this_vram.mem_out_bus6_3\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__8117\,
            I => \this_vram.mem_mem_4_1_RNI14P11Z0Z_0_cascade_\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \this_vram.mem_N_2336_cascade_\
        );

    \I__1366\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__8108\,
            I => \this_vram.mem_N_2335\
        );

    \I__1364\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__8102\,
            I => \N__8099\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__8099\,
            I => \N__8096\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__8096\,
            I => \this_vram.mem_out_bus3_2\
        );

    \I__1360\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__8090\,
            I => \this_vram.mem_out_bus2_2\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__8087\,
            I => \this_vram.mem_mem_2_1_RNIROJZ0Z11_cascade_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__8075\,
            I => \this_vram.mem_mem_0_1_RNINGFZ0Z11\
        );

    \I__1353\ : InMux
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__1351\ : Span4Mux_v
    port map (
            O => \N__8066\,
            I => \N__8063\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__8063\,
            I => \this_vram.mem_out_bus3_5\
        );

    \I__1349\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8057\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__8057\,
            I => \this_vram.mem_out_bus2_5\
        );

    \I__1347\ : InMux
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1345\ : Span4Mux_v
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__8045\,
            I => \this_vram.mem_mem_0_2_RNIPGF11Z0Z_0\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__8042\,
            I => \this_vram.mem_mem_2_2_RNITOJ11Z0Z_0_cascade_\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__8039\,
            I => \this_vram.mem_N_2371_cascade_\
        );

    \I__1341\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__8033\,
            I => \N__8030\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__8030\,
            I => \N__8027\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__8027\,
            I => \this_vram.mem_out_bus0_3\
        );

    \I__1337\ : InMux
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__8021\,
            I => \this_vram.mem_out_bus1_3\
        );

    \I__1335\ : InMux
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__8009\,
            I => \this_vram.mem_out_bus0_4\
        );

    \I__1331\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__8003\,
            I => \this_vram.mem_out_bus1_4\
        );

    \I__1329\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7997\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7997\,
            I => \this_vram.mem_out_bus1_5\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7991\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__7985\,
            I => \this_vram.mem_out_bus0_5\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7979\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1321\ : Span4Mux_v
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1320\ : Odrv4
    port map (
            O => \N__7973\,
            I => \this_vram.mem_out_bus3_0\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7967\,
            I => \this_vram.mem_out_bus2_0\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1315\ : Odrv12
    port map (
            O => \N__7958\,
            I => \this_vram.mem_mem_0_0_RNILGFZ0Z11\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__7955\,
            I => \this_vram.mem_mem_2_0_RNIPOJZ0Z11_cascade_\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__7946\,
            I => \this_vram.mem_N_2362\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__7943\,
            I => \this_vram.mem_N_2364_cascade_\
        );

    \I__1309\ : IoInMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__1307\ : Span12Mux_s6_h
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1306\ : Odrv12
    port map (
            O => \N__7931\,
            I => \M_this_vram_read_data_0\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1303\ : Span4Mux_v
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__7919\,
            I => \this_vram.mem_out_bus3_3\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7913\,
            I => \this_vram.mem_out_bus2_3\
        );

    \I__1299\ : IoInMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1297\ : Span12Mux_s0_h
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__1296\ : Odrv12
    port map (
            O => \N__7901\,
            I => \this_vga_signals_N_170_i\
        );

    \I__1295\ : IoInMux
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__7895\,
            I => \this_vga_signals_N_171_i\
        );

    \I__1293\ : IoInMux
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7889\,
            I => \N__7884\
        );

    \I__1291\ : IoInMux
    port map (
            O => \N__7888\,
            I => \N__7881\
        );

    \I__1290\ : IoInMux
    port map (
            O => \N__7887\,
            I => \N__7878\
        );

    \I__1289\ : Span4Mux_s0_h
    port map (
            O => \N__7884\,
            I => \N__7874\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7869\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7878\,
            I => \N__7869\
        );

    \I__1286\ : IoInMux
    port map (
            O => \N__7877\,
            I => \N__7866\
        );

    \I__1285\ : Span4Mux_v
    port map (
            O => \N__7874\,
            I => \N__7863\
        );

    \I__1284\ : IoSpan4Mux
    port map (
            O => \N__7869\,
            I => \N__7858\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7866\,
            I => \N__7858\
        );

    \I__1282\ : Span4Mux_v
    port map (
            O => \N__7863\,
            I => \N__7855\
        );

    \I__1281\ : IoSpan4Mux
    port map (
            O => \N__7858\,
            I => \N__7852\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__7855\,
            I => \N__7847\
        );

    \I__1279\ : Span4Mux_s0_h
    port map (
            O => \N__7852\,
            I => \N__7847\
        );

    \I__1278\ : Span4Mux_v
    port map (
            O => \N__7847\,
            I => \N__7842\
        );

    \I__1277\ : IoInMux
    port map (
            O => \N__7846\,
            I => \N__7839\
        );

    \I__1276\ : IoInMux
    port map (
            O => \N__7845\,
            I => \N__7836\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__7842\,
            I => rgb5_i
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7839\,
            I => rgb5_i
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__7836\,
            I => rgb5_i
        );

    \I__1272\ : IoInMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7826\,
            I => vsync_c
        );

    \I__1270\ : IoInMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__1268\ : Span4Mux_s1_h
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__7814\,
            I => \N__7811\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__7811\,
            I => \this_vga_signals_N_94_i\
        );

    \I__1265\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__7799\,
            I => \this_vram.mem_out_bus0_0\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7793\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__7793\,
            I => \this_vram.mem_out_bus1_0\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7787\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__7787\,
            I => \N__7784\
        );

    \I__1257\ : Span4Mux_v
    port map (
            O => \N__7784\,
            I => \N__7781\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__7781\,
            I => \this_vram.mem_out_bus0_2\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7778\,
            I => \N__7775\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7775\,
            I => \this_vram.mem_out_bus1_2\
        );

    \I__1253\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7767\
        );

    \I__1252\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7762\
        );

    \I__1251\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7759\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__7767\,
            I => \N__7755\
        );

    \I__1249\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7752\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7765\,
            I => \N__7749\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__7762\,
            I => \N__7745\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__7759\,
            I => \N__7742\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7739\
        );

    \I__1244\ : Span12Mux_s9_h
    port map (
            O => \N__7755\,
            I => \N__7735\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__7752\,
            I => \N__7732\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7749\,
            I => \N__7729\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7726\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__7745\,
            I => \N__7723\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__7742\,
            I => \N__7720\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__7739\,
            I => \N__7717\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7738\,
            I => \N__7714\
        );

    \I__1236\ : Span12Mux_h
    port map (
            O => \N__7735\,
            I => \N__7709\
        );

    \I__1235\ : Span12Mux_s9_h
    port map (
            O => \N__7732\,
            I => \N__7706\
        );

    \I__1234\ : Span4Mux_h
    port map (
            O => \N__7729\,
            I => \N__7703\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7700\
        );

    \I__1232\ : Sp12to4
    port map (
            O => \N__7723\,
            I => \N__7697\
        );

    \I__1231\ : Span4Mux_h
    port map (
            O => \N__7720\,
            I => \N__7694\
        );

    \I__1230\ : Span12Mux_s10_h
    port map (
            O => \N__7717\,
            I => \N__7691\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7714\,
            I => \N__7688\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7685\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7682\
        );

    \I__1226\ : Span12Mux_v
    port map (
            O => \N__7709\,
            I => \N__7677\
        );

    \I__1225\ : Span12Mux_h
    port map (
            O => \N__7706\,
            I => \N__7677\
        );

    \I__1224\ : Sp12to4
    port map (
            O => \N__7703\,
            I => \N__7674\
        );

    \I__1223\ : Span4Mux_h
    port map (
            O => \N__7700\,
            I => \N__7671\
        );

    \I__1222\ : Span12Mux_v
    port map (
            O => \N__7697\,
            I => \N__7666\
        );

    \I__1221\ : Sp12to4
    port map (
            O => \N__7694\,
            I => \N__7666\
        );

    \I__1220\ : Span12Mux_v
    port map (
            O => \N__7691\,
            I => \N__7661\
        );

    \I__1219\ : Span12Mux_s10_h
    port map (
            O => \N__7688\,
            I => \N__7661\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7658\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__7682\,
            I => \N__7655\
        );

    \I__1216\ : Span12Mux_v
    port map (
            O => \N__7677\,
            I => \N__7652\
        );

    \I__1215\ : Span12Mux_v
    port map (
            O => \N__7674\,
            I => \N__7647\
        );

    \I__1214\ : Sp12to4
    port map (
            O => \N__7671\,
            I => \N__7647\
        );

    \I__1213\ : Span12Mux_h
    port map (
            O => \N__7666\,
            I => \N__7640\
        );

    \I__1212\ : Span12Mux_v
    port map (
            O => \N__7661\,
            I => \N__7640\
        );

    \I__1211\ : Span12Mux_s10_h
    port map (
            O => \N__7658\,
            I => \N__7640\
        );

    \I__1210\ : Span4Mux_h
    port map (
            O => \N__7655\,
            I => \N__7637\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__7652\,
            I => write_data_c_1
        );

    \I__1208\ : Odrv12
    port map (
            O => \N__7647\,
            I => write_data_c_1
        );

    \I__1207\ : Odrv12
    port map (
            O => \N__7640\,
            I => write_data_c_1
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__7637\,
            I => write_data_c_1
        );

    \I__1205\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__7625\,
            I => \N__7621\
        );

    \I__1203\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7618\
        );

    \I__1202\ : Span4Mux_h
    port map (
            O => \N__7621\,
            I => \N__7615\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__7618\,
            I => \N__7611\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__7615\,
            I => \N__7607\
        );

    \I__1199\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7604\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__7611\,
            I => \N__7601\
        );

    \I__1197\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7597\
        );

    \I__1196\ : Span4Mux_v
    port map (
            O => \N__7607\,
            I => \N__7594\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__7604\,
            I => \N__7591\
        );

    \I__1194\ : Span4Mux_v
    port map (
            O => \N__7601\,
            I => \N__7587\
        );

    \I__1193\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7584\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7581\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__7594\,
            I => \N__7575\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__7591\,
            I => \N__7575\
        );

    \I__1189\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7572\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__7587\,
            I => \N__7569\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__7584\,
            I => \N__7566\
        );

    \I__1186\ : Span4Mux_s2_v
    port map (
            O => \N__7581\,
            I => \N__7562\
        );

    \I__1185\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7559\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__7575\,
            I => \N__7556\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7572\,
            I => \N__7553\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__7569\,
            I => \N__7548\
        );

    \I__1181\ : Span4Mux_h
    port map (
            O => \N__7566\,
            I => \N__7548\
        );

    \I__1180\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7545\
        );

    \I__1179\ : Span4Mux_v
    port map (
            O => \N__7562\,
            I => \N__7540\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__7559\,
            I => \N__7540\
        );

    \I__1177\ : Span4Mux_h
    port map (
            O => \N__7556\,
            I => \N__7537\
        );

    \I__1176\ : Span4Mux_h
    port map (
            O => \N__7553\,
            I => \N__7534\
        );

    \I__1175\ : Span4Mux_h
    port map (
            O => \N__7548\,
            I => \N__7530\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__7545\,
            I => \N__7527\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__7540\,
            I => \N__7524\
        );

    \I__1172\ : Span4Mux_h
    port map (
            O => \N__7537\,
            I => \N__7519\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__7534\,
            I => \N__7519\
        );

    \I__1170\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7516\
        );

    \I__1169\ : Span4Mux_h
    port map (
            O => \N__7530\,
            I => \N__7513\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__7527\,
            I => \N__7510\
        );

    \I__1167\ : Sp12to4
    port map (
            O => \N__7524\,
            I => \N__7506\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__7519\,
            I => \N__7503\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__7516\,
            I => \N__7500\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__7513\,
            I => \N__7495\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__7510\,
            I => \N__7495\
        );

    \I__1162\ : InMux
    port map (
            O => \N__7509\,
            I => \N__7492\
        );

    \I__1161\ : Span12Mux_s10_h
    port map (
            O => \N__7506\,
            I => \N__7489\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__7503\,
            I => \N__7484\
        );

    \I__1159\ : Span4Mux_h
    port map (
            O => \N__7500\,
            I => \N__7484\
        );

    \I__1158\ : Span4Mux_v
    port map (
            O => \N__7495\,
            I => \N__7481\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__7492\,
            I => \N__7478\
        );

    \I__1156\ : Span12Mux_v
    port map (
            O => \N__7489\,
            I => \N__7475\
        );

    \I__1155\ : Span4Mux_v
    port map (
            O => \N__7484\,
            I => \N__7472\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__7481\,
            I => \N__7467\
        );

    \I__1153\ : Span4Mux_h
    port map (
            O => \N__7478\,
            I => \N__7467\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__7475\,
            I => write_data_c_0
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__7472\,
            I => write_data_c_0
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__7467\,
            I => write_data_c_0
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__7460\,
            I => \N__7457\
        );

    \I__1148\ : CascadeBuf
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1146\ : CascadeBuf
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__1144\ : CascadeBuf
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__7442\,
            I => \N__7438\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__7441\,
            I => \N__7435\
        );

    \I__1141\ : CascadeBuf
    port map (
            O => \N__7438\,
            I => \N__7432\
        );

    \I__1140\ : CascadeBuf
    port map (
            O => \N__7435\,
            I => \N__7429\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__7432\,
            I => \N__7426\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__7429\,
            I => \N__7423\
        );

    \I__1137\ : CascadeBuf
    port map (
            O => \N__7426\,
            I => \N__7420\
        );

    \I__1136\ : CascadeBuf
    port map (
            O => \N__7423\,
            I => \N__7417\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__7420\,
            I => \N__7414\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__7417\,
            I => \N__7411\
        );

    \I__1133\ : CascadeBuf
    port map (
            O => \N__7414\,
            I => \N__7408\
        );

    \I__1132\ : CascadeBuf
    port map (
            O => \N__7411\,
            I => \N__7405\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__7408\,
            I => \N__7402\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__7405\,
            I => \N__7399\
        );

    \I__1129\ : CascadeBuf
    port map (
            O => \N__7402\,
            I => \N__7396\
        );

    \I__1128\ : CascadeBuf
    port map (
            O => \N__7399\,
            I => \N__7393\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__7396\,
            I => \N__7390\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1125\ : CascadeBuf
    port map (
            O => \N__7390\,
            I => \N__7384\
        );

    \I__1124\ : CascadeBuf
    port map (
            O => \N__7387\,
            I => \N__7381\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__7384\,
            I => \N__7378\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__7381\,
            I => \N__7375\
        );

    \I__1121\ : CascadeBuf
    port map (
            O => \N__7378\,
            I => \N__7372\
        );

    \I__1120\ : CascadeBuf
    port map (
            O => \N__7375\,
            I => \N__7369\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__7372\,
            I => \N__7366\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__7369\,
            I => \N__7363\
        );

    \I__1117\ : CascadeBuf
    port map (
            O => \N__7366\,
            I => \N__7360\
        );

    \I__1116\ : CascadeBuf
    port map (
            O => \N__7363\,
            I => \N__7357\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__7360\,
            I => \N__7354\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__7357\,
            I => \N__7351\
        );

    \I__1113\ : CascadeBuf
    port map (
            O => \N__7354\,
            I => \N__7348\
        );

    \I__1112\ : CascadeBuf
    port map (
            O => \N__7351\,
            I => \N__7345\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__7348\,
            I => \N__7342\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__7345\,
            I => \N__7339\
        );

    \I__1109\ : CascadeBuf
    port map (
            O => \N__7342\,
            I => \N__7336\
        );

    \I__1108\ : CascadeBuf
    port map (
            O => \N__7339\,
            I => \N__7333\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__7336\,
            I => \N__7330\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__7333\,
            I => \N__7327\
        );

    \I__1105\ : CascadeBuf
    port map (
            O => \N__7330\,
            I => \N__7324\
        );

    \I__1104\ : CascadeBuf
    port map (
            O => \N__7327\,
            I => \N__7321\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__7324\,
            I => \N__7318\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__7321\,
            I => \N__7315\
        );

    \I__1101\ : CascadeBuf
    port map (
            O => \N__7318\,
            I => \N__7312\
        );

    \I__1100\ : CascadeBuf
    port map (
            O => \N__7315\,
            I => \N__7309\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__7312\,
            I => \N__7306\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__7309\,
            I => \N__7303\
        );

    \I__1097\ : CascadeBuf
    port map (
            O => \N__7306\,
            I => \N__7300\
        );

    \I__1096\ : CascadeBuf
    port map (
            O => \N__7303\,
            I => \N__7297\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__7300\,
            I => \N__7294\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__7297\,
            I => \N__7291\
        );

    \I__1093\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7288\
        );

    \I__1092\ : CascadeBuf
    port map (
            O => \N__7291\,
            I => \N__7285\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__7288\,
            I => \N__7282\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__7285\,
            I => \N__7279\
        );

    \I__1089\ : Span4Mux_s3_v
    port map (
            O => \N__7282\,
            I => \N__7276\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7273\
        );

    \I__1087\ : Span4Mux_h
    port map (
            O => \N__7276\,
            I => \N__7270\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__7273\,
            I => \N__7267\
        );

    \I__1085\ : Sp12to4
    port map (
            O => \N__7270\,
            I => \N__7264\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__7267\,
            I => \N__7261\
        );

    \I__1083\ : Span12Mux_h
    port map (
            O => \N__7264\,
            I => \N__7258\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__7261\,
            I => write_address_c_9
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__7258\,
            I => write_address_c_9
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__7253\,
            I => \N__7250\
        );

    \I__1079\ : CascadeBuf
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1077\ : CascadeBuf
    port map (
            O => \N__7244\,
            I => \N__7240\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__7243\,
            I => \N__7237\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__7240\,
            I => \N__7234\
        );

    \I__1074\ : CascadeBuf
    port map (
            O => \N__7237\,
            I => \N__7231\
        );

    \I__1073\ : CascadeBuf
    port map (
            O => \N__7234\,
            I => \N__7228\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__7231\,
            I => \N__7225\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__7228\,
            I => \N__7222\
        );

    \I__1070\ : CascadeBuf
    port map (
            O => \N__7225\,
            I => \N__7219\
        );

    \I__1069\ : CascadeBuf
    port map (
            O => \N__7222\,
            I => \N__7216\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__7219\,
            I => \N__7213\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__7216\,
            I => \N__7210\
        );

    \I__1066\ : CascadeBuf
    port map (
            O => \N__7213\,
            I => \N__7207\
        );

    \I__1065\ : CascadeBuf
    port map (
            O => \N__7210\,
            I => \N__7204\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__7207\,
            I => \N__7201\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__7204\,
            I => \N__7198\
        );

    \I__1062\ : CascadeBuf
    port map (
            O => \N__7201\,
            I => \N__7195\
        );

    \I__1061\ : CascadeBuf
    port map (
            O => \N__7198\,
            I => \N__7192\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__7195\,
            I => \N__7189\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__7192\,
            I => \N__7186\
        );

    \I__1058\ : CascadeBuf
    port map (
            O => \N__7189\,
            I => \N__7183\
        );

    \I__1057\ : CascadeBuf
    port map (
            O => \N__7186\,
            I => \N__7180\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__7183\,
            I => \N__7177\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__7180\,
            I => \N__7174\
        );

    \I__1054\ : CascadeBuf
    port map (
            O => \N__7177\,
            I => \N__7171\
        );

    \I__1053\ : CascadeBuf
    port map (
            O => \N__7174\,
            I => \N__7168\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__7171\,
            I => \N__7165\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__7168\,
            I => \N__7162\
        );

    \I__1050\ : CascadeBuf
    port map (
            O => \N__7165\,
            I => \N__7159\
        );

    \I__1049\ : CascadeBuf
    port map (
            O => \N__7162\,
            I => \N__7156\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__7159\,
            I => \N__7153\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__7156\,
            I => \N__7150\
        );

    \I__1046\ : CascadeBuf
    port map (
            O => \N__7153\,
            I => \N__7147\
        );

    \I__1045\ : CascadeBuf
    port map (
            O => \N__7150\,
            I => \N__7144\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \N__7141\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__7144\,
            I => \N__7138\
        );

    \I__1042\ : CascadeBuf
    port map (
            O => \N__7141\,
            I => \N__7135\
        );

    \I__1041\ : CascadeBuf
    port map (
            O => \N__7138\,
            I => \N__7132\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__7135\,
            I => \N__7129\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__7132\,
            I => \N__7126\
        );

    \I__1038\ : CascadeBuf
    port map (
            O => \N__7129\,
            I => \N__7123\
        );

    \I__1037\ : CascadeBuf
    port map (
            O => \N__7126\,
            I => \N__7120\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__7123\,
            I => \N__7117\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__7120\,
            I => \N__7114\
        );

    \I__1034\ : CascadeBuf
    port map (
            O => \N__7117\,
            I => \N__7111\
        );

    \I__1033\ : CascadeBuf
    port map (
            O => \N__7114\,
            I => \N__7108\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__7111\,
            I => \N__7105\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__7108\,
            I => \N__7102\
        );

    \I__1030\ : CascadeBuf
    port map (
            O => \N__7105\,
            I => \N__7099\
        );

    \I__1029\ : CascadeBuf
    port map (
            O => \N__7102\,
            I => \N__7096\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__7099\,
            I => \N__7093\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__7096\,
            I => \N__7090\
        );

    \I__1026\ : CascadeBuf
    port map (
            O => \N__7093\,
            I => \N__7087\
        );

    \I__1025\ : CascadeBuf
    port map (
            O => \N__7090\,
            I => \N__7084\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__7087\,
            I => \N__7081\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__7084\,
            I => \N__7078\
        );

    \I__1022\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7075\
        );

    \I__1021\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7072\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__7075\,
            I => \N__7069\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__7072\,
            I => \N__7066\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__7069\,
            I => \N__7063\
        );

    \I__1017\ : IoSpan4Mux
    port map (
            O => \N__7066\,
            I => \N__7060\
        );

    \I__1016\ : IoSpan4Mux
    port map (
            O => \N__7063\,
            I => \N__7057\
        );

    \I__1015\ : IoSpan4Mux
    port map (
            O => \N__7060\,
            I => \N__7054\
        );

    \I__1014\ : IoSpan4Mux
    port map (
            O => \N__7057\,
            I => \N__7051\
        );

    \I__1013\ : IoSpan4Mux
    port map (
            O => \N__7054\,
            I => \N__7048\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__7051\,
            I => write_address_c_8
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__7048\,
            I => write_address_c_8
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__1009\ : CascadeBuf
    port map (
            O => \N__7040\,
            I => \N__7037\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__1007\ : CascadeBuf
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__7031\,
            I => \N__7027\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__7030\,
            I => \N__7024\
        );

    \I__1004\ : CascadeBuf
    port map (
            O => \N__7027\,
            I => \N__7021\
        );

    \I__1003\ : CascadeBuf
    port map (
            O => \N__7024\,
            I => \N__7018\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__7021\,
            I => \N__7015\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__7018\,
            I => \N__7012\
        );

    \I__1000\ : CascadeBuf
    port map (
            O => \N__7015\,
            I => \N__7009\
        );

    \I__999\ : CascadeBuf
    port map (
            O => \N__7012\,
            I => \N__7006\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__7009\,
            I => \N__7003\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__7006\,
            I => \N__7000\
        );

    \I__996\ : CascadeBuf
    port map (
            O => \N__7003\,
            I => \N__6997\
        );

    \I__995\ : CascadeBuf
    port map (
            O => \N__7000\,
            I => \N__6994\
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__6997\,
            I => \N__6991\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__6994\,
            I => \N__6988\
        );

    \I__992\ : CascadeBuf
    port map (
            O => \N__6991\,
            I => \N__6985\
        );

    \I__991\ : CascadeBuf
    port map (
            O => \N__6988\,
            I => \N__6982\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__6985\,
            I => \N__6979\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__6982\,
            I => \N__6976\
        );

    \I__988\ : CascadeBuf
    port map (
            O => \N__6979\,
            I => \N__6973\
        );

    \I__987\ : CascadeBuf
    port map (
            O => \N__6976\,
            I => \N__6970\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__6973\,
            I => \N__6967\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__6970\,
            I => \N__6964\
        );

    \I__984\ : CascadeBuf
    port map (
            O => \N__6967\,
            I => \N__6961\
        );

    \I__983\ : CascadeBuf
    port map (
            O => \N__6964\,
            I => \N__6958\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__6961\,
            I => \N__6955\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__6958\,
            I => \N__6952\
        );

    \I__980\ : CascadeBuf
    port map (
            O => \N__6955\,
            I => \N__6949\
        );

    \I__979\ : CascadeBuf
    port map (
            O => \N__6952\,
            I => \N__6946\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__6949\,
            I => \N__6943\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__6946\,
            I => \N__6940\
        );

    \I__976\ : CascadeBuf
    port map (
            O => \N__6943\,
            I => \N__6937\
        );

    \I__975\ : CascadeBuf
    port map (
            O => \N__6940\,
            I => \N__6934\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__6937\,
            I => \N__6931\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__6934\,
            I => \N__6928\
        );

    \I__972\ : CascadeBuf
    port map (
            O => \N__6931\,
            I => \N__6925\
        );

    \I__971\ : CascadeBuf
    port map (
            O => \N__6928\,
            I => \N__6922\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__6925\,
            I => \N__6919\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__6922\,
            I => \N__6916\
        );

    \I__968\ : CascadeBuf
    port map (
            O => \N__6919\,
            I => \N__6913\
        );

    \I__967\ : CascadeBuf
    port map (
            O => \N__6916\,
            I => \N__6910\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__6913\,
            I => \N__6907\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__6910\,
            I => \N__6904\
        );

    \I__964\ : CascadeBuf
    port map (
            O => \N__6907\,
            I => \N__6901\
        );

    \I__963\ : CascadeBuf
    port map (
            O => \N__6904\,
            I => \N__6898\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__6901\,
            I => \N__6895\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6898\,
            I => \N__6892\
        );

    \I__960\ : CascadeBuf
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__959\ : CascadeBuf
    port map (
            O => \N__6892\,
            I => \N__6886\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__6889\,
            I => \N__6883\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__6886\,
            I => \N__6880\
        );

    \I__956\ : CascadeBuf
    port map (
            O => \N__6883\,
            I => \N__6877\
        );

    \I__955\ : CascadeBuf
    port map (
            O => \N__6880\,
            I => \N__6874\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__6877\,
            I => \N__6871\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__6874\,
            I => \N__6868\
        );

    \I__952\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6865\
        );

    \I__951\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6862\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6859\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6862\,
            I => \N__6856\
        );

    \I__948\ : Span4Mux_s2_v
    port map (
            O => \N__6859\,
            I => \N__6853\
        );

    \I__947\ : Span4Mux_h
    port map (
            O => \N__6856\,
            I => \N__6850\
        );

    \I__946\ : Sp12to4
    port map (
            O => \N__6853\,
            I => \N__6847\
        );

    \I__945\ : Sp12to4
    port map (
            O => \N__6850\,
            I => \N__6842\
        );

    \I__944\ : Span12Mux_h
    port map (
            O => \N__6847\,
            I => \N__6842\
        );

    \I__943\ : Span12Mux_v
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__942\ : Span12Mux_v
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__941\ : Odrv12
    port map (
            O => \N__6836\,
            I => write_address_c_7
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__6833\,
            I => \N__6830\
        );

    \I__939\ : CascadeBuf
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__937\ : CascadeBuf
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__6821\,
            I => \N__6818\
        );

    \I__935\ : CascadeBuf
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__6815\,
            I => \N__6811\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__6814\,
            I => \N__6808\
        );

    \I__932\ : CascadeBuf
    port map (
            O => \N__6811\,
            I => \N__6805\
        );

    \I__931\ : CascadeBuf
    port map (
            O => \N__6808\,
            I => \N__6802\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__6805\,
            I => \N__6799\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__6802\,
            I => \N__6796\
        );

    \I__928\ : CascadeBuf
    port map (
            O => \N__6799\,
            I => \N__6793\
        );

    \I__927\ : CascadeBuf
    port map (
            O => \N__6796\,
            I => \N__6790\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__6793\,
            I => \N__6787\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__6790\,
            I => \N__6784\
        );

    \I__924\ : CascadeBuf
    port map (
            O => \N__6787\,
            I => \N__6781\
        );

    \I__923\ : CascadeBuf
    port map (
            O => \N__6784\,
            I => \N__6778\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__6781\,
            I => \N__6775\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__6778\,
            I => \N__6772\
        );

    \I__920\ : CascadeBuf
    port map (
            O => \N__6775\,
            I => \N__6769\
        );

    \I__919\ : CascadeBuf
    port map (
            O => \N__6772\,
            I => \N__6766\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__6769\,
            I => \N__6763\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__6766\,
            I => \N__6760\
        );

    \I__916\ : CascadeBuf
    port map (
            O => \N__6763\,
            I => \N__6757\
        );

    \I__915\ : CascadeBuf
    port map (
            O => \N__6760\,
            I => \N__6754\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__6757\,
            I => \N__6751\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__6754\,
            I => \N__6748\
        );

    \I__912\ : CascadeBuf
    port map (
            O => \N__6751\,
            I => \N__6745\
        );

    \I__911\ : CascadeBuf
    port map (
            O => \N__6748\,
            I => \N__6742\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__6745\,
            I => \N__6739\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__6742\,
            I => \N__6736\
        );

    \I__908\ : CascadeBuf
    port map (
            O => \N__6739\,
            I => \N__6733\
        );

    \I__907\ : CascadeBuf
    port map (
            O => \N__6736\,
            I => \N__6730\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__6733\,
            I => \N__6727\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__6730\,
            I => \N__6724\
        );

    \I__904\ : CascadeBuf
    port map (
            O => \N__6727\,
            I => \N__6721\
        );

    \I__903\ : CascadeBuf
    port map (
            O => \N__6724\,
            I => \N__6718\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__6721\,
            I => \N__6715\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__6718\,
            I => \N__6712\
        );

    \I__900\ : CascadeBuf
    port map (
            O => \N__6715\,
            I => \N__6709\
        );

    \I__899\ : CascadeBuf
    port map (
            O => \N__6712\,
            I => \N__6706\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__6709\,
            I => \N__6703\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__6706\,
            I => \N__6700\
        );

    \I__896\ : CascadeBuf
    port map (
            O => \N__6703\,
            I => \N__6697\
        );

    \I__895\ : CascadeBuf
    port map (
            O => \N__6700\,
            I => \N__6694\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__6697\,
            I => \N__6691\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__6694\,
            I => \N__6688\
        );

    \I__892\ : CascadeBuf
    port map (
            O => \N__6691\,
            I => \N__6685\
        );

    \I__891\ : CascadeBuf
    port map (
            O => \N__6688\,
            I => \N__6682\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__6685\,
            I => \N__6679\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__6682\,
            I => \N__6676\
        );

    \I__888\ : CascadeBuf
    port map (
            O => \N__6679\,
            I => \N__6673\
        );

    \I__887\ : CascadeBuf
    port map (
            O => \N__6676\,
            I => \N__6670\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__6673\,
            I => \N__6667\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__6670\,
            I => \N__6664\
        );

    \I__884\ : InMux
    port map (
            O => \N__6667\,
            I => \N__6661\
        );

    \I__883\ : CascadeBuf
    port map (
            O => \N__6664\,
            I => \N__6658\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__6661\,
            I => \N__6655\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__6658\,
            I => \N__6652\
        );

    \I__880\ : Span4Mux_v
    port map (
            O => \N__6655\,
            I => \N__6649\
        );

    \I__879\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6646\
        );

    \I__878\ : Sp12to4
    port map (
            O => \N__6649\,
            I => \N__6643\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__6646\,
            I => \N__6640\
        );

    \I__876\ : Span12Mux_h
    port map (
            O => \N__6643\,
            I => \N__6637\
        );

    \I__875\ : Span12Mux_h
    port map (
            O => \N__6640\,
            I => \N__6634\
        );

    \I__874\ : Span12Mux_v
    port map (
            O => \N__6637\,
            I => \N__6631\
        );

    \I__873\ : Span12Mux_v
    port map (
            O => \N__6634\,
            I => \N__6626\
        );

    \I__872\ : Span12Mux_h
    port map (
            O => \N__6631\,
            I => \N__6626\
        );

    \I__871\ : Odrv12
    port map (
            O => \N__6626\,
            I => write_address_c_6
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__6623\,
            I => \N__6620\
        );

    \I__869\ : CascadeBuf
    port map (
            O => \N__6620\,
            I => \N__6617\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__6617\,
            I => \N__6614\
        );

    \I__867\ : CascadeBuf
    port map (
            O => \N__6614\,
            I => \N__6611\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__6611\,
            I => \N__6608\
        );

    \I__865\ : CascadeBuf
    port map (
            O => \N__6608\,
            I => \N__6605\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__6605\,
            I => \N__6601\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__6604\,
            I => \N__6598\
        );

    \I__862\ : CascadeBuf
    port map (
            O => \N__6601\,
            I => \N__6595\
        );

    \I__861\ : CascadeBuf
    port map (
            O => \N__6598\,
            I => \N__6592\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__6595\,
            I => \N__6589\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__6592\,
            I => \N__6586\
        );

    \I__858\ : CascadeBuf
    port map (
            O => \N__6589\,
            I => \N__6583\
        );

    \I__857\ : CascadeBuf
    port map (
            O => \N__6586\,
            I => \N__6580\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__6583\,
            I => \N__6577\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__6580\,
            I => \N__6574\
        );

    \I__854\ : CascadeBuf
    port map (
            O => \N__6577\,
            I => \N__6571\
        );

    \I__853\ : CascadeBuf
    port map (
            O => \N__6574\,
            I => \N__6568\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__6571\,
            I => \N__6565\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__6568\,
            I => \N__6562\
        );

    \I__850\ : CascadeBuf
    port map (
            O => \N__6565\,
            I => \N__6559\
        );

    \I__849\ : CascadeBuf
    port map (
            O => \N__6562\,
            I => \N__6556\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__846\ : CascadeBuf
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__845\ : CascadeBuf
    port map (
            O => \N__6550\,
            I => \N__6544\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__6547\,
            I => \N__6541\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__6544\,
            I => \N__6538\
        );

    \I__842\ : CascadeBuf
    port map (
            O => \N__6541\,
            I => \N__6535\
        );

    \I__841\ : CascadeBuf
    port map (
            O => \N__6538\,
            I => \N__6532\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__6535\,
            I => \N__6529\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__6532\,
            I => \N__6526\
        );

    \I__838\ : CascadeBuf
    port map (
            O => \N__6529\,
            I => \N__6523\
        );

    \I__837\ : CascadeBuf
    port map (
            O => \N__6526\,
            I => \N__6520\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__6523\,
            I => \N__6517\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__6520\,
            I => \N__6514\
        );

    \I__834\ : CascadeBuf
    port map (
            O => \N__6517\,
            I => \N__6511\
        );

    \I__833\ : CascadeBuf
    port map (
            O => \N__6514\,
            I => \N__6508\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__6511\,
            I => \N__6505\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__830\ : CascadeBuf
    port map (
            O => \N__6505\,
            I => \N__6499\
        );

    \I__829\ : CascadeBuf
    port map (
            O => \N__6502\,
            I => \N__6496\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__6499\,
            I => \N__6493\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__6496\,
            I => \N__6490\
        );

    \I__826\ : CascadeBuf
    port map (
            O => \N__6493\,
            I => \N__6487\
        );

    \I__825\ : CascadeBuf
    port map (
            O => \N__6490\,
            I => \N__6484\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__6487\,
            I => \N__6481\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__6484\,
            I => \N__6478\
        );

    \I__822\ : CascadeBuf
    port map (
            O => \N__6481\,
            I => \N__6475\
        );

    \I__821\ : CascadeBuf
    port map (
            O => \N__6478\,
            I => \N__6472\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__6475\,
            I => \N__6469\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__6472\,
            I => \N__6466\
        );

    \I__818\ : CascadeBuf
    port map (
            O => \N__6469\,
            I => \N__6463\
        );

    \I__817\ : CascadeBuf
    port map (
            O => \N__6466\,
            I => \N__6460\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__6463\,
            I => \N__6457\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__6460\,
            I => \N__6454\
        );

    \I__814\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6451\
        );

    \I__813\ : CascadeBuf
    port map (
            O => \N__6454\,
            I => \N__6448\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__6451\,
            I => \N__6445\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__6448\,
            I => \N__6442\
        );

    \I__810\ : Span4Mux_s3_v
    port map (
            O => \N__6445\,
            I => \N__6439\
        );

    \I__809\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6436\
        );

    \I__808\ : Span4Mux_v
    port map (
            O => \N__6439\,
            I => \N__6433\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__806\ : Span4Mux_v
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__805\ : Sp12to4
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__804\ : Sp12to4
    port map (
            O => \N__6427\,
            I => \N__6421\
        );

    \I__803\ : Span12Mux_s11_v
    port map (
            O => \N__6424\,
            I => \N__6418\
        );

    \I__802\ : Span12Mux_h
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__801\ : Odrv12
    port map (
            O => \N__6418\,
            I => write_address_c_5
        );

    \I__800\ : Odrv12
    port map (
            O => \N__6415\,
            I => write_address_c_5
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__798\ : CascadeBuf
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__796\ : CascadeBuf
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__794\ : CascadeBuf
    port map (
            O => \N__6395\,
            I => \N__6391\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__6394\,
            I => \N__6388\
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__6391\,
            I => \N__6385\
        );

    \I__791\ : CascadeBuf
    port map (
            O => \N__6388\,
            I => \N__6382\
        );

    \I__790\ : CascadeBuf
    port map (
            O => \N__6385\,
            I => \N__6379\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__6382\,
            I => \N__6376\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__6379\,
            I => \N__6373\
        );

    \I__787\ : CascadeBuf
    port map (
            O => \N__6376\,
            I => \N__6370\
        );

    \I__786\ : CascadeBuf
    port map (
            O => \N__6373\,
            I => \N__6367\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__6370\,
            I => \N__6364\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__783\ : CascadeBuf
    port map (
            O => \N__6364\,
            I => \N__6358\
        );

    \I__782\ : CascadeBuf
    port map (
            O => \N__6361\,
            I => \N__6355\
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__6358\,
            I => \N__6352\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__6355\,
            I => \N__6349\
        );

    \I__779\ : CascadeBuf
    port map (
            O => \N__6352\,
            I => \N__6346\
        );

    \I__778\ : CascadeBuf
    port map (
            O => \N__6349\,
            I => \N__6343\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__6346\,
            I => \N__6340\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__6343\,
            I => \N__6337\
        );

    \I__775\ : CascadeBuf
    port map (
            O => \N__6340\,
            I => \N__6334\
        );

    \I__774\ : CascadeBuf
    port map (
            O => \N__6337\,
            I => \N__6331\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__6334\,
            I => \N__6328\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__6331\,
            I => \N__6325\
        );

    \I__771\ : CascadeBuf
    port map (
            O => \N__6328\,
            I => \N__6322\
        );

    \I__770\ : CascadeBuf
    port map (
            O => \N__6325\,
            I => \N__6319\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__6322\,
            I => \N__6316\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__6319\,
            I => \N__6313\
        );

    \I__767\ : CascadeBuf
    port map (
            O => \N__6316\,
            I => \N__6310\
        );

    \I__766\ : CascadeBuf
    port map (
            O => \N__6313\,
            I => \N__6307\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__6310\,
            I => \N__6304\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__6307\,
            I => \N__6301\
        );

    \I__763\ : CascadeBuf
    port map (
            O => \N__6304\,
            I => \N__6298\
        );

    \I__762\ : CascadeBuf
    port map (
            O => \N__6301\,
            I => \N__6295\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__6298\,
            I => \N__6292\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__6295\,
            I => \N__6289\
        );

    \I__759\ : CascadeBuf
    port map (
            O => \N__6292\,
            I => \N__6286\
        );

    \I__758\ : CascadeBuf
    port map (
            O => \N__6289\,
            I => \N__6283\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__6286\,
            I => \N__6280\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__6283\,
            I => \N__6277\
        );

    \I__755\ : CascadeBuf
    port map (
            O => \N__6280\,
            I => \N__6274\
        );

    \I__754\ : CascadeBuf
    port map (
            O => \N__6277\,
            I => \N__6271\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__6274\,
            I => \N__6268\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__6271\,
            I => \N__6265\
        );

    \I__751\ : CascadeBuf
    port map (
            O => \N__6268\,
            I => \N__6262\
        );

    \I__750\ : CascadeBuf
    port map (
            O => \N__6265\,
            I => \N__6259\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__6262\,
            I => \N__6256\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__6259\,
            I => \N__6253\
        );

    \I__747\ : CascadeBuf
    port map (
            O => \N__6256\,
            I => \N__6250\
        );

    \I__746\ : CascadeBuf
    port map (
            O => \N__6253\,
            I => \N__6247\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__6250\,
            I => \N__6244\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__6247\,
            I => \N__6241\
        );

    \I__743\ : CascadeBuf
    port map (
            O => \N__6244\,
            I => \N__6238\
        );

    \I__742\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6235\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__6238\,
            I => \N__6232\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6229\
        );

    \I__739\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6226\
        );

    \I__738\ : Span4Mux_v
    port map (
            O => \N__6229\,
            I => \N__6223\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__6226\,
            I => \N__6220\
        );

    \I__736\ : Span4Mux_v
    port map (
            O => \N__6223\,
            I => \N__6217\
        );

    \I__735\ : Span4Mux_v
    port map (
            O => \N__6220\,
            I => \N__6214\
        );

    \I__734\ : Sp12to4
    port map (
            O => \N__6217\,
            I => \N__6211\
        );

    \I__733\ : Sp12to4
    port map (
            O => \N__6214\,
            I => \N__6206\
        );

    \I__732\ : Span12Mux_h
    port map (
            O => \N__6211\,
            I => \N__6206\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__6206\,
            I => write_address_c_4
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__729\ : CascadeBuf
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__6197\,
            I => \N__6194\
        );

    \I__727\ : CascadeBuf
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__6191\,
            I => \N__6188\
        );

    \I__725\ : CascadeBuf
    port map (
            O => \N__6188\,
            I => \N__6184\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__6187\,
            I => \N__6181\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__6184\,
            I => \N__6178\
        );

    \I__722\ : CascadeBuf
    port map (
            O => \N__6181\,
            I => \N__6175\
        );

    \I__721\ : CascadeBuf
    port map (
            O => \N__6178\,
            I => \N__6172\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__6175\,
            I => \N__6169\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__6172\,
            I => \N__6166\
        );

    \I__718\ : CascadeBuf
    port map (
            O => \N__6169\,
            I => \N__6163\
        );

    \I__717\ : CascadeBuf
    port map (
            O => \N__6166\,
            I => \N__6160\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__6163\,
            I => \N__6157\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__6160\,
            I => \N__6154\
        );

    \I__714\ : CascadeBuf
    port map (
            O => \N__6157\,
            I => \N__6151\
        );

    \I__713\ : CascadeBuf
    port map (
            O => \N__6154\,
            I => \N__6148\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__6151\,
            I => \N__6145\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__6148\,
            I => \N__6142\
        );

    \I__710\ : CascadeBuf
    port map (
            O => \N__6145\,
            I => \N__6139\
        );

    \I__709\ : CascadeBuf
    port map (
            O => \N__6142\,
            I => \N__6136\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__6139\,
            I => \N__6133\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__6136\,
            I => \N__6130\
        );

    \I__706\ : CascadeBuf
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__705\ : CascadeBuf
    port map (
            O => \N__6130\,
            I => \N__6124\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__6127\,
            I => \N__6121\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__6124\,
            I => \N__6118\
        );

    \I__702\ : CascadeBuf
    port map (
            O => \N__6121\,
            I => \N__6115\
        );

    \I__701\ : CascadeBuf
    port map (
            O => \N__6118\,
            I => \N__6112\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__6115\,
            I => \N__6109\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__6112\,
            I => \N__6106\
        );

    \I__698\ : CascadeBuf
    port map (
            O => \N__6109\,
            I => \N__6103\
        );

    \I__697\ : CascadeBuf
    port map (
            O => \N__6106\,
            I => \N__6100\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__6103\,
            I => \N__6097\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__6100\,
            I => \N__6094\
        );

    \I__694\ : CascadeBuf
    port map (
            O => \N__6097\,
            I => \N__6091\
        );

    \I__693\ : CascadeBuf
    port map (
            O => \N__6094\,
            I => \N__6088\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__6091\,
            I => \N__6085\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__6088\,
            I => \N__6082\
        );

    \I__690\ : CascadeBuf
    port map (
            O => \N__6085\,
            I => \N__6079\
        );

    \I__689\ : CascadeBuf
    port map (
            O => \N__6082\,
            I => \N__6076\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__6079\,
            I => \N__6073\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__6076\,
            I => \N__6070\
        );

    \I__686\ : CascadeBuf
    port map (
            O => \N__6073\,
            I => \N__6067\
        );

    \I__685\ : CascadeBuf
    port map (
            O => \N__6070\,
            I => \N__6064\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__6067\,
            I => \N__6061\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__6064\,
            I => \N__6058\
        );

    \I__682\ : CascadeBuf
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__681\ : CascadeBuf
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__6055\,
            I => \N__6049\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__6052\,
            I => \N__6046\
        );

    \I__678\ : CascadeBuf
    port map (
            O => \N__6049\,
            I => \N__6043\
        );

    \I__677\ : CascadeBuf
    port map (
            O => \N__6046\,
            I => \N__6040\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__6043\,
            I => \N__6037\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__6040\,
            I => \N__6034\
        );

    \I__674\ : CascadeBuf
    port map (
            O => \N__6037\,
            I => \N__6031\
        );

    \I__673\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6028\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__6028\,
            I => \N__6022\
        );

    \I__670\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6019\
        );

    \I__669\ : Span4Mux_s1_v
    port map (
            O => \N__6022\,
            I => \N__6016\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__6019\,
            I => \N__6013\
        );

    \I__667\ : Sp12to4
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__665\ : Span12Mux_h
    port map (
            O => \N__6010\,
            I => \N__6004\
        );

    \I__664\ : Span4Mux_h
    port map (
            O => \N__6007\,
            I => \N__6001\
        );

    \I__663\ : Span12Mux_h
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__662\ : Odrv4
    port map (
            O => \N__6001\,
            I => write_address_c_3
        );

    \I__661\ : Odrv12
    port map (
            O => \N__5998\,
            I => write_address_c_3
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__659\ : CascadeBuf
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__5987\,
            I => \N__5983\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__5986\,
            I => \N__5980\
        );

    \I__656\ : CascadeBuf
    port map (
            O => \N__5983\,
            I => \N__5977\
        );

    \I__655\ : CascadeBuf
    port map (
            O => \N__5980\,
            I => \N__5974\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__5977\,
            I => \N__5971\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__5974\,
            I => \N__5968\
        );

    \I__652\ : CascadeBuf
    port map (
            O => \N__5971\,
            I => \N__5965\
        );

    \I__651\ : CascadeBuf
    port map (
            O => \N__5968\,
            I => \N__5962\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \N__5959\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__5962\,
            I => \N__5956\
        );

    \I__648\ : CascadeBuf
    port map (
            O => \N__5959\,
            I => \N__5953\
        );

    \I__647\ : CascadeBuf
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__5953\,
            I => \N__5947\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__5950\,
            I => \N__5944\
        );

    \I__644\ : CascadeBuf
    port map (
            O => \N__5947\,
            I => \N__5941\
        );

    \I__643\ : CascadeBuf
    port map (
            O => \N__5944\,
            I => \N__5938\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__5941\,
            I => \N__5935\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__5938\,
            I => \N__5932\
        );

    \I__640\ : CascadeBuf
    port map (
            O => \N__5935\,
            I => \N__5929\
        );

    \I__639\ : CascadeBuf
    port map (
            O => \N__5932\,
            I => \N__5926\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__5929\,
            I => \N__5923\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__636\ : CascadeBuf
    port map (
            O => \N__5923\,
            I => \N__5917\
        );

    \I__635\ : CascadeBuf
    port map (
            O => \N__5920\,
            I => \N__5914\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__5917\,
            I => \N__5911\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__632\ : CascadeBuf
    port map (
            O => \N__5911\,
            I => \N__5905\
        );

    \I__631\ : CascadeBuf
    port map (
            O => \N__5908\,
            I => \N__5902\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__5905\,
            I => \N__5899\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__5902\,
            I => \N__5896\
        );

    \I__628\ : CascadeBuf
    port map (
            O => \N__5899\,
            I => \N__5893\
        );

    \I__627\ : CascadeBuf
    port map (
            O => \N__5896\,
            I => \N__5890\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__5893\,
            I => \N__5887\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__5890\,
            I => \N__5884\
        );

    \I__624\ : CascadeBuf
    port map (
            O => \N__5887\,
            I => \N__5881\
        );

    \I__623\ : CascadeBuf
    port map (
            O => \N__5884\,
            I => \N__5878\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__5881\,
            I => \N__5875\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__5878\,
            I => \N__5872\
        );

    \I__620\ : CascadeBuf
    port map (
            O => \N__5875\,
            I => \N__5869\
        );

    \I__619\ : CascadeBuf
    port map (
            O => \N__5872\,
            I => \N__5866\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__5869\,
            I => \N__5863\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__5866\,
            I => \N__5860\
        );

    \I__616\ : CascadeBuf
    port map (
            O => \N__5863\,
            I => \N__5857\
        );

    \I__615\ : CascadeBuf
    port map (
            O => \N__5860\,
            I => \N__5854\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__5857\,
            I => \N__5851\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__5854\,
            I => \N__5848\
        );

    \I__612\ : CascadeBuf
    port map (
            O => \N__5851\,
            I => \N__5845\
        );

    \I__611\ : CascadeBuf
    port map (
            O => \N__5848\,
            I => \N__5842\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__5842\,
            I => \N__5836\
        );

    \I__608\ : CascadeBuf
    port map (
            O => \N__5839\,
            I => \N__5833\
        );

    \I__607\ : CascadeBuf
    port map (
            O => \N__5836\,
            I => \N__5830\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__5833\,
            I => \N__5827\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__5830\,
            I => \N__5824\
        );

    \I__604\ : CascadeBuf
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__603\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5818\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__5821\,
            I => \N__5815\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__5818\,
            I => \N__5812\
        );

    \I__600\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5809\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__5812\,
            I => \N__5806\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5809\,
            I => \N__5803\
        );

    \I__597\ : Sp12to4
    port map (
            O => \N__5806\,
            I => \N__5800\
        );

    \I__596\ : Span12Mux_s1_v
    port map (
            O => \N__5803\,
            I => \N__5797\
        );

    \I__595\ : Span12Mux_h
    port map (
            O => \N__5800\,
            I => \N__5792\
        );

    \I__594\ : Span12Mux_h
    port map (
            O => \N__5797\,
            I => \N__5792\
        );

    \I__593\ : Odrv12
    port map (
            O => \N__5792\,
            I => write_address_c_2
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__5789\,
            I => \N__5786\
        );

    \I__591\ : CascadeBuf
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__589\ : CascadeBuf
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__5777\,
            I => \N__5773\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__5776\,
            I => \N__5770\
        );

    \I__586\ : CascadeBuf
    port map (
            O => \N__5773\,
            I => \N__5767\
        );

    \I__585\ : CascadeBuf
    port map (
            O => \N__5770\,
            I => \N__5764\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__5767\,
            I => \N__5761\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__5764\,
            I => \N__5758\
        );

    \I__582\ : CascadeBuf
    port map (
            O => \N__5761\,
            I => \N__5755\
        );

    \I__581\ : CascadeBuf
    port map (
            O => \N__5758\,
            I => \N__5752\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__5755\,
            I => \N__5749\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__578\ : CascadeBuf
    port map (
            O => \N__5749\,
            I => \N__5743\
        );

    \I__577\ : CascadeBuf
    port map (
            O => \N__5746\,
            I => \N__5740\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__5743\,
            I => \N__5737\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__5740\,
            I => \N__5734\
        );

    \I__574\ : CascadeBuf
    port map (
            O => \N__5737\,
            I => \N__5731\
        );

    \I__573\ : CascadeBuf
    port map (
            O => \N__5734\,
            I => \N__5728\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__5731\,
            I => \N__5725\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__5728\,
            I => \N__5722\
        );

    \I__570\ : CascadeBuf
    port map (
            O => \N__5725\,
            I => \N__5719\
        );

    \I__569\ : CascadeBuf
    port map (
            O => \N__5722\,
            I => \N__5716\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__5716\,
            I => \N__5710\
        );

    \I__566\ : CascadeBuf
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__565\ : CascadeBuf
    port map (
            O => \N__5710\,
            I => \N__5704\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__5704\,
            I => \N__5698\
        );

    \I__562\ : CascadeBuf
    port map (
            O => \N__5701\,
            I => \N__5695\
        );

    \I__561\ : CascadeBuf
    port map (
            O => \N__5698\,
            I => \N__5692\
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__5695\,
            I => \N__5689\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__5692\,
            I => \N__5686\
        );

    \I__558\ : CascadeBuf
    port map (
            O => \N__5689\,
            I => \N__5683\
        );

    \I__557\ : CascadeBuf
    port map (
            O => \N__5686\,
            I => \N__5680\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__5680\,
            I => \N__5674\
        );

    \I__554\ : CascadeBuf
    port map (
            O => \N__5677\,
            I => \N__5671\
        );

    \I__553\ : CascadeBuf
    port map (
            O => \N__5674\,
            I => \N__5668\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__5671\,
            I => \N__5665\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__5668\,
            I => \N__5662\
        );

    \I__550\ : CascadeBuf
    port map (
            O => \N__5665\,
            I => \N__5659\
        );

    \I__549\ : CascadeBuf
    port map (
            O => \N__5662\,
            I => \N__5656\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__5659\,
            I => \N__5653\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__5656\,
            I => \N__5650\
        );

    \I__546\ : CascadeBuf
    port map (
            O => \N__5653\,
            I => \N__5647\
        );

    \I__545\ : CascadeBuf
    port map (
            O => \N__5650\,
            I => \N__5644\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__5647\,
            I => \N__5641\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__5644\,
            I => \N__5638\
        );

    \I__542\ : CascadeBuf
    port map (
            O => \N__5641\,
            I => \N__5635\
        );

    \I__541\ : CascadeBuf
    port map (
            O => \N__5638\,
            I => \N__5632\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__5635\,
            I => \N__5629\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \N__5626\
        );

    \I__538\ : CascadeBuf
    port map (
            O => \N__5629\,
            I => \N__5623\
        );

    \I__537\ : CascadeBuf
    port map (
            O => \N__5626\,
            I => \N__5620\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__5623\,
            I => \N__5617\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__5620\,
            I => \N__5614\
        );

    \I__534\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5611\
        );

    \I__533\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5608\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5602\
        );

    \I__530\ : Span4Mux_s1_v
    port map (
            O => \N__5605\,
            I => \N__5599\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__5602\,
            I => \N__5596\
        );

    \I__528\ : Sp12to4
    port map (
            O => \N__5599\,
            I => \N__5593\
        );

    \I__527\ : IoSpan4Mux
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__526\ : Span12Mux_h
    port map (
            O => \N__5593\,
            I => \N__5587\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__5590\,
            I => write_address_c_10
        );

    \I__524\ : Odrv12
    port map (
            O => \N__5587\,
            I => write_address_c_10
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__522\ : CascadeBuf
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__520\ : CascadeBuf
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__518\ : CascadeBuf
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__516\ : CascadeBuf
    port map (
            O => \N__5561\,
            I => \N__5557\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__5560\,
            I => \N__5554\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__5557\,
            I => \N__5551\
        );

    \I__513\ : CascadeBuf
    port map (
            O => \N__5554\,
            I => \N__5548\
        );

    \I__512\ : CascadeBuf
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__5548\,
            I => \N__5542\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__5545\,
            I => \N__5539\
        );

    \I__509\ : CascadeBuf
    port map (
            O => \N__5542\,
            I => \N__5536\
        );

    \I__508\ : CascadeBuf
    port map (
            O => \N__5539\,
            I => \N__5533\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__5533\,
            I => \N__5527\
        );

    \I__505\ : CascadeBuf
    port map (
            O => \N__5530\,
            I => \N__5524\
        );

    \I__504\ : CascadeBuf
    port map (
            O => \N__5527\,
            I => \N__5521\
        );

    \I__503\ : CascadeMux
    port map (
            O => \N__5524\,
            I => \N__5518\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__5521\,
            I => \N__5515\
        );

    \I__501\ : CascadeBuf
    port map (
            O => \N__5518\,
            I => \N__5512\
        );

    \I__500\ : CascadeBuf
    port map (
            O => \N__5515\,
            I => \N__5509\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__5512\,
            I => \N__5506\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__5509\,
            I => \N__5503\
        );

    \I__497\ : CascadeBuf
    port map (
            O => \N__5506\,
            I => \N__5500\
        );

    \I__496\ : CascadeBuf
    port map (
            O => \N__5503\,
            I => \N__5497\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__5500\,
            I => \N__5494\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__5497\,
            I => \N__5491\
        );

    \I__493\ : CascadeBuf
    port map (
            O => \N__5494\,
            I => \N__5488\
        );

    \I__492\ : CascadeBuf
    port map (
            O => \N__5491\,
            I => \N__5485\
        );

    \I__491\ : CascadeMux
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__5485\,
            I => \N__5479\
        );

    \I__489\ : CascadeBuf
    port map (
            O => \N__5482\,
            I => \N__5476\
        );

    \I__488\ : CascadeBuf
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__5476\,
            I => \N__5470\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__5473\,
            I => \N__5467\
        );

    \I__485\ : CascadeBuf
    port map (
            O => \N__5470\,
            I => \N__5464\
        );

    \I__484\ : CascadeBuf
    port map (
            O => \N__5467\,
            I => \N__5461\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__5464\,
            I => \N__5458\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__5461\,
            I => \N__5455\
        );

    \I__481\ : CascadeBuf
    port map (
            O => \N__5458\,
            I => \N__5452\
        );

    \I__480\ : CascadeBuf
    port map (
            O => \N__5455\,
            I => \N__5449\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__5452\,
            I => \N__5446\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__5449\,
            I => \N__5443\
        );

    \I__477\ : CascadeBuf
    port map (
            O => \N__5446\,
            I => \N__5440\
        );

    \I__476\ : CascadeBuf
    port map (
            O => \N__5443\,
            I => \N__5437\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__5440\,
            I => \N__5434\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__5437\,
            I => \N__5431\
        );

    \I__473\ : CascadeBuf
    port map (
            O => \N__5434\,
            I => \N__5428\
        );

    \I__472\ : CascadeBuf
    port map (
            O => \N__5431\,
            I => \N__5425\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__5428\,
            I => \N__5422\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__5425\,
            I => \N__5419\
        );

    \I__469\ : CascadeBuf
    port map (
            O => \N__5422\,
            I => \N__5416\
        );

    \I__468\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5413\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__5416\,
            I => \N__5410\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__5413\,
            I => \N__5407\
        );

    \I__465\ : CascadeBuf
    port map (
            O => \N__5410\,
            I => \N__5404\
        );

    \I__464\ : Span4Mux_s3_v
    port map (
            O => \N__5407\,
            I => \N__5401\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__5404\,
            I => \N__5398\
        );

    \I__462\ : Span4Mux_h
    port map (
            O => \N__5401\,
            I => \N__5395\
        );

    \I__461\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5392\
        );

    \I__460\ : Sp12to4
    port map (
            O => \N__5395\,
            I => \N__5389\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5386\
        );

    \I__458\ : Span12Mux_h
    port map (
            O => \N__5389\,
            I => \N__5383\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__5386\,
            I => write_address_c_1
        );

    \I__456\ : Odrv12
    port map (
            O => \N__5383\,
            I => write_address_c_1
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__454\ : CascadeBuf
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__5372\,
            I => \N__5368\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__451\ : CascadeBuf
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__450\ : CascadeBuf
    port map (
            O => \N__5365\,
            I => \N__5359\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \N__5356\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__447\ : CascadeBuf
    port map (
            O => \N__5356\,
            I => \N__5350\
        );

    \I__446\ : CascadeBuf
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__5347\,
            I => \N__5341\
        );

    \I__443\ : CascadeBuf
    port map (
            O => \N__5344\,
            I => \N__5338\
        );

    \I__442\ : CascadeBuf
    port map (
            O => \N__5341\,
            I => \N__5335\
        );

    \I__441\ : CascadeMux
    port map (
            O => \N__5338\,
            I => \N__5332\
        );

    \I__440\ : CascadeMux
    port map (
            O => \N__5335\,
            I => \N__5329\
        );

    \I__439\ : CascadeBuf
    port map (
            O => \N__5332\,
            I => \N__5326\
        );

    \I__438\ : CascadeBuf
    port map (
            O => \N__5329\,
            I => \N__5323\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__5326\,
            I => \N__5320\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__5323\,
            I => \N__5317\
        );

    \I__435\ : CascadeBuf
    port map (
            O => \N__5320\,
            I => \N__5314\
        );

    \I__434\ : CascadeBuf
    port map (
            O => \N__5317\,
            I => \N__5311\
        );

    \I__433\ : CascadeMux
    port map (
            O => \N__5314\,
            I => \N__5308\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__5311\,
            I => \N__5305\
        );

    \I__431\ : CascadeBuf
    port map (
            O => \N__5308\,
            I => \N__5302\
        );

    \I__430\ : CascadeBuf
    port map (
            O => \N__5305\,
            I => \N__5299\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__5302\,
            I => \N__5296\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__5299\,
            I => \N__5293\
        );

    \I__427\ : CascadeBuf
    port map (
            O => \N__5296\,
            I => \N__5290\
        );

    \I__426\ : CascadeBuf
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__5287\,
            I => \N__5281\
        );

    \I__423\ : CascadeBuf
    port map (
            O => \N__5284\,
            I => \N__5278\
        );

    \I__422\ : CascadeBuf
    port map (
            O => \N__5281\,
            I => \N__5275\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__5278\,
            I => \N__5272\
        );

    \I__420\ : CascadeMux
    port map (
            O => \N__5275\,
            I => \N__5269\
        );

    \I__419\ : CascadeBuf
    port map (
            O => \N__5272\,
            I => \N__5266\
        );

    \I__418\ : CascadeBuf
    port map (
            O => \N__5269\,
            I => \N__5263\
        );

    \I__417\ : CascadeMux
    port map (
            O => \N__5266\,
            I => \N__5260\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__5263\,
            I => \N__5257\
        );

    \I__415\ : CascadeBuf
    port map (
            O => \N__5260\,
            I => \N__5254\
        );

    \I__414\ : CascadeBuf
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__5254\,
            I => \N__5248\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__5251\,
            I => \N__5245\
        );

    \I__411\ : CascadeBuf
    port map (
            O => \N__5248\,
            I => \N__5242\
        );

    \I__410\ : CascadeBuf
    port map (
            O => \N__5245\,
            I => \N__5239\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__5242\,
            I => \N__5236\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__5239\,
            I => \N__5233\
        );

    \I__407\ : CascadeBuf
    port map (
            O => \N__5236\,
            I => \N__5230\
        );

    \I__406\ : CascadeBuf
    port map (
            O => \N__5233\,
            I => \N__5227\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__5230\,
            I => \N__5224\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__5227\,
            I => \N__5221\
        );

    \I__403\ : CascadeBuf
    port map (
            O => \N__5224\,
            I => \N__5218\
        );

    \I__402\ : CascadeBuf
    port map (
            O => \N__5221\,
            I => \N__5215\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__5218\,
            I => \N__5212\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__5215\,
            I => \N__5209\
        );

    \I__399\ : CascadeBuf
    port map (
            O => \N__5212\,
            I => \N__5206\
        );

    \I__398\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5203\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__5206\,
            I => \N__5200\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5197\
        );

    \I__395\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5194\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__5197\,
            I => \N__5191\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__5194\,
            I => \N__5188\
        );

    \I__392\ : Sp12to4
    port map (
            O => \N__5191\,
            I => \N__5185\
        );

    \I__391\ : Span4Mux_h
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__390\ : Span12Mux_h
    port map (
            O => \N__5185\,
            I => \N__5179\
        );

    \I__389\ : Span4Mux_h
    port map (
            O => \N__5182\,
            I => \N__5176\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__5179\,
            I => write_address_c_0
        );

    \I__387\ : Odrv4
    port map (
            O => \N__5176\,
            I => write_address_c_0
        );

    \I__386\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__384\ : Span4Mux_s3_v
    port map (
            O => \N__5165\,
            I => \N__5161\
        );

    \I__383\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5158\
        );

    \I__382\ : Span4Mux_v
    port map (
            O => \N__5161\,
            I => \N__5151\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__5158\,
            I => \N__5151\
        );

    \I__380\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5148\
        );

    \I__379\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5145\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__5151\,
            I => \N__5139\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__5148\,
            I => \N__5139\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__5145\,
            I => \N__5136\
        );

    \I__375\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5133\
        );

    \I__374\ : Span4Mux_v
    port map (
            O => \N__5139\,
            I => \N__5130\
        );

    \I__373\ : Span4Mux_v
    port map (
            O => \N__5136\,
            I => \N__5125\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__5133\,
            I => \N__5125\
        );

    \I__371\ : Span4Mux_v
    port map (
            O => \N__5130\,
            I => \N__5119\
        );

    \I__370\ : Span4Mux_v
    port map (
            O => \N__5125\,
            I => \N__5119\
        );

    \I__369\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5114\
        );

    \I__368\ : Span4Mux_h
    port map (
            O => \N__5119\,
            I => \N__5109\
        );

    \I__367\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5106\
        );

    \I__366\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5103\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__5114\,
            I => \N__5100\
        );

    \I__364\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5097\
        );

    \I__363\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5094\
        );

    \I__362\ : Sp12to4
    port map (
            O => \N__5109\,
            I => \N__5091\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__5106\,
            I => \N__5086\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__5103\,
            I => \N__5086\
        );

    \I__359\ : Span12Mux_s7_v
    port map (
            O => \N__5100\,
            I => \N__5079\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__5097\,
            I => \N__5079\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__5094\,
            I => \N__5079\
        );

    \I__356\ : Span12Mux_h
    port map (
            O => \N__5091\,
            I => \N__5072\
        );

    \I__355\ : Span12Mux_v
    port map (
            O => \N__5086\,
            I => \N__5072\
        );

    \I__354\ : Span12Mux_v
    port map (
            O => \N__5079\,
            I => \N__5072\
        );

    \I__353\ : Odrv12
    port map (
            O => \N__5072\,
            I => write_data_c_5
        );

    \I__352\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__5066\,
            I => \N__5062\
        );

    \I__350\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5059\
        );

    \I__349\ : Span4Mux_v
    port map (
            O => \N__5062\,
            I => \N__5054\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__5059\,
            I => \N__5054\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__346\ : Span4Mux_v
    port map (
            O => \N__5051\,
            I => \N__5047\
        );

    \I__345\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5044\
        );

    \I__344\ : Span4Mux_v
    port map (
            O => \N__5047\,
            I => \N__5038\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__5044\,
            I => \N__5038\
        );

    \I__342\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5033\
        );

    \I__341\ : Span4Mux_v
    port map (
            O => \N__5038\,
            I => \N__5030\
        );

    \I__340\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5026\
        );

    \I__339\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5022\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__5033\,
            I => \N__5019\
        );

    \I__337\ : Span4Mux_h
    port map (
            O => \N__5030\,
            I => \N__5016\
        );

    \I__336\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5013\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__5026\,
            I => \N__5010\
        );

    \I__334\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5007\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__5022\,
            I => \N__5004\
        );

    \I__332\ : Span12Mux_h
    port map (
            O => \N__5019\,
            I => \N__4999\
        );

    \I__331\ : Span4Mux_v
    port map (
            O => \N__5016\,
            I => \N__4996\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__5013\,
            I => \N__4993\
        );

    \I__329\ : Span12Mux_s4_v
    port map (
            O => \N__5010\,
            I => \N__4988\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__5007\,
            I => \N__4988\
        );

    \I__327\ : Span4Mux_v
    port map (
            O => \N__5004\,
            I => \N__4985\
        );

    \I__326\ : InMux
    port map (
            O => \N__5003\,
            I => \N__4982\
        );

    \I__325\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4979\
        );

    \I__324\ : Span12Mux_v
    port map (
            O => \N__4999\,
            I => \N__4972\
        );

    \I__323\ : Sp12to4
    port map (
            O => \N__4996\,
            I => \N__4972\
        );

    \I__322\ : Span12Mux_h
    port map (
            O => \N__4993\,
            I => \N__4972\
        );

    \I__321\ : Span12Mux_v
    port map (
            O => \N__4988\,
            I => \N__4963\
        );

    \I__320\ : Sp12to4
    port map (
            O => \N__4985\,
            I => \N__4963\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__4982\,
            I => \N__4963\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4963\
        );

    \I__317\ : Span12Mux_h
    port map (
            O => \N__4972\,
            I => \N__4958\
        );

    \I__316\ : Span12Mux_v
    port map (
            O => \N__4963\,
            I => \N__4958\
        );

    \I__315\ : Odrv12
    port map (
            O => \N__4958\,
            I => write_data_c_4
        );

    \I__314\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4951\
        );

    \I__313\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4948\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__4951\,
            I => \N__4945\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__4948\,
            I => \N__4941\
        );

    \I__310\ : Span4Mux_s2_v
    port map (
            O => \N__4945\,
            I => \N__4937\
        );

    \I__309\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4934\
        );

    \I__308\ : Span4Mux_s3_v
    port map (
            O => \N__4941\,
            I => \N__4931\
        );

    \I__307\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4928\
        );

    \I__306\ : Span4Mux_v
    port map (
            O => \N__4937\,
            I => \N__4921\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__4934\,
            I => \N__4921\
        );

    \I__304\ : Span4Mux_v
    port map (
            O => \N__4931\,
            I => \N__4914\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4914\
        );

    \I__302\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4911\
        );

    \I__301\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4908\
        );

    \I__300\ : Span4Mux_h
    port map (
            O => \N__4921\,
            I => \N__4904\
        );

    \I__299\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4901\
        );

    \I__298\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4898\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__4914\,
            I => \N__4893\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4893\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4890\
        );

    \I__294\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4887\
        );

    \I__293\ : Span4Mux_v
    port map (
            O => \N__4904\,
            I => \N__4882\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4882\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4879\
        );

    \I__290\ : Span4Mux_v
    port map (
            O => \N__4893\,
            I => \N__4875\
        );

    \I__289\ : Span4Mux_v
    port map (
            O => \N__4890\,
            I => \N__4870\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__4887\,
            I => \N__4870\
        );

    \I__287\ : Span4Mux_v
    port map (
            O => \N__4882\,
            I => \N__4867\
        );

    \I__286\ : Span4Mux_v
    port map (
            O => \N__4879\,
            I => \N__4864\
        );

    \I__285\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4861\
        );

    \I__284\ : Span4Mux_v
    port map (
            O => \N__4875\,
            I => \N__4856\
        );

    \I__283\ : Span4Mux_v
    port map (
            O => \N__4870\,
            I => \N__4856\
        );

    \I__282\ : Span4Mux_v
    port map (
            O => \N__4867\,
            I => \N__4849\
        );

    \I__281\ : Span4Mux_v
    port map (
            O => \N__4864\,
            I => \N__4849\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__4861\,
            I => \N__4849\
        );

    \I__279\ : Sp12to4
    port map (
            O => \N__4856\,
            I => \N__4846\
        );

    \I__278\ : Span4Mux_h
    port map (
            O => \N__4849\,
            I => \N__4843\
        );

    \I__277\ : Span12Mux_h
    port map (
            O => \N__4846\,
            I => \N__4840\
        );

    \I__276\ : IoSpan4Mux
    port map (
            O => \N__4843\,
            I => \N__4837\
        );

    \I__275\ : Odrv12
    port map (
            O => \N__4840\,
            I => write_data_c_3
        );

    \I__274\ : Odrv4
    port map (
            O => \N__4837\,
            I => write_data_c_3
        );

    \I__273\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__4829\,
            I => \N__4825\
        );

    \I__271\ : InMux
    port map (
            O => \N__4828\,
            I => \N__4822\
        );

    \I__270\ : Span4Mux_v
    port map (
            O => \N__4825\,
            I => \N__4817\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__4822\,
            I => \N__4817\
        );

    \I__268\ : Span4Mux_v
    port map (
            O => \N__4817\,
            I => \N__4812\
        );

    \I__267\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4809\
        );

    \I__266\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4805\
        );

    \I__265\ : Span4Mux_v
    port map (
            O => \N__4812\,
            I => \N__4799\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4799\
        );

    \I__263\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4796\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4793\
        );

    \I__261\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4790\
        );

    \I__260\ : Span4Mux_v
    port map (
            O => \N__4799\,
            I => \N__4785\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__4796\,
            I => \N__4785\
        );

    \I__258\ : Span4Mux_v
    port map (
            O => \N__4793\,
            I => \N__4779\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__4790\,
            I => \N__4779\
        );

    \I__256\ : Span4Mux_v
    port map (
            O => \N__4785\,
            I => \N__4775\
        );

    \I__255\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4772\
        );

    \I__254\ : Span4Mux_v
    port map (
            O => \N__4779\,
            I => \N__4769\
        );

    \I__253\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4766\
        );

    \I__252\ : Span4Mux_v
    port map (
            O => \N__4775\,
            I => \N__4760\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4760\
        );

    \I__250\ : Span4Mux_v
    port map (
            O => \N__4769\,
            I => \N__4755\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__4766\,
            I => \N__4755\
        );

    \I__248\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4752\
        );

    \I__247\ : Span4Mux_v
    port map (
            O => \N__4760\,
            I => \N__4749\
        );

    \I__246\ : Span4Mux_v
    port map (
            O => \N__4755\,
            I => \N__4744\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__4752\,
            I => \N__4744\
        );

    \I__244\ : Span4Mux_h
    port map (
            O => \N__4749\,
            I => \N__4740\
        );

    \I__243\ : Span4Mux_v
    port map (
            O => \N__4744\,
            I => \N__4737\
        );

    \I__242\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4734\
        );

    \I__241\ : Sp12to4
    port map (
            O => \N__4740\,
            I => \N__4731\
        );

    \I__240\ : Span4Mux_v
    port map (
            O => \N__4737\,
            I => \N__4726\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__4734\,
            I => \N__4726\
        );

    \I__238\ : Span12Mux_h
    port map (
            O => \N__4731\,
            I => \N__4723\
        );

    \I__237\ : Span4Mux_v
    port map (
            O => \N__4726\,
            I => \N__4720\
        );

    \I__236\ : Odrv12
    port map (
            O => \N__4723\,
            I => write_data_c_2
        );

    \I__235\ : Odrv4
    port map (
            O => \N__4720\,
            I => write_data_c_2
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_6_cry_7\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.address_1_0_8\,
            carryinitout => \bfn_13_18_0_\
        );

    \this_reset_cond.M_stage_q_RNI6VB7_3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12070\,
            GLOBALBUFFEROUTPUT => \N_112_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNI1P4R_0_0_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__11797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12139\,
            lcout => \this_vga_signals_N_170_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11784\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12126\,
            lcout => \this_vga_signals_N_171_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNIUAUT_0_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12140\,
            in1 => \N__10471\,
            in2 => \N__10520\,
            in3 => \N__11798\,
            lcout => rgb5_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNITHP2_0_0_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__10472\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10519\,
            lcout => vsync_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNITHP2_0_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10465\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10515\,
            lcout => \this_vga_signals_N_94_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNILGF11_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14436\,
            in1 => \N__7808\,
            in2 => \_gnd_net_\,
            in3 => \N__7796\,
            lcout => \this_vram.mem_mem_0_0_RNILGFZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNINGF11_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7790\,
            in1 => \N__14477\,
            in2 => \_gnd_net_\,
            in3 => \N__7778\,
            lcout => \this_vram.mem_mem_0_1_RNINGFZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNINGF11_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14476\,
            in1 => \N__8036\,
            in2 => \_gnd_net_\,
            in3 => \N__8024\,
            lcout => \this_vram.mem_mem_0_1_RNINGF11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_2_RNIPGF11_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8018\,
            in1 => \N__14463\,
            in2 => \_gnd_net_\,
            in3 => \N__8006\,
            lcout => \this_vram.mem_mem_0_2_RNIPGFZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_2_RNIPGF11_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14462\,
            in1 => \N__8000\,
            in2 => \_gnd_net_\,
            in3 => \N__7994\,
            lcout => \this_vram.mem_mem_0_2_RNIPGF11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIPOJ11_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7982\,
            in1 => \N__14456\,
            in2 => \_gnd_net_\,
            in3 => \N__7970\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_0_RNIPOJZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNINVA72_0_12_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__7964\,
            in1 => \_gnd_net_\,
            in2 => \N__7955\,
            in3 => \N__14175\,
            lcout => \this_vram.mem_N_2362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OEJ4_0_13_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8381\,
            in1 => \N__7952\,
            in2 => \_gnd_net_\,
            in3 => \N__10273\,
            lcout => OPEN,
            ltout => \this_vram.mem_N_2364_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIN7E66_0_14_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__8732\,
            in1 => \N__13946\,
            in2 => \N__7943\,
            in3 => \N__10202\,
            lcout => \M_this_vram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNIROJ11_0_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7928\,
            in1 => \N__14361\,
            in2 => \_gnd_net_\,
            in3 => \N__7916\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_1_RNIROJ11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIRVA72_12_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__8165\,
            in1 => \_gnd_net_\,
            in2 => \N__8156\,
            in3 => \N__14097\,
            lcout => \this_vram.mem_N_2335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_1_RNI14P11_0_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14171\,
            in1 => \N__8153\,
            in2 => \_gnd_net_\,
            in3 => \N__8138\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_4_1_RNI14P11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIC1S72_11_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__12749\,
            in1 => \_gnd_net_\,
            in2 => \N__8117\,
            in3 => \N__14453\,
            lcout => OPEN,
            ltout => \this_vram.mem_N_2336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIHOEJ4_13_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10293\,
            in1 => \_gnd_net_\,
            in2 => \N__8114\,
            in3 => \N__8111\,
            lcout => \this_vram.mem_N_2337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNIROJ11_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8105\,
            in1 => \N__14452\,
            in2 => \_gnd_net_\,
            in3 => \N__8093\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_1_RNIROJZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIRVA72_0_12_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__14172\,
            in1 => \_gnd_net_\,
            in2 => \N__8087\,
            in3 => \N__8084\,
            lcout => \this_vram.mem_N_2344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_2_RNITOJ11_0_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8072\,
            in1 => \N__14454\,
            in2 => \_gnd_net_\,
            in3 => \N__8060\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_2_RNITOJ11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIVVA72_12_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8054\,
            in2 => \N__8042\,
            in3 => \N__14173\,
            lcout => OPEN,
            ltout => \this_vram.mem_N_2371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIPOEJ4_13_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__10294\,
            in1 => \_gnd_net_\,
            in2 => \N__8039\,
            in3 => \N__13466\,
            lcout => \this_vram.mem_N_2373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_2_RNITOJ11_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8318\,
            in1 => \N__14455\,
            in2 => \_gnd_net_\,
            in3 => \N__8312\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_2_RNITOJZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIVVA72_0_12_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__14174\,
            in1 => \N__8300\,
            in2 => \N__8288\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_vram.mem_N_2326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIPOEJ4_0_13_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__10295\,
            in1 => \N__8765\,
            in2 => \N__8285\,
            in3 => \_gnd_net_\,
            lcout => \this_vram.mem_N_2328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIB8E66_14_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__10230\,
            in1 => \N__12827\,
            in2 => \N__8282\,
            in3 => \N__8733\,
            lcout => \M_this_vram_read_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIB8E66_0_14_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__8252\,
            in1 => \N__14267\,
            in2 => \N__8741\,
            in3 => \N__10232\,
            lcout => \M_this_vram_read_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI18E66_14_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__8225\,
            in1 => \N__14492\,
            in2 => \N__8740\,
            in3 => \N__10231\,
            lcout => \M_this_vram_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNILGF11_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14435\,
            in1 => \N__8201\,
            in2 => \_gnd_net_\,
            in3 => \N__8189\,
            lcout => \this_vram.mem_mem_0_0_RNILGF11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIPOJ11_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8183\,
            in1 => \N__14425\,
            in2 => \_gnd_net_\,
            in3 => \N__8171\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_0_RNIPOJ11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNINVA72_12_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8507\,
            in2 => \N__8498\,
            in3 => \N__14157\,
            lcout => \this_vram.mem_N_2353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_RNIV3P11_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8495\,
            in1 => \N__14095\,
            in2 => \_gnd_net_\,
            in3 => \N__8474\,
            lcout => \this_vram.mem_mem_4_0_RNIV3PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_wclke_0_a2_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14804\,
            in1 => \N__14900\,
            in2 => \N__14681\,
            in3 => \N__13864\,
            lcout => \this_vram.mem_WE_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_0_RNI18R11_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14096\,
            in1 => \N__8429\,
            in2 => \_gnd_net_\,
            in3 => \N__8408\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_5_0_RNI18RZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI81S72_0_11_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__14357\,
            in1 => \_gnd_net_\,
            in2 => \N__8390\,
            in3 => \N__8387\,
            lcout => \this_vram.mem_N_2363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIHOEJ4_0_13_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10281\,
            in1 => \N__8813\,
            in2 => \_gnd_net_\,
            in3 => \N__8369\,
            lcout => \this_vram.mem_N_2346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIU5NC_13_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__10215\,
            in1 => \N__10282\,
            in2 => \_gnd_net_\,
            in3 => \N__14161\,
            lcout => \this_vram.mem_G_25_0\,
            ltout => \this_vram.mem_G_25_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI18E66_0_14_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__13880\,
            in1 => \N__8360\,
            in2 => \N__8354\,
            in3 => \N__10214\,
            lcout => \M_this_vram_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_wclke_0_a2_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__14803\,
            in1 => \N__14895\,
            in2 => \N__13860\,
            in3 => \N__14676\,
            lcout => \this_vram.mem_WE_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIG1S72_0_11_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14201\,
            in1 => \N__8654\,
            in2 => \_gnd_net_\,
            in3 => \N__14431\,
            lcout => \this_vram.mem_N_2327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OEJ4_13_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10283\,
            in1 => \N__8543\,
            in2 => \_gnd_net_\,
            in3 => \N__8756\,
            lcout => OPEN,
            ltout => \this_vram.mem_N_2355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIN7E66_14_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__10216\,
            in1 => \N__13913\,
            in2 => \N__8744\,
            in3 => \N__8712\,
            lcout => \M_this_vram_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_2_RNI34P11_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8690\,
            in1 => \N__14170\,
            in2 => \_gnd_net_\,
            in3 => \N__8675\,
            lcout => \this_vram.mem_mem_4_2_RNI34PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_wclke_0_a2_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14793\,
            in1 => \N__14885\,
            in2 => \N__13859\,
            in3 => \N__14675\,
            lcout => \this_vram.mem_WE_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_RNIV3P11_0_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8621\,
            in1 => \N__8600\,
            in2 => \_gnd_net_\,
            in3 => \N__14176\,
            lcout => \this_vram.mem_mem_4_0_RNIV3P11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_0_RNI18R11_0_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8588\,
            in1 => \N__14177\,
            in2 => \_gnd_net_\,
            in3 => \N__8573\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_5_0_RNI18R11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI81S72_11_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__8552\,
            in1 => \_gnd_net_\,
            in2 => \N__8546\,
            in3 => \N__14464\,
            lcout => \this_vram.mem_N_2354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_wclke_0_a2_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__14680\,
            in1 => \N__14899\,
            in2 => \N__13865\,
            in3 => \N__14784\,
            lcout => \this_vram.mem_WE_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_1_RNI14P11_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8852\,
            in1 => \N__14141\,
            in2 => \_gnd_net_\,
            in3 => \N__8837\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_4_1_RNI14PZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIC1S72_0_11_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__12788\,
            in1 => \_gnd_net_\,
            in2 => \N__8816\,
            in3 => \N__14407\,
            lcout => \this_vram.mem_N_2345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_wclke_0_a2_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__14774\,
            in1 => \N__14864\,
            in2 => \N__13858\,
            in3 => \N__14659\,
            lcout => \this_vram.mem_WE_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m24_0_o2_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10792\,
            in2 => \_gnd_net_\,
            in3 => \N__10729\,
            lcout => \this_vga_signals.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_1_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__10730\,
            in1 => \N__10834\,
            in2 => \_gnd_net_\,
            in3 => \N__10793\,
            lcout => \this_vga_signals.m27_0_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__10539\,
            in1 => \N__10409\,
            in2 => \N__10462\,
            in3 => \N__10309\,
            lcout => OPEN,
            ltout => \this_vga_signals.m24_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m24_0_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111001"
        )
    port map (
            in0 => \N__10500\,
            in1 => \N__8771\,
            in2 => \N__8777\,
            in3 => \N__9715\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_0_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__12076\,
            in1 => \N__10501\,
            in2 => \N__8774\,
            in3 => \N__10680\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_0_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001010110"
        )
    port map (
            in0 => \N__10498\,
            in1 => \N__9730\,
            in2 => \N__10464\,
            in3 => \N__10842\,
            lcout => \this_vga_signals.m24_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m27_0_0_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101100000011"
        )
    port map (
            in0 => \N__10540\,
            in1 => \N__10499\,
            in2 => \N__10463\,
            in3 => \N__10310\,
            lcout => OPEN,
            ltout => \this_vga_signals.m27_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m27_0_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110100"
        )
    port map (
            in0 => \N__10453\,
            in1 => \N__9731\,
            in2 => \N__9722\,
            in3 => \N__9716\,
            lcout => OPEN,
            ltout => \this_vga_signals.i9_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_1_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__12077\,
            in1 => \N__10454\,
            in2 => \N__9719\,
            in3 => \N__10681\,
            lcout => \this_vga_signals.M_vstate_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__11986\,
            in1 => \N__10933\,
            in2 => \_gnd_net_\,
            in3 => \N__10322\,
            lcout => \this_vga_signals.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI8NSN1_2_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10788\,
            in2 => \N__9758\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \this_vga_signals.address_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_cry_0_c_RNI17SC1_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10728\,
            in2 => \N__9743\,
            in3 => \N__9293\,
            lcout => \M_this_vga_signals_address_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_cry_0\,
            carryout => \this_vga_signals.address_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_cry_1_c_RNI5DUC1_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10682\,
            in2 => \N__10388\,
            in3 => \N__9074\,
            lcout => \M_this_vga_signals_address_9\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_cry_1\,
            carryout => \this_vga_signals.address_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_cry_2_c_RNI9J0D1_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10637\,
            in2 => \N__10373\,
            in3 => \N__8858\,
            lcout => \M_this_vga_signals_address_10\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_cry_2\,
            carryout => \this_vga_signals.address_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_11_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10358\,
            in2 => \N__10601\,
            in3 => \N__8855\,
            lcout => \this_vram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_cry_3\,
            carryout => \this_vga_signals.address_1_cry_4\,
            clk => \N__13676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_12_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10346\,
            in2 => \N__10973\,
            in3 => \N__10298\,
            lcout => \this_vram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_cry_4\,
            carryout => \this_vga_signals.address_1_cry_5\,
            clk => \N__13676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_13_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10331\,
            in2 => \N__10934\,
            in3 => \N__10238\,
            lcout => \this_vram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_cry_5\,
            carryout => \this_vga_signals.address_1_cry_6\,
            clk => \N__13676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_14_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11987\,
            in2 => \_gnd_net_\,
            in3 => \N__10235\,
            lcout => \this_vram.mem_radregZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_2_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__12015\,
            in1 => \N__10797\,
            in2 => \N__11936\,
            in3 => \N__10751\,
            lcout => \this_vga_signals.address_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_3_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__10737\,
            in1 => \N__12016\,
            in2 => \N__10697\,
            in3 => \N__11933\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNINV7N_9_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10787\,
            in2 => \N__11747\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \this_vga_signals.address_1_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_cry_0_c_RNIM2N91_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10727\,
            in2 => \N__11712\,
            in3 => \N__9761\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_0_cry_0\,
            carryout => \this_vga_signals.address_1_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_cry_1_c_RNIP6O91_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10666\,
            in2 => \N__12490\,
            in3 => \N__9746\,
            lcout => \this_vga_signals.address_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_0_cry_1\,
            carryout => \this_vga_signals.address_1_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_cry_2_c_RNIADGT_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10636\,
            in3 => \N__10391\,
            lcout => \this_vga_signals.address_1_0_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_0_cry_2\,
            carryout => \this_vga_signals.address_1_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_cry_3_c_RNICGHT_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10588\,
            in2 => \_gnd_net_\,
            in3 => \N__10376\,
            lcout => \this_vga_signals.address_1_0_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_0_cry_3\,
            carryout => \this_vga_signals.address_1_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_cry_4_c_RNIEJIT_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10960\,
            in2 => \_gnd_net_\,
            in3 => \N__10361\,
            lcout => \this_vga_signals.address_1_0_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_0_cry_4\,
            carryout => \this_vga_signals.address_1_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_cry_5_c_RNIGMJT_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10923\,
            in2 => \_gnd_net_\,
            in3 => \N__10349\,
            lcout => \this_vga_signals.address_1_0_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_0_cry_5\,
            carryout => \this_vga_signals.address_1_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_cry_6_c_RNIIPKT_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11984\,
            in2 => \_gnd_net_\,
            in3 => \N__10337\,
            lcout => \this_vga_signals.address_1_0_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.address_1_0_cry_6\,
            carryout => \this_vga_signals.address_1_0_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.address_1_0_8_THRU_LUT4_0_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10334\,
            lcout => \this_vga_signals.address_1_0_8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_3_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__10961\,
            in1 => \N__10589\,
            in2 => \N__10869\,
            in3 => \N__10630\,
            lcout => \this_vga_signals.m27_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_5_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10631\,
            in1 => \N__10862\,
            in2 => \N__10843\,
            in3 => \N__10316\,
            lcout => \this_vga_signals.m27_0_a2_1_5\,
            ltout => \this_vga_signals.m27_0_a2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNICG7G4_1_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10443\,
            in1 => \N__10526\,
            in2 => \N__10301\,
            in3 => \N__10541\,
            lcout => \this_vga_signals.N_68\,
            ltout => \this_vga_signals.N_68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_1_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__10838\,
            in1 => \N__11929\,
            in2 => \N__10544\,
            in3 => \N__10811\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_4_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10962\,
            in1 => \N__10918\,
            in2 => \N__11985\,
            in3 => \N__10590\,
            lcout => \this_vga_signals.m27_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_RNIVAHF_0_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10496\,
            in2 => \_gnd_net_\,
            in3 => \N__10670\,
            lcout => \this_vga_signals.M_vcounter_q_0_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vstate_q_ns_1_0__m24_0_0_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010100"
        )
    port map (
            in0 => \N__10497\,
            in1 => \N__10799\,
            in2 => \N__10461\,
            in3 => \N__10739\,
            lcout => \this_vga_signals.m24_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11865\,
            in2 => \N__11834\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11846\,
            in2 => \_gnd_net_\,
            in3 => \N__10403\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__13673\,
            ce => 'H',
            sr => \N__11908\
        );

    \this_vga_signals.M_hcounter_q_3_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11810\,
            in2 => \_gnd_net_\,
            in3 => \N__10400\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__13673\,
            ce => 'H',
            sr => \N__11908\
        );

    \this_vga_signals.M_hcounter_q_4_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12520\,
            in2 => \_gnd_net_\,
            in3 => \N__10397\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__13673\,
            ce => 'H',
            sr => \N__11908\
        );

    \this_vga_signals.M_hcounter_q_5_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12271\,
            in2 => \_gnd_net_\,
            in3 => \N__10394\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__13673\,
            ce => 'H',
            sr => \N__11908\
        );

    \this_vga_signals.M_hcounter_q_6_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11481\,
            in2 => \_gnd_net_\,
            in3 => \N__10562\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__13673\,
            ce => 'H',
            sr => \N__11908\
        );

    \this_vga_signals.M_hcounter_q_7_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12227\,
            in1 => \N__11251\,
            in2 => \_gnd_net_\,
            in3 => \N__10559\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__13673\,
            ce => 'H',
            sr => \N__11908\
        );

    \this_vga_signals.M_hcounter_q_8_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11010\,
            in2 => \_gnd_net_\,
            in3 => \N__10556\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__13673\,
            ce => 'H',
            sr => \N__11908\
        );

    \this_vga_signals.M_hcounter_q_9_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11745\,
            in2 => \_gnd_net_\,
            in3 => \N__10553\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_9\,
            clk => \N__13677\,
            ce => 'H',
            sr => \N__11906\
        );

    \this_vga_signals.M_hcounter_q_10_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12224\,
            in1 => \N__11711\,
            in2 => \_gnd_net_\,
            in3 => \N__10550\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_10\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_9\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_10\,
            clk => \N__13677\,
            ce => 'H',
            sr => \N__11906\
        );

    \this_vga_signals.M_hcounter_q_11_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12223\,
            in1 => \N__12489\,
            in2 => \_gnd_net_\,
            in3 => \N__10547\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13677\,
            ce => 'H',
            sr => \N__11906\
        );

    \this_vga_signals.M_vcounter_q_0_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__10871\,
            in1 => \N__12011\,
            in2 => \N__11935\,
            in3 => \N__12225\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_2_0_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__12111\,
            in1 => \N__11744\,
            in2 => \_gnd_net_\,
            in3 => \N__11493\,
            lcout => \this_vga_signals.M_hstate_q_ns_i_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_1_0_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__11255\,
            in1 => \N__11018\,
            in2 => \N__11714\,
            in3 => \N__11768\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_0_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__11769\,
            in1 => \N__10886\,
            in2 => \N__10877\,
            in3 => \N__12731\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_0_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000100"
        )
    port map (
            in0 => \N__12066\,
            in1 => \N__12191\,
            in2 => \N__10874\,
            in3 => \N__11770\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_0_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10870\,
            in2 => \N__12226\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_LUT4_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10844\,
            in3 => \N__10802\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_LUT4_0_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10798\,
            in2 => \_gnd_net_\,
            in3 => \N__10742\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_LUT4_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10738\,
            in2 => \_gnd_net_\,
            in3 => \N__10685\,
            lcout => \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10671\,
            in2 => \_gnd_net_\,
            in3 => \N__10640\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_4\,
            clk => \N__13685\,
            ce => 'H',
            sr => \N__11905\
        );

    \this_vga_signals.M_vcounter_q_5_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10632\,
            in2 => \_gnd_net_\,
            in3 => \N__10604\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_5\,
            clk => \N__13685\,
            ce => 'H',
            sr => \N__11905\
        );

    \this_vga_signals.M_vcounter_q_6_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10591\,
            in2 => \_gnd_net_\,
            in3 => \N__10565\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_6\,
            clk => \N__13685\,
            ce => 'H',
            sr => \N__11905\
        );

    \this_vga_signals.M_vcounter_q_7_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10963\,
            in2 => \_gnd_net_\,
            in3 => \N__10937\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_7\,
            clk => \N__13685\,
            ce => 'H',
            sr => \N__11905\
        );

    \this_vga_signals.M_vcounter_q_8_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10922\,
            in2 => \_gnd_net_\,
            in3 => \N__10889\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8\,
            clk => \N__13689\,
            ce => 'H',
            sr => \N__11904\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_0_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13017\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_8\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__13084\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_0_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13021\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_1_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_3_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__13085\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_2_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_4_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13025\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_3_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_5_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__13086\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_4_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_6_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13029\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_5_THRU_CO\,
            carryout => \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__11971\,
            in1 => \N__12017\,
            in2 => \N__11934\,
            in3 => \N__11990\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11866\,
            in2 => \_gnd_net_\,
            in3 => \N__11832\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13669\,
            ce => 'H',
            sr => \N__11907\
        );

    \this_vga_signals.M_hcounter_q_0_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13669\,
            ce => 'H',
            sr => \N__11907\
        );

    \this_vga_signals.M_hcounter_q_RNI2UC41_1_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11864\,
            in1 => \N__11845\,
            in2 => \N__11833\,
            in3 => \N__11809\,
            lcout => \this_vga_signals.N_169_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNITMFU_0_9_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__11704\,
            in1 => \_gnd_net_\,
            in2 => \N__11746\,
            in3 => \N__11486\,
            lcout => \this_vga_signals.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNID7PV_0_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__11767\,
            in1 => \N__11250\,
            in2 => \_gnd_net_\,
            in3 => \N__11014\,
            lcout => \this_vga_signals.N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNITMFU_9_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__11740\,
            in1 => \_gnd_net_\,
            in2 => \N__11713\,
            in3 => \N__11485\,
            lcout => \this_vga_signals.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_4_0_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11259\,
            in2 => \_gnd_net_\,
            in3 => \N__11022\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_3_0_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000011"
        )
    port map (
            in0 => \N__12151\,
            in1 => \N__12163\,
            in2 => \N__12734\,
            in3 => \N__12108\,
            lcout => \this_vga_signals.M_hstate_q_ns_i_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12539\,
            in1 => \N__12278\,
            in2 => \N__12491\,
            in3 => \N__12236\,
            lcout => \this_vga_signals.N_169\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIPU1C1_11_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12540\,
            in1 => \N__12485\,
            in2 => \N__12288\,
            in3 => \N__12107\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_hstate_d_0_sqmuxa_0_a2_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__12175\,
            in1 => \N__12150\,
            in2 => \N__12239\,
            in3 => \N__12235\,
            lcout => \this_vga_signals.M_hstate_d_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_1_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000010"
        )
    port map (
            in0 => \N__12187\,
            in1 => \N__12083\,
            in2 => \N__12065\,
            in3 => \N__12110\,
            lcout => \this_vga_signals.M_hstate_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hstate_q_RNO_0_1_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111110"
        )
    port map (
            in0 => \N__12176\,
            in1 => \N__12164\,
            in2 => \N__12155\,
            in3 => \N__12109\,
            lcout => \this_vga_signals.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13758\,
            in2 => \_gnd_net_\,
            in3 => \N__13733\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13760\,
            in2 => \_gnd_net_\,
            in3 => \N__12023\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__13759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12029\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13757\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_2_RNI34P11_0_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13502\,
            in1 => \N__13490\,
            in2 => \_gnd_net_\,
            in3 => \N__14156\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_4_2_RNI34P11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIG1S72_11_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__14009\,
            in1 => \_gnd_net_\,
            in2 => \N__13469\,
            in3 => \N__14406\,
            lcout => \this_vram.mem_N_2372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_0_wclke_0_a2_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14650\,
            in1 => \N__14870\,
            in2 => \N__13828\,
            in3 => \N__14802\,
            lcout => \this_vram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_22_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_2_RNI9H021_0_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14478\,
            in1 => \N__12851\,
            in2 => \_gnd_net_\,
            in3 => \N__12836\,
            lcout => \this_vram.mem_mem_8_2_RNI9H021Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_1_RNI38R11_LC_24_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14169\,
            in1 => \N__12809\,
            in2 => \_gnd_net_\,
            in3 => \N__12794\,
            lcout => \this_vram.mem_mem_5_1_RNI38RZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_1_RNI38R11_0_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12770\,
            in1 => \N__14168\,
            in2 => \_gnd_net_\,
            in3 => \N__12755\,
            lcout => \this_vram.mem_mem_5_1_RNI38R11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_6_0_wclke_0_a2_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__14800\,
            in1 => \N__14845\,
            in2 => \N__13804\,
            in3 => \N__14629\,
            lcout => \this_vram.mem_WE_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_2_RNI58R11_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14225\,
            in1 => \N__14140\,
            in2 => \_gnd_net_\,
            in3 => \N__14216\,
            lcout => \this_vram.mem_mem_5_2_RNI58RZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_2_RNI58R11_0_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14183\,
            in1 => \N__14139\,
            in2 => \_gnd_net_\,
            in3 => \N__14024\,
            lcout => \this_vram.mem_mem_5_2_RNI58R11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_7_0_wclke_0_a2_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14801\,
            in1 => \N__14846\,
            in2 => \N__13805\,
            in3 => \N__14630\,
            lcout => \this_vram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_0_RNI5H021_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13964\,
            in1 => \N__14465\,
            in2 => \_gnd_net_\,
            in3 => \N__13952\,
            lcout => \this_vram.mem_mem_8_0_RNI5HZ0Z021\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_0_RNI5H021_0_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13931\,
            in1 => \N__14466\,
            in2 => \_gnd_net_\,
            in3 => \N__13925\,
            lcout => \this_vram.mem_mem_8_0_RNI5H021Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_1_RNI7H021_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13898\,
            in1 => \N__14467\,
            in2 => \_gnd_net_\,
            in3 => \N__13892\,
            lcout => \this_vram.mem_mem_8_1_RNI7HZ0Z021\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_wclke_0_a2_1_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14697\,
            lcout => \this_vram.mem_N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_9_0_wclke_0_a2_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14699\,
            in1 => \N__14705\,
            in2 => \N__14570\,
            in3 => \N__14614\,
            lcout => \this_vram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_0_wclke_0_a2_0_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__14844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14767\,
            lcout => \this_vram.mem_N_29\,
            ltout => \this_vram.mem_N_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_0_wclke_0_a2_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14698\,
            in1 => \N__14613\,
            in2 => \N__14573\,
            in3 => \N__14566\,
            lcout => \this_vram.mem_WE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_1_RNI7H021_0_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14513\,
            in1 => \N__14479\,
            in2 => \_gnd_net_\,
            in3 => \N__14501\,
            lcout => \this_vram.mem_mem_8_1_RNI7H021Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_8_2_RNI9H021_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__14480\,
            in1 => \_gnd_net_\,
            in2 => \N__14288\,
            in3 => \N__14279\,
            lcout => \this_vram.mem_mem_8_2_RNI9HZ0Z021\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
