// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 21 2022 22:52:11

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__25733;
    wire N__25732;
    wire N__25731;
    wire N__25722;
    wire N__25721;
    wire N__25720;
    wire N__25713;
    wire N__25712;
    wire N__25711;
    wire N__25704;
    wire N__25703;
    wire N__25702;
    wire N__25695;
    wire N__25694;
    wire N__25693;
    wire N__25686;
    wire N__25685;
    wire N__25684;
    wire N__25677;
    wire N__25676;
    wire N__25675;
    wire N__25668;
    wire N__25667;
    wire N__25666;
    wire N__25659;
    wire N__25658;
    wire N__25657;
    wire N__25650;
    wire N__25649;
    wire N__25648;
    wire N__25641;
    wire N__25640;
    wire N__25639;
    wire N__25632;
    wire N__25631;
    wire N__25630;
    wire N__25623;
    wire N__25622;
    wire N__25621;
    wire N__25614;
    wire N__25613;
    wire N__25612;
    wire N__25605;
    wire N__25604;
    wire N__25603;
    wire N__25596;
    wire N__25595;
    wire N__25594;
    wire N__25587;
    wire N__25586;
    wire N__25585;
    wire N__25578;
    wire N__25577;
    wire N__25576;
    wire N__25569;
    wire N__25568;
    wire N__25567;
    wire N__25560;
    wire N__25559;
    wire N__25558;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25542;
    wire N__25541;
    wire N__25540;
    wire N__25533;
    wire N__25532;
    wire N__25531;
    wire N__25524;
    wire N__25523;
    wire N__25522;
    wire N__25515;
    wire N__25514;
    wire N__25513;
    wire N__25506;
    wire N__25505;
    wire N__25504;
    wire N__25497;
    wire N__25496;
    wire N__25495;
    wire N__25488;
    wire N__25487;
    wire N__25486;
    wire N__25479;
    wire N__25478;
    wire N__25477;
    wire N__25470;
    wire N__25469;
    wire N__25468;
    wire N__25461;
    wire N__25460;
    wire N__25459;
    wire N__25452;
    wire N__25451;
    wire N__25450;
    wire N__25443;
    wire N__25442;
    wire N__25441;
    wire N__25434;
    wire N__25433;
    wire N__25432;
    wire N__25425;
    wire N__25424;
    wire N__25423;
    wire N__25416;
    wire N__25415;
    wire N__25414;
    wire N__25407;
    wire N__25406;
    wire N__25405;
    wire N__25398;
    wire N__25397;
    wire N__25396;
    wire N__25389;
    wire N__25388;
    wire N__25387;
    wire N__25380;
    wire N__25379;
    wire N__25378;
    wire N__25371;
    wire N__25370;
    wire N__25369;
    wire N__25362;
    wire N__25361;
    wire N__25360;
    wire N__25353;
    wire N__25352;
    wire N__25351;
    wire N__25344;
    wire N__25343;
    wire N__25342;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25280;
    wire N__25277;
    wire N__25276;
    wire N__25275;
    wire N__25274;
    wire N__25265;
    wire N__25264;
    wire N__25263;
    wire N__25262;
    wire N__25261;
    wire N__25260;
    wire N__25259;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25255;
    wire N__25254;
    wire N__25253;
    wire N__25252;
    wire N__25251;
    wire N__25248;
    wire N__25239;
    wire N__25230;
    wire N__25221;
    wire N__25220;
    wire N__25219;
    wire N__25216;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25212;
    wire N__25209;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25197;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25165;
    wire N__25162;
    wire N__25161;
    wire N__25160;
    wire N__25159;
    wire N__25156;
    wire N__25155;
    wire N__25154;
    wire N__25153;
    wire N__25152;
    wire N__25147;
    wire N__25144;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25097;
    wire N__25092;
    wire N__25089;
    wire N__25082;
    wire N__25079;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25037;
    wire N__25036;
    wire N__25035;
    wire N__25034;
    wire N__25033;
    wire N__25032;
    wire N__25031;
    wire N__25030;
    wire N__25029;
    wire N__25028;
    wire N__25027;
    wire N__25026;
    wire N__25025;
    wire N__25024;
    wire N__25023;
    wire N__25022;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25017;
    wire N__25016;
    wire N__25015;
    wire N__25014;
    wire N__25013;
    wire N__25012;
    wire N__25011;
    wire N__25010;
    wire N__25009;
    wire N__25008;
    wire N__25007;
    wire N__25006;
    wire N__25005;
    wire N__25004;
    wire N__25003;
    wire N__25002;
    wire N__25001;
    wire N__25000;
    wire N__24999;
    wire N__24998;
    wire N__24997;
    wire N__24996;
    wire N__24995;
    wire N__24994;
    wire N__24993;
    wire N__24992;
    wire N__24991;
    wire N__24990;
    wire N__24989;
    wire N__24988;
    wire N__24987;
    wire N__24986;
    wire N__24985;
    wire N__24984;
    wire N__24983;
    wire N__24982;
    wire N__24981;
    wire N__24980;
    wire N__24979;
    wire N__24978;
    wire N__24977;
    wire N__24976;
    wire N__24975;
    wire N__24974;
    wire N__24973;
    wire N__24972;
    wire N__24971;
    wire N__24970;
    wire N__24969;
    wire N__24968;
    wire N__24967;
    wire N__24966;
    wire N__24965;
    wire N__24964;
    wire N__24963;
    wire N__24962;
    wire N__24961;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24799;
    wire N__24798;
    wire N__24795;
    wire N__24794;
    wire N__24793;
    wire N__24792;
    wire N__24791;
    wire N__24790;
    wire N__24789;
    wire N__24788;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24770;
    wire N__24765;
    wire N__24762;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24746;
    wire N__24745;
    wire N__24744;
    wire N__24743;
    wire N__24742;
    wire N__24741;
    wire N__24740;
    wire N__24739;
    wire N__24738;
    wire N__24737;
    wire N__24736;
    wire N__24735;
    wire N__24734;
    wire N__24733;
    wire N__24732;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24362;
    wire N__24359;
    wire N__24358;
    wire N__24355;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24321;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24302;
    wire N__24299;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24281;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24265;
    wire N__24262;
    wire N__24257;
    wire N__24254;
    wire N__24249;
    wire N__24248;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24230;
    wire N__24227;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24209;
    wire N__24208;
    wire N__24207;
    wire N__24206;
    wire N__24203;
    wire N__24198;
    wire N__24195;
    wire N__24194;
    wire N__24191;
    wire N__24186;
    wire N__24183;
    wire N__24176;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24164;
    wire N__24161;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24149;
    wire N__24146;
    wire N__24141;
    wire N__24134;
    wire N__24131;
    wire N__24130;
    wire N__24129;
    wire N__24124;
    wire N__24121;
    wire N__24120;
    wire N__24115;
    wire N__24112;
    wire N__24107;
    wire N__24104;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24096;
    wire N__24095;
    wire N__24094;
    wire N__24089;
    wire N__24084;
    wire N__24081;
    wire N__24080;
    wire N__24079;
    wire N__24076;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24056;
    wire N__24055;
    wire N__24054;
    wire N__24053;
    wire N__24052;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24034;
    wire N__24031;
    wire N__24030;
    wire N__24027;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23989;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23950;
    wire N__23947;
    wire N__23942;
    wire N__23941;
    wire N__23940;
    wire N__23935;
    wire N__23932;
    wire N__23931;
    wire N__23930;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23919;
    wire N__23918;
    wire N__23913;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23892;
    wire N__23889;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23860;
    wire N__23859;
    wire N__23858;
    wire N__23857;
    wire N__23856;
    wire N__23855;
    wire N__23854;
    wire N__23853;
    wire N__23852;
    wire N__23851;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23843;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23831;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23823;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23760;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23739;
    wire N__23736;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23718;
    wire N__23709;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23692;
    wire N__23691;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23548;
    wire N__23547;
    wire N__23546;
    wire N__23545;
    wire N__23544;
    wire N__23543;
    wire N__23542;
    wire N__23541;
    wire N__23540;
    wire N__23537;
    wire N__23536;
    wire N__23535;
    wire N__23534;
    wire N__23531;
    wire N__23530;
    wire N__23527;
    wire N__23526;
    wire N__23523;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23505;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23474;
    wire N__23471;
    wire N__23470;
    wire N__23467;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23431;
    wire N__23430;
    wire N__23425;
    wire N__23422;
    wire N__23415;
    wire N__23408;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23198;
    wire N__23195;
    wire N__23194;
    wire N__23193;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23107;
    wire N__23104;
    wire N__23103;
    wire N__23100;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23085;
    wire N__23080;
    wire N__23077;
    wire N__23076;
    wire N__23071;
    wire N__23068;
    wire N__23067;
    wire N__23062;
    wire N__23059;
    wire N__23054;
    wire N__23051;
    wire N__23046;
    wire N__23041;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22914;
    wire N__22911;
    wire N__22910;
    wire N__22909;
    wire N__22908;
    wire N__22907;
    wire N__22906;
    wire N__22905;
    wire N__22904;
    wire N__22899;
    wire N__22898;
    wire N__22897;
    wire N__22896;
    wire N__22895;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22883;
    wire N__22880;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22855;
    wire N__22850;
    wire N__22841;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22819;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22788;
    wire N__22783;
    wire N__22780;
    wire N__22779;
    wire N__22774;
    wire N__22771;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22759;
    wire N__22756;
    wire N__22755;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22740;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22712;
    wire N__22711;
    wire N__22708;
    wire N__22703;
    wire N__22700;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22664;
    wire N__22661;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22387;
    wire N__22386;
    wire N__22385;
    wire N__22384;
    wire N__22379;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22365;
    wire N__22364;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22341;
    wire N__22338;
    wire N__22331;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22300;
    wire N__22299;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22265;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22238;
    wire N__22233;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22217;
    wire N__22214;
    wire N__22213;
    wire N__22212;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22165;
    wire N__22162;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22055;
    wire N__22054;
    wire N__22053;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22045;
    wire N__22044;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22040;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22032;
    wire N__22031;
    wire N__22030;
    wire N__22029;
    wire N__22028;
    wire N__22027;
    wire N__22026;
    wire N__22023;
    wire N__22022;
    wire N__22021;
    wire N__22018;
    wire N__22011;
    wire N__22004;
    wire N__22003;
    wire N__22000;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21978;
    wire N__21977;
    wire N__21976;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21956;
    wire N__21953;
    wire N__21948;
    wire N__21939;
    wire N__21936;
    wire N__21929;
    wire N__21922;
    wire N__21917;
    wire N__21912;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21890;
    wire N__21887;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21661;
    wire N__21660;
    wire N__21653;
    wire N__21650;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21638;
    wire N__21637;
    wire N__21636;
    wire N__21635;
    wire N__21634;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21626;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21602;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21587;
    wire N__21584;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21572;
    wire N__21567;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21542;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21517;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21280;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21232;
    wire N__21231;
    wire N__21226;
    wire N__21225;
    wire N__21224;
    wire N__21223;
    wire N__21220;
    wire N__21219;
    wire N__21216;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21212;
    wire N__21207;
    wire N__21204;
    wire N__21199;
    wire N__21198;
    wire N__21197;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21183;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21171;
    wire N__21170;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21155;
    wire N__21152;
    wire N__21147;
    wire N__21142;
    wire N__21139;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21115;
    wire N__21114;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21092;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21078;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21047;
    wire N__21044;
    wire N__21043;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20972;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20956;
    wire N__20953;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20927;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20902;
    wire N__20899;
    wire N__20894;
    wire N__20887;
    wire N__20882;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20874;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20850;
    wire N__20847;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20831;
    wire N__20828;
    wire N__20827;
    wire N__20824;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20789;
    wire N__20786;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20778;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20767;
    wire N__20764;
    wire N__20763;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20745;
    wire N__20744;
    wire N__20739;
    wire N__20736;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20630;
    wire N__20627;
    wire N__20626;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20611;
    wire N__20608;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20590;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20544;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20532;
    wire N__20529;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20506;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20491;
    wire N__20488;
    wire N__20487;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20462;
    wire N__20459;
    wire N__20458;
    wire N__20453;
    wire N__20450;
    wire N__20449;
    wire N__20448;
    wire N__20447;
    wire N__20446;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20428;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20245;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20218;
    wire N__20215;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20167;
    wire N__20162;
    wire N__20157;
    wire N__20154;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19861;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19843;
    wire N__19840;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19821;
    wire N__19816;
    wire N__19813;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19801;
    wire N__19800;
    wire N__19799;
    wire N__19798;
    wire N__19795;
    wire N__19794;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19778;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19756;
    wire N__19755;
    wire N__19754;
    wire N__19751;
    wire N__19746;
    wire N__19743;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19571;
    wire N__19568;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19556;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19544;
    wire N__19541;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19514;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19499;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19487;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19475;
    wire N__19472;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19460;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19442;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19430;
    wire N__19427;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19415;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19403;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19388;
    wire N__19385;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19351;
    wire N__19346;
    wire N__19345;
    wire N__19344;
    wire N__19341;
    wire N__19336;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19216;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19077;
    wire N__19074;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18784;
    wire N__18781;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18759;
    wire N__18758;
    wire N__18753;
    wire N__18750;
    wire N__18749;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18741;
    wire N__18740;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18716;
    wire N__18715;
    wire N__18714;
    wire N__18711;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18653;
    wire N__18650;
    wire N__18643;
    wire N__18642;
    wire N__18639;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18585;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18472;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18346;
    wire N__18343;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18328;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18286;
    wire N__18285;
    wire N__18282;
    wire N__18277;
    wire N__18272;
    wire N__18269;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18250;
    wire N__18249;
    wire N__18248;
    wire N__18247;
    wire N__18246;
    wire N__18245;
    wire N__18244;
    wire N__18241;
    wire N__18232;
    wire N__18229;
    wire N__18224;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18106;
    wire N__18105;
    wire N__18102;
    wire N__18101;
    wire N__18100;
    wire N__18099;
    wire N__18098;
    wire N__18097;
    wire N__18094;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18083;
    wire N__18082;
    wire N__18079;
    wire N__18076;
    wire N__18071;
    wire N__18068;
    wire N__18067;
    wire N__18066;
    wire N__18063;
    wire N__18062;
    wire N__18057;
    wire N__18054;
    wire N__18049;
    wire N__18046;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18013;
    wire N__17996;
    wire N__17995;
    wire N__17994;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17979;
    wire N__17974;
    wire N__17971;
    wire N__17966;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17954;
    wire N__17953;
    wire N__17952;
    wire N__17951;
    wire N__17946;
    wire N__17941;
    wire N__17936;
    wire N__17935;
    wire N__17934;
    wire N__17933;
    wire N__17930;
    wire N__17929;
    wire N__17928;
    wire N__17927;
    wire N__17920;
    wire N__17917;
    wire N__17910;
    wire N__17903;
    wire N__17902;
    wire N__17901;
    wire N__17898;
    wire N__17897;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17889;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17871;
    wire N__17870;
    wire N__17869;
    wire N__17866;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17839;
    wire N__17832;
    wire N__17829;
    wire N__17820;
    wire N__17807;
    wire N__17804;
    wire N__17803;
    wire N__17802;
    wire N__17801;
    wire N__17800;
    wire N__17799;
    wire N__17796;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17775;
    wire N__17774;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17751;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17735;
    wire N__17728;
    wire N__17717;
    wire N__17714;
    wire N__17713;
    wire N__17712;
    wire N__17709;
    wire N__17704;
    wire N__17699;
    wire N__17696;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17675;
    wire N__17674;
    wire N__17673;
    wire N__17672;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17661;
    wire N__17660;
    wire N__17659;
    wire N__17658;
    wire N__17655;
    wire N__17652;
    wire N__17649;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17637;
    wire N__17636;
    wire N__17635;
    wire N__17632;
    wire N__17631;
    wire N__17630;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17604;
    wire N__17603;
    wire N__17602;
    wire N__17599;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17591;
    wire N__17590;
    wire N__17589;
    wire N__17586;
    wire N__17585;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17560;
    wire N__17559;
    wire N__17556;
    wire N__17553;
    wire N__17550;
    wire N__17549;
    wire N__17544;
    wire N__17541;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17523;
    wire N__17522;
    wire N__17519;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17503;
    wire N__17502;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17492;
    wire N__17489;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17458;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17435;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17423;
    wire N__17416;
    wire N__17409;
    wire N__17406;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17379;
    wire N__17372;
    wire N__17369;
    wire N__17364;
    wire N__17361;
    wire N__17354;
    wire N__17349;
    wire N__17348;
    wire N__17347;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17329;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17273;
    wire N__17272;
    wire N__17267;
    wire N__17264;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17200;
    wire N__17195;
    wire N__17194;
    wire N__17191;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17179;
    wire N__17174;
    wire N__17173;
    wire N__17172;
    wire N__17171;
    wire N__17170;
    wire N__17165;
    wire N__17160;
    wire N__17157;
    wire N__17150;
    wire N__17149;
    wire N__17148;
    wire N__17147;
    wire N__17146;
    wire N__17145;
    wire N__17144;
    wire N__17143;
    wire N__17142;
    wire N__17141;
    wire N__17140;
    wire N__17133;
    wire N__17128;
    wire N__17123;
    wire N__17120;
    wire N__17119;
    wire N__17118;
    wire N__17111;
    wire N__17108;
    wire N__17103;
    wire N__17100;
    wire N__17095;
    wire N__17092;
    wire N__17087;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17057;
    wire N__17056;
    wire N__17055;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17029;
    wire N__17026;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17006;
    wire N__17003;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16997;
    wire N__16996;
    wire N__16993;
    wire N__16992;
    wire N__16989;
    wire N__16988;
    wire N__16987;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16974;
    wire N__16971;
    wire N__16968;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16956;
    wire N__16955;
    wire N__16948;
    wire N__16943;
    wire N__16940;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16888;
    wire N__16887;
    wire N__16884;
    wire N__16879;
    wire N__16874;
    wire N__16871;
    wire N__16870;
    wire N__16869;
    wire N__16868;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16853;
    wire N__16850;
    wire N__16845;
    wire N__16842;
    wire N__16835;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16816;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16774;
    wire N__16773;
    wire N__16770;
    wire N__16765;
    wire N__16764;
    wire N__16763;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16748;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16726;
    wire N__16725;
    wire N__16722;
    wire N__16717;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16700;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16662;
    wire N__16661;
    wire N__16656;
    wire N__16651;
    wire N__16646;
    wire N__16643;
    wire N__16642;
    wire N__16641;
    wire N__16640;
    wire N__16639;
    wire N__16638;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16616;
    wire N__16615;
    wire N__16614;
    wire N__16613;
    wire N__16612;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16592;
    wire N__16589;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16562;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16544;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16342;
    wire N__16339;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16319;
    wire N__16318;
    wire N__16317;
    wire N__16316;
    wire N__16315;
    wire N__16314;
    wire N__16311;
    wire N__16310;
    wire N__16309;
    wire N__16304;
    wire N__16301;
    wire N__16292;
    wire N__16291;
    wire N__16290;
    wire N__16287;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16268;
    wire N__16257;
    wire N__16254;
    wire N__16241;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16233;
    wire N__16230;
    wire N__16225;
    wire N__16220;
    wire N__16217;
    wire N__16216;
    wire N__16215;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16207;
    wire N__16206;
    wire N__16205;
    wire N__16204;
    wire N__16203;
    wire N__16202;
    wire N__16199;
    wire N__16198;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16172;
    wire N__16171;
    wire N__16170;
    wire N__16169;
    wire N__16168;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16148;
    wire N__16141;
    wire N__16130;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16102;
    wire N__16101;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16093;
    wire N__16092;
    wire N__16089;
    wire N__16086;
    wire N__16085;
    wire N__16082;
    wire N__16077;
    wire N__16074;
    wire N__16069;
    wire N__16066;
    wire N__16065;
    wire N__16064;
    wire N__16063;
    wire N__16062;
    wire N__16057;
    wire N__16056;
    wire N__16053;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16023;
    wire N__16018;
    wire N__16007;
    wire N__16004;
    wire N__16003;
    wire N__16002;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15992;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15984;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15976;
    wire N__15973;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15961;
    wire N__15960;
    wire N__15959;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15943;
    wire N__15940;
    wire N__15939;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15924;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15889;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15878;
    wire N__15877;
    wire N__15876;
    wire N__15875;
    wire N__15870;
    wire N__15867;
    wire N__15864;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15854;
    wire N__15847;
    wire N__15846;
    wire N__15845;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15806;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15794;
    wire N__15793;
    wire N__15792;
    wire N__15791;
    wire N__15790;
    wire N__15785;
    wire N__15782;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15774;
    wire N__15769;
    wire N__15768;
    wire N__15767;
    wire N__15766;
    wire N__15765;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15731;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15707;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15686;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15661;
    wire N__15658;
    wire N__15657;
    wire N__15654;
    wire N__15651;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15623;
    wire N__15622;
    wire N__15621;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15613;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15552;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15529;
    wire N__15524;
    wire N__15523;
    wire N__15522;
    wire N__15521;
    wire N__15520;
    wire N__15519;
    wire N__15518;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15493;
    wire N__15492;
    wire N__15491;
    wire N__15490;
    wire N__15489;
    wire N__15488;
    wire N__15487;
    wire N__15486;
    wire N__15483;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15451;
    wire N__15450;
    wire N__15449;
    wire N__15448;
    wire N__15447;
    wire N__15446;
    wire N__15443;
    wire N__15442;
    wire N__15441;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15433;
    wire N__15432;
    wire N__15431;
    wire N__15430;
    wire N__15429;
    wire N__15428;
    wire N__15427;
    wire N__15426;
    wire N__15425;
    wire N__15424;
    wire N__15423;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15415;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15403;
    wire N__15402;
    wire N__15399;
    wire N__15398;
    wire N__15397;
    wire N__15394;
    wire N__15389;
    wire N__15384;
    wire N__15381;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15362;
    wire N__15359;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15340;
    wire N__15339;
    wire N__15334;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15315;
    wire N__15308;
    wire N__15301;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15285;
    wire N__15280;
    wire N__15277;
    wire N__15272;
    wire N__15265;
    wire N__15264;
    wire N__15261;
    wire N__15256;
    wire N__15251;
    wire N__15244;
    wire N__15237;
    wire N__15236;
    wire N__15233;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15203;
    wire N__15202;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15155;
    wire N__15154;
    wire N__15153;
    wire N__15152;
    wire N__15151;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15143;
    wire N__15142;
    wire N__15141;
    wire N__15138;
    wire N__15137;
    wire N__15136;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15128;
    wire N__15127;
    wire N__15126;
    wire N__15125;
    wire N__15122;
    wire N__15119;
    wire N__15110;
    wire N__15107;
    wire N__15106;
    wire N__15105;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15094;
    wire N__15093;
    wire N__15092;
    wire N__15087;
    wire N__15084;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15064;
    wire N__15063;
    wire N__15060;
    wire N__15053;
    wire N__15050;
    wire N__15045;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15030;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15018;
    wire N__15011;
    wire N__15006;
    wire N__14997;
    wire N__14994;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14908;
    wire N__14907;
    wire N__14904;
    wire N__14899;
    wire N__14894;
    wire N__14891;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14863;
    wire N__14862;
    wire N__14859;
    wire N__14854;
    wire N__14849;
    wire N__14846;
    wire N__14845;
    wire N__14844;
    wire N__14843;
    wire N__14840;
    wire N__14833;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14803;
    wire N__14802;
    wire N__14801;
    wire N__14794;
    wire N__14791;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14716;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14686;
    wire N__14685;
    wire N__14682;
    wire N__14677;
    wire N__14672;
    wire N__14671;
    wire N__14670;
    wire N__14665;
    wire N__14662;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14581;
    wire N__14580;
    wire N__14579;
    wire N__14578;
    wire N__14577;
    wire N__14576;
    wire N__14575;
    wire N__14574;
    wire N__14573;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14565;
    wire N__14564;
    wire N__14563;
    wire N__14562;
    wire N__14561;
    wire N__14558;
    wire N__14557;
    wire N__14556;
    wire N__14555;
    wire N__14552;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14541;
    wire N__14540;
    wire N__14535;
    wire N__14532;
    wire N__14531;
    wire N__14526;
    wire N__14519;
    wire N__14514;
    wire N__14513;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14499;
    wire N__14498;
    wire N__14495;
    wire N__14488;
    wire N__14483;
    wire N__14480;
    wire N__14475;
    wire N__14472;
    wire N__14471;
    wire N__14470;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14454;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14420;
    wire N__14415;
    wire N__14410;
    wire N__14403;
    wire N__14400;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14384;
    wire N__14383;
    wire N__14380;
    wire N__14379;
    wire N__14378;
    wire N__14377;
    wire N__14376;
    wire N__14375;
    wire N__14374;
    wire N__14373;
    wire N__14372;
    wire N__14371;
    wire N__14370;
    wire N__14369;
    wire N__14368;
    wire N__14367;
    wire N__14366;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14351;
    wire N__14348;
    wire N__14347;
    wire N__14346;
    wire N__14345;
    wire N__14344;
    wire N__14343;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14335;
    wire N__14334;
    wire N__14333;
    wire N__14330;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14312;
    wire N__14307;
    wire N__14306;
    wire N__14305;
    wire N__14304;
    wire N__14303;
    wire N__14302;
    wire N__14301;
    wire N__14296;
    wire N__14291;
    wire N__14284;
    wire N__14281;
    wire N__14276;
    wire N__14271;
    wire N__14270;
    wire N__14267;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14255;
    wire N__14254;
    wire N__14251;
    wire N__14242;
    wire N__14237;
    wire N__14234;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14214;
    wire N__14207;
    wire N__14204;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14180;
    wire N__14173;
    wire N__14164;
    wire N__14157;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14131;
    wire N__14130;
    wire N__14129;
    wire N__14128;
    wire N__14127;
    wire N__14126;
    wire N__14123;
    wire N__14122;
    wire N__14119;
    wire N__14118;
    wire N__14115;
    wire N__14114;
    wire N__14113;
    wire N__14110;
    wire N__14109;
    wire N__14108;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14075;
    wire N__14068;
    wire N__14067;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14022;
    wire N__14017;
    wire N__14014;
    wire N__14007;
    wire N__14004;
    wire N__13991;
    wire N__13988;
    wire N__13987;
    wire N__13986;
    wire N__13985;
    wire N__13982;
    wire N__13981;
    wire N__13978;
    wire N__13977;
    wire N__13974;
    wire N__13967;
    wire N__13966;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13943;
    wire N__13938;
    wire N__13931;
    wire N__13930;
    wire N__13929;
    wire N__13928;
    wire N__13927;
    wire N__13926;
    wire N__13925;
    wire N__13924;
    wire N__13923;
    wire N__13920;
    wire N__13913;
    wire N__13912;
    wire N__13911;
    wire N__13908;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13892;
    wire N__13887;
    wire N__13886;
    wire N__13885;
    wire N__13884;
    wire N__13881;
    wire N__13874;
    wire N__13869;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13804;
    wire N__13803;
    wire N__13802;
    wire N__13801;
    wire N__13800;
    wire N__13799;
    wire N__13798;
    wire N__13797;
    wire N__13794;
    wire N__13793;
    wire N__13792;
    wire N__13791;
    wire N__13790;
    wire N__13789;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13777;
    wire N__13774;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13751;
    wire N__13746;
    wire N__13743;
    wire N__13736;
    wire N__13733;
    wire N__13728;
    wire N__13723;
    wire N__13706;
    wire N__13705;
    wire N__13702;
    wire N__13701;
    wire N__13700;
    wire N__13699;
    wire N__13698;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13683;
    wire N__13678;
    wire N__13677;
    wire N__13676;
    wire N__13675;
    wire N__13674;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13657;
    wire N__13656;
    wire N__13655;
    wire N__13652;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13642;
    wire N__13637;
    wire N__13634;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13601;
    wire N__13586;
    wire N__13585;
    wire N__13584;
    wire N__13583;
    wire N__13582;
    wire N__13579;
    wire N__13578;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13568;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13558;
    wire N__13557;
    wire N__13556;
    wire N__13555;
    wire N__13554;
    wire N__13551;
    wire N__13546;
    wire N__13545;
    wire N__13544;
    wire N__13539;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13523;
    wire N__13520;
    wire N__13515;
    wire N__13510;
    wire N__13507;
    wire N__13490;
    wire N__13487;
    wire N__13486;
    wire N__13485;
    wire N__13482;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13458;
    wire N__13453;
    wire N__13450;
    wire N__13447;
    wire N__13444;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13402;
    wire N__13399;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13369;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13359;
    wire N__13358;
    wire N__13355;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13331;
    wire N__13322;
    wire N__13321;
    wire N__13318;
    wire N__13317;
    wire N__13316;
    wire N__13315;
    wire N__13314;
    wire N__13311;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13297;
    wire N__13294;
    wire N__13293;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13250;
    wire N__13245;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13207;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13174;
    wire N__13173;
    wire N__13170;
    wire N__13165;
    wire N__13160;
    wire N__13159;
    wire N__13156;
    wire N__13155;
    wire N__13154;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13146;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13131;
    wire N__13128;
    wire N__13119;
    wire N__13112;
    wire N__13111;
    wire N__13108;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13085;
    wire N__13082;
    wire N__13081;
    wire N__13080;
    wire N__13077;
    wire N__13072;
    wire N__13067;
    wire N__13066;
    wire N__13065;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13049;
    wire N__13046;
    wire N__13045;
    wire N__13042;
    wire N__13039;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13022;
    wire N__13021;
    wire N__13020;
    wire N__13019;
    wire N__13018;
    wire N__13017;
    wire N__13016;
    wire N__13011;
    wire N__13000;
    wire N__12999;
    wire N__12994;
    wire N__12993;
    wire N__12992;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12977;
    wire N__12968;
    wire N__12967;
    wire N__12962;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12947;
    wire N__12944;
    wire N__12943;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12901;
    wire N__12898;
    wire N__12895;
    wire N__12890;
    wire N__12887;
    wire N__12886;
    wire N__12881;
    wire N__12878;
    wire N__12877;
    wire N__12874;
    wire N__12871;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12856;
    wire N__12853;
    wire N__12852;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12840;
    wire N__12833;
    wire N__12830;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12818;
    wire N__12817;
    wire N__12816;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12774;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12724;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12706;
    wire N__12705;
    wire N__12704;
    wire N__12699;
    wire N__12694;
    wire N__12687;
    wire N__12680;
    wire N__12679;
    wire N__12674;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12662;
    wire N__12661;
    wire N__12660;
    wire N__12657;
    wire N__12652;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12640;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12632;
    wire N__12631;
    wire N__12630;
    wire N__12629;
    wire N__12628;
    wire N__12625;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12568;
    wire N__12567;
    wire N__12562;
    wire N__12561;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12553;
    wire N__12552;
    wire N__12551;
    wire N__12550;
    wire N__12549;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12538;
    wire N__12537;
    wire N__12536;
    wire N__12535;
    wire N__12534;
    wire N__12533;
    wire N__12532;
    wire N__12529;
    wire N__12522;
    wire N__12515;
    wire N__12510;
    wire N__12507;
    wire N__12498;
    wire N__12491;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12466;
    wire N__12461;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12453;
    wire N__12448;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12406;
    wire N__12405;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12376;
    wire N__12375;
    wire N__12374;
    wire N__12373;
    wire N__12372;
    wire N__12369;
    wire N__12368;
    wire N__12367;
    wire N__12366;
    wire N__12365;
    wire N__12364;
    wire N__12363;
    wire N__12362;
    wire N__12361;
    wire N__12358;
    wire N__12357;
    wire N__12348;
    wire N__12345;
    wire N__12340;
    wire N__12337;
    wire N__12330;
    wire N__12323;
    wire N__12320;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12287;
    wire N__12284;
    wire N__12281;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12269;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12235;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12199;
    wire N__12198;
    wire N__12195;
    wire N__12194;
    wire N__12193;
    wire N__12192;
    wire N__12191;
    wire N__12190;
    wire N__12189;
    wire N__12184;
    wire N__12181;
    wire N__12176;
    wire N__12175;
    wire N__12174;
    wire N__12173;
    wire N__12172;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12164;
    wire N__12161;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12145;
    wire N__12140;
    wire N__12137;
    wire N__12126;
    wire N__12117;
    wire N__12114;
    wire N__12095;
    wire N__12092;
    wire N__12091;
    wire N__12090;
    wire N__12089;
    wire N__12088;
    wire N__12085;
    wire N__12084;
    wire N__12083;
    wire N__12082;
    wire N__12079;
    wire N__12074;
    wire N__12073;
    wire N__12072;
    wire N__12071;
    wire N__12070;
    wire N__12069;
    wire N__12068;
    wire N__12067;
    wire N__12066;
    wire N__12065;
    wire N__12062;
    wire N__12061;
    wire N__12058;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12036;
    wire N__12029;
    wire N__12020;
    wire N__12017;
    wire N__11996;
    wire N__11995;
    wire N__11992;
    wire N__11989;
    wire N__11986;
    wire N__11983;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11956;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11950;
    wire N__11943;
    wire N__11940;
    wire N__11933;
    wire N__11930;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11918;
    wire N__11917;
    wire N__11916;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11900;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11888;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11880;
    wire N__11879;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11861;
    wire N__11858;
    wire N__11857;
    wire N__11854;
    wire N__11853;
    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11845;
    wire N__11844;
    wire N__11841;
    wire N__11836;
    wire N__11835;
    wire N__11832;
    wire N__11831;
    wire N__11830;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11806;
    wire N__11803;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11767;
    wire N__11764;
    wire N__11761;
    wire N__11756;
    wire N__11755;
    wire N__11754;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11728;
    wire N__11727;
    wire N__11726;
    wire N__11725;
    wire N__11716;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11699;
    wire N__11698;
    wire N__11697;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11685;
    wire N__11680;
    wire N__11675;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11620;
    wire N__11617;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11592;
    wire N__11585;
    wire N__11580;
    wire N__11573;
    wire N__11570;
    wire N__11569;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11543;
    wire N__11540;
    wire N__11539;
    wire N__11538;
    wire N__11535;
    wire N__11530;
    wire N__11525;
    wire N__11524;
    wire N__11521;
    wire N__11520;
    wire N__11517;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11464;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11443;
    wire N__11440;
    wire N__11439;
    wire N__11436;
    wire N__11435;
    wire N__11432;
    wire N__11425;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11398;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11381;
    wire N__11380;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11329;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11300;
    wire N__11291;
    wire N__11288;
    wire N__11287;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11283;
    wire N__11280;
    wire N__11279;
    wire N__11278;
    wire N__11277;
    wire N__11276;
    wire N__11275;
    wire N__11274;
    wire N__11273;
    wire N__11272;
    wire N__11271;
    wire N__11266;
    wire N__11263;
    wire N__11258;
    wire N__11249;
    wire N__11244;
    wire N__11235;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11200;
    wire N__11195;
    wire N__11194;
    wire N__11193;
    wire N__11190;
    wire N__11185;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10977;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10842;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10587;
    wire N__10580;
    wire N__10577;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10535;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10523;
    wire N__10520;
    wire N__10519;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10504;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10492;
    wire N__10491;
    wire N__10486;
    wire N__10483;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10365;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10347;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10224;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10056;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9936;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9851;
    wire N__9848;
    wire N__9847;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9803;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9788;
    wire N__9785;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9653;
    wire N__9650;
    wire N__9649;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9505;
    wire N__9504;
    wire N__9501;
    wire N__9496;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9475;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9394;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9301;
    wire N__9300;
    wire N__9295;
    wire N__9292;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9271;
    wire N__9266;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9223;
    wire N__9222;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9177;
    wire N__9172;
    wire N__9169;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9145;
    wire N__9144;
    wire N__9141;
    wire N__9136;
    wire N__9131;
    wire N__9130;
    wire N__9129;
    wire N__9126;
    wire N__9121;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9079;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8905;
    wire N__8904;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8892;
    wire N__8891;
    wire N__8890;
    wire N__8885;
    wire N__8882;
    wire N__8877;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8863;
    wire N__8862;
    wire N__8861;
    wire N__8856;
    wire N__8851;
    wire N__8850;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8838;
    wire N__8835;
    wire N__8830;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8808;
    wire N__8805;
    wire N__8800;
    wire N__8795;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8779;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8763;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8744;
    wire N__8743;
    wire N__8740;
    wire N__8735;
    wire N__8732;
    wire N__8727;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8707;
    wire N__8706;
    wire N__8705;
    wire N__8704;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8690;
    wire N__8687;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire VCCG0;
    wire \this_vga_signals.N_517_1 ;
    wire N_205_i;
    wire \this_vga_ramdac.M_this_rgb_d_3_0_dreg ;
    wire \this_vga_ramdac.m5_cascade_ ;
    wire \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_0 ;
    wire \this_vga_ramdac.m16 ;
    wire \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_2 ;
    wire \this_vga_ramdac.m19 ;
    wire \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_3 ;
    wire \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_1 ;
    wire \this_vga_ramdac.i2_mux ;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_1;
    wire M_this_vram_read_data_3;
    wire \this_vga_ramdac.N_706_0 ;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire \this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_4 ;
    wire N_94;
    wire N_274_i;
    wire \this_vga_signals.if_N_6_mux_0_0_cascade_ ;
    wire M_this_vga_signals_address_8;
    wire M_this_vga_signals_address_11;
    wire \this_vga_signals.g0_0_a2_1 ;
    wire M_this_vga_signals_address_9;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1 ;
    wire \this_vga_signals.g2_0_x1 ;
    wire \this_vga_signals.g2_0_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0 ;
    wire \this_vga_signals.g2_0 ;
    wire M_this_vga_signals_address_12;
    wire \this_vga_signals.g0_2 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_1 ;
    wire bfn_9_12_0_;
    wire \this_vga_signals.mult1_un40_sum_cry_0 ;
    wire \this_vga_signals.mult1_un40_sum_cry_1 ;
    wire \this_vga_signals.mult1_un40_sum_cry_2 ;
    wire N_70_cascade_;
    wire \this_vga_signals.mult1_un40_sum_cry_1_THRU_CO ;
    wire G_501;
    wire N_70;
    wire N_26;
    wire bfn_9_14_0_;
    wire \this_vga_signals.mult1_un47_sum_cry_0 ;
    wire \this_vga_signals.mult1_un40_sum_cry_1_s ;
    wire \this_vga_signals.mult1_un47_sum_cry_1 ;
    wire \this_vga_signals.mult1_un47_sum_axb_3 ;
    wire \this_vga_signals.mult1_un47_sum_cry_2 ;
    wire \this_vga_signals.mult1_un40_sum_axb_2 ;
    wire \this_vga_signals.mult1_un40_sum_axb_1_l_fx ;
    wire \this_vga_signals.mult1_un40_sum_cry_2_THRU_CO ;
    wire \this_vga_signals.mult1_un40_sum_s_3 ;
    wire bfn_9_15_0_;
    wire \this_vga_signals.mult1_un61_sum_cry_0 ;
    wire \this_vga_signals.mult1_un61_sum_cry_1 ;
    wire \this_vga_signals.mult1_un61_sum_cry_2 ;
    wire \this_vga_signals.N_70_0 ;
    wire \this_vga_signals.mult1_un54_sum_i_3 ;
    wire bfn_9_16_0_;
    wire \this_vga_signals.mult1_un54_sum_cry_1_s ;
    wire \this_vga_signals.mult1_un54_sum_cry_0 ;
    wire \this_vga_signals.mult1_un47_sum_cry_1_s ;
    wire \this_vga_signals.mult1_un61_sum_axb_3 ;
    wire \this_vga_signals.mult1_un54_sum_cry_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb_3 ;
    wire \this_vga_signals.mult1_un54_sum_cry_2 ;
    wire \this_vga_signals.mult1_un54_sum_s_3 ;
    wire \this_vga_signals.M_hcounter_q_i_0_5 ;
    wire \this_vga_signals.mult1_un47_sum_s_3 ;
    wire \this_vga_signals.mult1_un47_sum_i_3 ;
    wire \this_ppu.M_N_6_0_cascade_ ;
    wire \this_ppu.M_N_13_mux ;
    wire \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_0 ;
    wire \this_ppu.M_N_15_mux_cascade_ ;
    wire \this_ppu.M_m12_0_x3_s_0_1Z0Z_0_cascade_ ;
    wire \this_ppu.M_m12_0_x3_out_0_cascade_ ;
    wire \this_vga_signals.if_m12_cascade_ ;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0_cascade_;
    wire \this_ppu.N_277 ;
    wire \this_ppu.M_mZ0Z1_cascade_ ;
    wire N_92;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_cascade_;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1;
    wire \this_ppu.M_N_16_1_cascade_ ;
    wire \this_ppu.M_m9_i_x3Z0Z_0 ;
    wire \this_ppu.M_mZ0Z1 ;
    wire \this_ppu.M_m1_e_0_1_0_cascade_ ;
    wire \this_ppu.M_m1_e_0_1_1 ;
    wire \this_ppu.M_m12_0_x3_out_0 ;
    wire \this_ppu.M_N_16_1 ;
    wire \this_ppu.M_m1_e_0_0 ;
    wire bfn_9_20_0_;
    wire \this_ppu.un1_M_current_q_cry_0 ;
    wire \this_ppu.un1_M_current_q_cry_1 ;
    wire \this_ppu.un1_M_current_q_cry_2 ;
    wire \this_ppu.un1_M_current_q_cry_3 ;
    wire \this_ppu.un1_M_current_q_cry_4 ;
    wire \this_ppu.un1_M_current_q_cry_5 ;
    wire \this_ppu.N_256_1_i ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0 ;
    wire M_this_vga_signals_address_10;
    wire \this_vga_signals.N_9_0_0 ;
    wire \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3Z0Z_5_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0Z0Z_5 ;
    wire \this_vga_signals.N_5 ;
    wire \this_vga_signals.g0_0_x2_0_0_a3_3_cascade_ ;
    wire \this_vga_signals.N_9_i_0_0_cascade_ ;
    wire \this_vga_signals.N_9_i_0_0 ;
    wire \this_vga_signals.g0_2_x0_cascade_ ;
    wire \this_vga_signals.g0_2_x1 ;
    wire \this_vga_signals.N_3_1 ;
    wire \this_vga_signals.m6_2 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_0_0 ;
    wire \this_vga_signals.if_i3_mux_0_0 ;
    wire \this_vga_signals.M_vcounter_q_RNI820378Z0Z_2 ;
    wire \this_vga_signals.N_3_0_cascade_ ;
    wire \this_vga_signals.g1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0 ;
    wire \this_vga_signals.M_vcounter_q_RNI820378_0Z0Z_2 ;
    wire \this_vga_signals.g0_3_0_a3_2_cascade_ ;
    wire \this_vga_signals.g2_1 ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire \this_vga_signals.N_188_0_cascade_ ;
    wire \this_vga_signals.if_m10_0_a4_0_0 ;
    wire \this_vga_signals.g1_3_0_cascade_ ;
    wire \this_vga_signals.if_m10_0_a4_1_1 ;
    wire \this_vga_signals.if_N_18_0 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_1_0_0 ;
    wire bfn_10_14_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_10_15_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.mult1_un40_sum_0_c3_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.mult1_un40_sum_0_c3_0 ;
    wire \this_vga_signals.mult1_un40_sum_1_c2_0 ;
    wire \this_vga_signals.mult1_un40_sum_m_x1_3_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_m_x0_3 ;
    wire \this_vga_signals.CO1_5_0 ;
    wire \this_vga_signals.mult1_un40_sum0_2_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_2_cascade_ ;
    wire \this_vga_signals.N_196_0 ;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0_cascade_;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_cascade_;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0;
    wire this_vga_signals_un4_lcounter_if_i1_mux_cascade_;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_cascade_;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1;
    wire \this_ppu.M_m7Z0Z_1 ;
    wire \this_ppu.M_m12_0_o2_381_10Z0Z_1 ;
    wire \this_ppu.M_N_11_mux_cascade_ ;
    wire \this_ppu.M_m12_0_o2_381_10 ;
    wire this_vga_signals_un4_lcounter_if_i1_mux;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_1;
    wire this_vga_signals_un4_lcounter_if_N_7_i_i;
    wire M_this_ppu_vram_addr_5;
    wire M_this_ppu_vram_addr_4;
    wire M_this_ppu_vram_addr_6;
    wire M_this_ppu_vram_addr_2;
    wire \this_ppu.un1_M_state_d8_4_0_cascade_ ;
    wire \this_ppu.M_N_3_mux_0_0 ;
    wire M_this_ppu_vram_addr_0;
    wire M_this_ppu_vram_addr_3;
    wire M_this_ppu_vram_addr_1;
    wire \this_ppu.un1_M_state_d8_5_0 ;
    wire M_this_sprites_ram_read_data_0_cascade_;
    wire M_this_vram_write_data_0;
    wire port_clk_c;
    wire \this_vga_signals.vsync_1_0_a2_6_a2_1_0 ;
    wire this_vga_signals_vsync_1_i;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire \this_vga_signals.g0_16_x0_cascade_ ;
    wire \this_vga_signals.g3_0 ;
    wire \this_vga_signals.N_57_i_i_0_0 ;
    wire \this_vga_signals.g0_1_0_cascade_ ;
    wire \this_vga_signals.N_5_0_0_1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_3_0_0_0_cascade_ ;
    wire this_vga_signals_address_0_i_7;
    wire \this_vga_signals.N_6_0_0 ;
    wire \this_vga_signals.mult1_un75_sum_c2_0_0_0_1 ;
    wire \this_vga_signals.g3_3_0 ;
    wire \this_vga_signals.g3_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_i_cascade_ ;
    wire \this_vga_signals.g1_2_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ;
    wire \this_vga_signals.g1_1 ;
    wire \this_vga_signals.N_4_i_0_x ;
    wire \this_vga_signals.N_4_i_0_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_3_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.if_m10_0_x2_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c2_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_c3_0_cascade_ ;
    wire \this_vga_signals.if_m2_1 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1 ;
    wire \this_vga_signals.if_m10_0_a4_1_0_x1 ;
    wire \this_vga_signals.if_m10_0_a4_1_0_x0_cascade_ ;
    wire \this_vga_signals.if_m10_0_a4_1 ;
    wire \this_vga_signals.mult1_un54_sum_c2_0 ;
    wire \this_vga_signals.g0_0_a3_0 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNISGOSZ0Z_4_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_1_x1 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_c ;
    wire N_475_cascade_;
    wire \this_vga_signals.if_N_3_mux_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axb2_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_x1 ;
    wire \this_vga_signals.mult1_un47_sum_axb2_0_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_x0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_ns ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_1_0_x1 ;
    wire this_vga_signals_M_vcounter_q_fast_6;
    wire \this_vga_signals.mult1_un40_sum_c3_0_1_0_x0 ;
    wire \this_vga_signals.mult1_un61_sum_axb2_i ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.if_m5_0_1 ;
    wire \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1 ;
    wire \this_vga_signals.mult1_un40_sum_0_axb1_i_cascade_ ;
    wire \this_vga_signals.N_81_0 ;
    wire \this_vga_signals.N_370_0 ;
    wire \this_vga_signals.mult1_un40_sum1_2 ;
    wire this_vga_signals_M_vcounter_q_7_rep1;
    wire this_vga_signals_M_vcounter_q_8_rep1;
    wire \this_vga_signals.N_330_0 ;
    wire \this_vga_signals.vsync_1_0_a2_6_a2_0 ;
    wire \this_vga_signals.if_m11_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_i_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_2_2_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_1_0_x1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_2_2_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_2_2_1_cascade_ ;
    wire this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0;
    wire \this_vga_signals.mult1_un54_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_2 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_sx ;
    wire \this_vga_signals.mult1_un61_sum_ac0_2_4_tz ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_3 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_2_cascade_ ;
    wire this_vga_signals_un4_lcounter_if_i3_mux;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_i ;
    wire \this_vga_signals.g0_16_x1 ;
    wire \this_vga_signals.N_81_1 ;
    wire \this_vga_signals.g1_2 ;
    wire \this_vga_signals.if_N_7_i ;
    wire \this_vga_signals.if_N_11 ;
    wire \this_vga_signals.if_i3_mux_0_1_cascade_ ;
    wire \this_vga_signals.m48_i_x4_3 ;
    wire \this_vga_signals.if_i3_mux_0_1 ;
    wire \this_vga_signals.mult1_un68_sum_axb1_0_0 ;
    wire \this_vga_signals.N_57_0 ;
    wire \this_vga_signals.N_57_i_i_0 ;
    wire \this_vga_signals.g1_0_cascade_ ;
    wire \this_vga_signals.if_N_6_mux_0_0_0 ;
    wire \this_vga_signals.g2_1_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.N_5_i_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i ;
    wire \this_vga_signals.g0_10_1_cascade_ ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_1 ;
    wire \this_vga_signals.if_N_18_1 ;
    wire \this_vga_signals.m48_i_x4_0 ;
    wire \this_vga_signals.mult1_un47_sum_c3_0 ;
    wire \this_vga_signals.g4_1_0 ;
    wire \this_vga_signals.g0_1 ;
    wire bfn_12_12_0_;
    wire \this_vga_signals.mult1_un68_sum_cry_0 ;
    wire \this_vga_signals.mult1_un61_sum_cry_1_s ;
    wire \this_vga_signals.mult1_un68_sum_cry_1 ;
    wire \this_vga_signals.mult1_un68_sum_axb_3 ;
    wire \this_vga_signals.mult1_un68_sum_cry_2 ;
    wire \this_vga_signals.vaddress_8 ;
    wire \this_vga_signals.N_3_2 ;
    wire \this_vga_signals.g1_4 ;
    wire \this_vga_signals.mult1_un61_sum_s_3 ;
    wire \this_vga_signals.mult1_un61_sum_i_3 ;
    wire \this_vga_signals.if_N_3_mux ;
    wire \this_vga_signals.g6_0 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire M_this_vga_signals_address_13;
    wire \this_vga_signals.g0_0 ;
    wire \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0ASZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.mult1_un47_sum_ac0_3_c_0_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ;
    wire \this_vga_signals.M_vcounter_q_9_repZ0Z1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.vaddress_7 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.N_188_0 ;
    wire \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0 ;
    wire \this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0_cascade_ ;
    wire \this_vga_signals.N_188_0_0_0 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_1_0_3 ;
    wire \this_vga_signals.N_188_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_1_0_2_cascade_ ;
    wire \this_vga_signals.g1_0_1 ;
    wire N_183_0;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_0_axb1_i ;
    wire \this_vga_signals.mult1_un40_sum_1_axb1 ;
    wire \this_vga_signals.mult1_un40_sum_m_x0_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_m_x1_1 ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_1 ;
    wire \this_vga_signals.mult1_un40_sum_m_ns_1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.if_N_8_0 ;
    wire \this_vga_signals.mult1_un54_sum_i_0 ;
    wire N_31;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire this_vga_signals_M_vcounter_q_6;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.N_177_0_cascade_ ;
    wire \this_vga_signals.CO0_i_0 ;
    wire \this_vga_signals.N_269_0 ;
    wire \this_vga_signals.N_286 ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1_cascade_;
    wire M_this_delay_clk_out_0;
    wire port_enb_c;
    wire this_start_data_delay_M_last_q;
    wire \this_vga_signals.mult1_un61_sum_i_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1_0 ;
    wire N_90_0;
    wire this_vga_signals_M_vcounter_q_2;
    wire this_vga_signals_M_vcounter_q_3;
    wire N_184_0;
    wire this_vga_signals_M_vcounter_q_1;
    wire N_184_0_cascade_;
    wire this_vga_signals_M_vcounter_q_0;
    wire bfn_13_15_0_;
    wire G_504;
    wire \this_vga_signals.mult1_un75_sum_cry_0 ;
    wire \this_vga_signals.mult1_un68_sum_cry_1_s ;
    wire G_503;
    wire \this_vga_signals.mult1_un75_sum_cry_1 ;
    wire \this_vga_signals.mult1_un75_sum_axb_3 ;
    wire \this_vga_signals.mult1_un75_sum_cry_2 ;
    wire \this_ppu.M_m12_0_o2_381Z0Z_4_cascade_ ;
    wire N_275;
    wire \this_ppu.M_m12_0_o2_381_5_cascade_ ;
    wire N_190_0;
    wire \this_ppu.M_m12_0_o2_381_8 ;
    wire \this_vga_signals.N_336_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.N_287 ;
    wire \this_vga_signals.N_287_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3_cascade_;
    wire \this_vga_signals.mult1_un68_sum_c3_0_1_cascade_ ;
    wire \this_vga_signals.SUM_7_i_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_1 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_2 ;
    wire \this_vga_signals.N_336_0 ;
    wire \this_vga_signals.N_3 ;
    wire \this_vga_signals.mult1_un68_sum_s_3 ;
    wire M_this_vga_signals_pixel_clk_0;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.N_517_1_g ;
    wire \this_vga_signals.N_684_g ;
    wire \this_vga_signals.N_272_0 ;
    wire this_vga_signals_M_vcounter_q_4;
    wire N_475;
    wire this_vga_signals_M_vcounter_q_5;
    wire \this_vga_signals.N_404_0 ;
    wire N_204_0;
    wire bfn_14_17_0_;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_5 ;
    wire this_vga_signals_M_hcounter_q_7;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_6 ;
    wire this_vga_signals_M_hcounter_q_8;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_8 ;
    wire bfn_14_18_0_;
    wire this_vga_signals_M_hcounter_q_9;
    wire \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0 ;
    wire this_vga_signals_M_hcounter_q_6;
    wire \this_vga_signals.N_517_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc1 ;
    wire \this_ppu.sprites_addr_1_i_2_1Z0Z_9 ;
    wire \this_ppu.sprites_addr_1_i_0_0Z0Z_9_cascade_ ;
    wire \this_ppu.sprites_addr_1_i_a0_2Z0Z_9 ;
    wire \this_ppu.sprites_addr_1_i_0_2Z0Z_9_cascade_ ;
    wire N_138_0;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_0_1 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_x0 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_x1 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_1 ;
    wire if_generate_plus_mult1_un68_sum_axbxc3_ns_cascade_;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_cascade_;
    wire this_vga_signals_M_hcounter_q_5;
    wire \this_vga_signals.mult1_un54_sum_axb1_0 ;
    wire this_vga_signals_M_hcounter_q_4;
    wire \this_vga_signals.if_N_8_i_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_axb1_1 ;
    wire M_counter_q_RNIFKS8_0;
    wire M_counter_q_RNIFKS8_0_cascade_;
    wire this_pixel_clk_M_counter_q_i_1;
    wire \this_vga_signals.N_455 ;
    wire \this_vga_signals.N_459 ;
    wire \this_vga_signals.GZ0Z_210_cascade_ ;
    wire this_vga_signals_M_vcounter_q_9;
    wire \this_vga_signals.M_vcounter_q_esr_RNIIRV75Z0Z_9 ;
    wire \this_pixel_clk.M_counter_qZ0Z_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire if_generate_plus_mult1_un75_sum_axbxc3_cascade_;
    wire \this_ppu.un5_sprites_addr_1_c2_cascade_ ;
    wire \this_ppu.N_4_0_1 ;
    wire \this_ppu.sprites_addr_1_i_7_tz_0_9 ;
    wire \this_ppu.sprites_addr_1_i_a7Z0Z_9 ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3;
    wire \this_ppu.un5_sprites_addr1_4 ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0;
    wire \this_vga_signals.GZ0Z_210 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9 ;
    wire this_vga_signals_M_hcounter_q_3;
    wire \this_vga_signals.if_N_9_1 ;
    wire \this_ppu.sprites_m1_0_xZ0Z1 ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3_cascade_;
    wire \this_ppu.sprites_m1_0_xZ0Z0 ;
    wire M_this_internal_address_q_3_ns_1_2;
    wire M_this_internal_address_q_3_ns_1_9;
    wire M_this_internal_address_q_3_ns_1_3_cascade_;
    wire M_this_internal_address_q_3_ns_1_8;
    wire bfn_15_23_0_;
    wire un1_M_this_data_count_q_cry_0;
    wire un1_M_this_data_count_q_cry_1;
    wire un1_M_this_data_count_q_cry_2;
    wire un1_M_this_data_count_q_cry_3;
    wire un1_M_this_data_count_q_cry_4;
    wire un1_M_this_data_count_q_cry_5;
    wire un1_M_this_data_count_q_cry_6;
    wire un1_M_this_data_count_q_cry_7;
    wire bfn_15_24_0_;
    wire un1_M_this_data_count_q_cry_8;
    wire un1_M_this_data_count_q_cry_9;
    wire un1_M_this_data_count_q_cry_10;
    wire un1_M_this_data_count_q_cry_11;
    wire M_this_state_q_RNI20CEZ0Z_0;
    wire un1_M_this_data_count_q_cry_12;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO;
    wire un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO;
    wire bfn_15_25_0_;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire N_13_0;
    wire M_this_vga_signals_address_5;
    wire \this_ppu.un5_sprites_addr_1_c4 ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0_cascade_;
    wire if_generate_plus_mult1_un89_sum_axbxc3;
    wire \this_ppu.sprites_N_7_0_cascade_ ;
    wire \this_ppu.un5_sprites_addr_1_c2 ;
    wire \this_ppu.sprites_m7Z0Z_0_cascade_ ;
    wire if_generate_plus_mult1_un68_sum_axbxc3_ns;
    wire N_140_i;
    wire this_vga_signals_M_hcounter_q_2;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3;
    wire if_generate_plus_mult1_un75_sum_axbxc3;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0;
    wire this_vga_signals_M_hcounter_q_1;
    wire this_vga_signals_M_hcounter_q_0;
    wire \this_ppu.sprites_mZ0Z1_cascade_ ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1;
    wire M_this_internal_address_q_3_ns_1_10_cascade_;
    wire bfn_16_21_0_;
    wire un1_M_this_internal_address_q_cry_0;
    wire M_this_internal_address_qZ0Z_2;
    wire M_this_internal_address_q_RNO_1Z0Z_2;
    wire un1_M_this_internal_address_q_cry_1;
    wire M_this_internal_address_qZ0Z_3;
    wire M_this_internal_address_q_RNO_1Z0Z_3;
    wire un1_M_this_internal_address_q_cry_2;
    wire un1_M_this_internal_address_q_cry_3;
    wire un1_M_this_internal_address_q_cry_4;
    wire un1_M_this_internal_address_q_cry_5;
    wire M_this_internal_address_q_RNO_1Z0Z_7;
    wire un1_M_this_internal_address_q_cry_6;
    wire un1_M_this_internal_address_q_cry_7;
    wire M_this_internal_address_qZ0Z_8;
    wire M_this_internal_address_q_RNO_1Z0Z_8;
    wire bfn_16_22_0_;
    wire M_this_internal_address_qZ0Z_9;
    wire M_this_internal_address_q_RNO_1Z0Z_9;
    wire un1_M_this_internal_address_q_cry_8;
    wire M_this_internal_address_qZ0Z_10;
    wire M_this_internal_address_q_RNO_1Z0Z_10;
    wire un1_M_this_internal_address_q_cry_9;
    wire un1_M_this_internal_address_q_cry_10;
    wire un1_M_this_internal_address_q_cry_11;
    wire un1_M_this_internal_address_q_cry_12;
    wire M_this_internal_address_q_RNO_1Z0Z_13;
    wire M_this_internal_address_qZ0Z_7;
    wire M_this_internal_address_q_3_ns_1_7;
    wire N_235_0_i;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_qZ0Z_0;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_qZ0Z_9;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_qZ0Z_4;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_state_q_srsts_0_a2_1_9_4;
    wire M_this_state_q_srsts_0_a2_1_7_4;
    wire M_this_state_q_srsts_0_a2_1_8_4_cascade_;
    wire M_this_state_q_srsts_0_a2_1_6_4;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0;
    wire this_ppu_sprites_N_2_1;
    wire N_134_0;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4 ;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4_cascade_ ;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_1Z0Z_4 ;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_0Z0Z_4 ;
    wire \this_vga_signals.N_224_0 ;
    wire M_this_state_q_nss_0;
    wire N_235_0;
    wire \this_vga_signals.N_319 ;
    wire un19_i_i_i_a2;
    wire M_this_internal_address_q_RNO_1Z0Z_11;
    wire M_this_internal_address_q_3_ns_1_0;
    wire M_this_internal_address_q_RNO_1Z0Z_0;
    wire M_this_internal_address_qZ0Z_0;
    wire M_this_internal_address_q_3_ns_1_1;
    wire M_this_internal_address_q_RNO_1Z0Z_1;
    wire M_this_internal_address_qZ0Z_1;
    wire N_476;
    wire N_240;
    wire M_this_state_qZ0Z_1;
    wire \this_vga_signals.N_343_cascade_ ;
    wire M_this_state_qZ0Z_2;
    wire M_this_internal_address_q_RNO_1Z0Z_5;
    wire M_this_internal_address_q_RNO_1Z0Z_6;
    wire M_this_internal_address_q_RNO_1Z0Z_12;
    wire M_this_internal_address_q_3_ns_1_11;
    wire M_this_internal_address_q_3_ns_1_4;
    wire M_this_internal_address_q_RNO_1Z0Z_4;
    wire M_this_internal_address_qZ0Z_4;
    wire M_this_vram_write_data_1;
    wire port_address_in_7;
    wire port_address_in_6;
    wire port_rw_in;
    wire \this_vga_signals.N_185_0 ;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4 ;
    wire M_this_state_qZ0Z_4;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4_cascade_ ;
    wire \this_vga_signals.N_490_cascade_ ;
    wire \this_vga_signals.N_386_cascade_ ;
    wire \this_vga_signals.N_387_cascade_ ;
    wire port_address_in_1;
    wire port_address_in_0;
    wire \this_vga_signals.N_391_cascade_ ;
    wire \this_vga_signals.N_490 ;
    wire M_this_state_qZ0Z_5;
    wire M_this_state_qZ0Z_6;
    wire N_14_0;
    wire M_this_internal_address_qZ0Z_5;
    wire M_this_internal_address_q_3_ns_1_5;
    wire M_this_internal_address_qZ0Z_6;
    wire M_this_internal_address_q_3_ns_1_6;
    wire M_this_internal_address_q_3_ns_1_13;
    wire N_355;
    wire M_this_internal_address_q_3_ns_1_12;
    wire M_this_state_qZ0Z_7;
    wire port_data_c_5;
    wire port_data_c_1;
    wire M_this_sprites_ram_write_data_1;
    wire port_data_c_0;
    wire port_data_c_4;
    wire M_this_sprites_ram_write_data_0;
    wire M_this_vram_write_data_2;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire \this_sprites_ram.mem_out_bus6_2 ;
    wire \this_sprites_ram.mem_out_bus2_2 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_ ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ;
    wire M_this_sprites_ram_read_data_2;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ;
    wire M_this_sprites_ram_read_data_1;
    wire \this_sprites_ram.mem_out_bus5_1 ;
    wire \this_sprites_ram.mem_out_bus1_1 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus4_0 ;
    wire \this_sprites_ram.mem_out_bus0_0 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ;
    wire M_this_sprites_ram_read_data_3_cascade_;
    wire M_this_ppu_vram_en_0;
    wire M_this_vram_write_data_3;
    wire \this_sprites_ram.mem_radregZ0Z_11 ;
    wire \this_sprites_ram.mem_radregZ0Z_12 ;
    wire \this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3 ;
    wire \this_sprites_ram.mem_out_bus6_0 ;
    wire \this_sprites_ram.mem_out_bus2_0 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ;
    wire \this_sprites_ram.mem_out_bus5_0 ;
    wire \this_sprites_ram.mem_out_bus1_0 ;
    wire \this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ;
    wire \this_vga_signals.N_483 ;
    wire N_175_0;
    wire \this_sprites_ram.mem_WE_0 ;
    wire \this_sprites_ram.mem_WE_14 ;
    wire \this_sprites_ram.mem_WE_10 ;
    wire \this_sprites_ram.mem_WE_12 ;
    wire \this_sprites_ram.mem_out_bus5_2 ;
    wire \this_sprites_ram.mem_out_bus1_2 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ;
    wire \this_sprites_ram.mem_out_bus4_1 ;
    wire \this_sprites_ram.mem_out_bus0_1 ;
    wire \this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus4_2 ;
    wire \this_sprites_ram.mem_out_bus0_2 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0 ;
    wire \this_sprites_ram.mem_WE_8 ;
    wire \this_sprites_ram.mem_out_bus7_2 ;
    wire \this_sprites_ram.mem_out_bus3_2 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ;
    wire \this_sprites_ram.mem_out_bus7_1 ;
    wire \this_sprites_ram.mem_out_bus3_1 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus6_1 ;
    wire \this_sprites_ram.mem_out_bus2_1 ;
    wire \this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus7_3 ;
    wire \this_sprites_ram.mem_out_bus3_3 ;
    wire \this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ;
    wire \this_sprites_ram.mem_WE_6 ;
    wire port_data_c_3;
    wire port_data_c_7;
    wire M_this_sprites_ram_write_data_3;
    wire \this_sprites_ram.mem_out_bus5_3 ;
    wire \this_sprites_ram.mem_out_bus1_3 ;
    wire \this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus0_3 ;
    wire \this_sprites_ram.mem_out_bus4_3 ;
    wire \this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus6_3 ;
    wire \this_sprites_ram.mem_out_bus2_3 ;
    wire \this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ;
    wire \this_sprites_ram.mem_out_bus7_0 ;
    wire \this_sprites_ram.mem_out_bus3_0 ;
    wire \this_sprites_ram.mem_radregZ0Z_13 ;
    wire \this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ;
    wire \this_vga_signals.N_481 ;
    wire port_data_c_2;
    wire port_data_c_6;
    wire \this_vga_signals.N_479 ;
    wire M_this_sprites_ram_write_data_2;
    wire \this_sprites_ram.mem_WE_4 ;
    wire M_this_internal_address_qZ0Z_12;
    wire M_this_internal_address_qZ0Z_11;
    wire M_this_internal_address_qZ0Z_13;
    wire N_24_0;
    wire \this_sprites_ram.mem_WE_2 ;
    wire N_192_0;
    wire this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2;
    wire \this_ppu.sprites_N_6 ;
    wire sprites_m7;
    wire M_this_state_qZ0Z_3;
    wire M_this_external_address_qZ0Z_0;
    wire bfn_31_23_0_;
    wire M_this_external_address_qZ0Z_1;
    wire un1_M_this_external_address_q_cry_0;
    wire M_this_external_address_qZ0Z_2;
    wire un1_M_this_external_address_q_cry_1;
    wire M_this_external_address_qZ0Z_3;
    wire un1_M_this_external_address_q_cry_2;
    wire M_this_external_address_qZ0Z_4;
    wire un1_M_this_external_address_q_cry_3;
    wire M_this_external_address_qZ0Z_5;
    wire un1_M_this_external_address_q_cry_4;
    wire M_this_external_address_qZ0Z_6;
    wire un1_M_this_external_address_q_cry_5;
    wire M_this_external_address_qZ0Z_7;
    wire un1_M_this_external_address_q_cry_6;
    wire un1_M_this_external_address_q_cry_7;
    wire M_this_external_address_qZ0Z_8;
    wire bfn_31_24_0_;
    wire M_this_external_address_qZ0Z_9;
    wire un1_M_this_external_address_q_cry_8;
    wire M_this_external_address_qZ0Z_10;
    wire un1_M_this_external_address_q_cry_9;
    wire M_this_external_address_qZ0Z_11;
    wire un1_M_this_external_address_q_cry_10;
    wire M_this_external_address_qZ0Z_12;
    wire un1_M_this_external_address_q_cry_11;
    wire M_this_external_address_qZ0Z_13;
    wire un1_M_this_external_address_q_cry_12;
    wire M_this_external_address_qZ0Z_14;
    wire un1_M_this_external_address_q_cry_13;
    wire M_this_state_qZ0Z_0;
    wire un1_M_this_external_address_q_cry_14;
    wire M_this_external_address_qZ0Z_15;
    wire clk_0_c_g;
    wire M_this_state_q_nss_g_0;
    wire port_address_in_2;
    wire port_address_in_3;
    wire port_address_in_4;
    wire port_address_in_5;
    wire \this_vga_signals.M_this_state_q_srsts_0_i_o4_5Z0Z_4 ;
    wire _gnd_net_;

    defparam \this_sprites_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,\this_sprites_ram.mem_out_bus0_1 ,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,\this_sprites_ram.mem_out_bus0_0 ,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__18215,N__16481,N__23654,N__19736,N__10196,N__10478,N__10340,N__10970,N__10049,N__10835,N__11111}),
            .WADDR({N__19058,N__19187,N__19313,N__18899,N__21374,N__21506,N__20366,N__18443,N__18575,N__19964,N__20105}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__20966,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__20789,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__24961),
            .RE(N__17674),
            .WCLKE(N__21866),
            .WCLK(N__24962),
            .WE(N__17492));
    defparam \this_sprites_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,\this_sprites_ram.mem_out_bus0_3 ,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,\this_sprites_ram.mem_out_bus0_2 ,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__18209,N__16475,N__23648,N__19730,N__10190,N__10472,N__10334,N__10964,N__10043,N__10829,N__11105}),
            .WADDR({N__19052,N__19181,N__19307,N__18893,N__21368,N__21500,N__20360,N__18437,N__18569,N__19958,N__20099}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__23107,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__24314,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__24963),
            .RE(N__17673),
            .WCLKE(N__21865),
            .WCLK(N__24964),
            .WE(N__17675));
    defparam \this_sprites_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,\this_sprites_ram.mem_out_bus1_1 ,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,\this_sprites_ram.mem_out_bus1_0 ,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__18203,N__16469,N__23642,N__19724,N__10184,N__10466,N__10328,N__10958,N__10037,N__10823,N__11099}),
            .WADDR({N__19046,N__19175,N__19301,N__18887,N__21362,N__21494,N__20354,N__18431,N__18563,N__19952,N__20093}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__20972,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__20785,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__24967),
            .RE(N__17661),
            .WCLKE(N__22661),
            .WCLK(N__24968),
            .WE(N__17672));
    defparam \this_sprites_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,\this_sprites_ram.mem_out_bus1_3 ,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,\this_sprites_ram.mem_out_bus1_2 ,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__18197,N__16463,N__23636,N__19718,N__10178,N__10460,N__10322,N__10952,N__10031,N__10817,N__11093}),
            .WADDR({N__19040,N__19169,N__19295,N__18881,N__21356,N__21488,N__20348,N__18425,N__18557,N__19946,N__20087}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__23099,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__24310,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__24971),
            .RE(N__17660),
            .WCLKE(N__22660),
            .WCLK(N__24972),
            .WE(N__17671));
    defparam \this_sprites_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,\this_sprites_ram.mem_out_bus2_1 ,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,\this_sprites_ram.mem_out_bus2_0 ,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__18191,N__16457,N__23630,N__19712,N__10172,N__10454,N__10316,N__10946,N__10025,N__10811,N__11087}),
            .WADDR({N__19034,N__19163,N__19289,N__18875,N__21350,N__21482,N__20342,N__18419,N__18551,N__19940,N__20081}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__20968,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__20778,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__24980),
            .RE(N__17637),
            .WCLKE(N__22676),
            .WCLK(N__24979),
            .WE(N__17659));
    defparam \this_sprites_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,\this_sprites_ram.mem_out_bus2_3 ,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,\this_sprites_ram.mem_out_bus2_2 ,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__18185,N__16451,N__23624,N__19706,N__10166,N__10448,N__10310,N__10940,N__10019,N__10805,N__11081}),
            .WADDR({N__19028,N__19157,N__19283,N__18869,N__21344,N__21476,N__20336,N__18413,N__18545,N__19934,N__20075}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__23085,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__24302,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__24992),
            .RE(N__17636),
            .WCLKE(N__22675),
            .WCLK(N__24993),
            .WE(N__17658));
    defparam \this_sprites_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,\this_sprites_ram.mem_out_bus3_1 ,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,\this_sprites_ram.mem_out_bus3_0 ,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__18179,N__16445,N__23618,N__19700,N__10160,N__10442,N__10304,N__10934,N__10013,N__10799,N__11075}),
            .WADDR({N__19022,N__19151,N__19277,N__18863,N__21338,N__21470,N__20330,N__18407,N__18539,N__19928,N__20069}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__20952,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__20767,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__25000),
            .RE(N__17604),
            .WCLKE(N__22537),
            .WCLK(N__25001),
            .WE(N__17631));
    defparam \this_sprites_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,\this_sprites_ram.mem_out_bus3_3 ,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,\this_sprites_ram.mem_out_bus3_2 ,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__18173,N__16439,N__23612,N__19694,N__10154,N__10436,N__10298,N__10928,N__10007,N__10793,N__11069}),
            .WADDR({N__19016,N__19145,N__19271,N__18857,N__21332,N__21464,N__20324,N__18401,N__18533,N__19922,N__20063}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__23067,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__24288,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__25010),
            .RE(N__17603),
            .WCLKE(N__22538),
            .WCLK(N__25011),
            .WE(N__17629));
    defparam \this_sprites_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,\this_sprites_ram.mem_out_bus4_1 ,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,\this_sprites_ram.mem_out_bus4_0 ,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__18167,N__16433,N__23606,N__19688,N__10148,N__10430,N__10292,N__10922,N__10001,N__10787,N__11063}),
            .WADDR({N__19010,N__19139,N__19265,N__18851,N__21326,N__21458,N__20318,N__18395,N__18527,N__19916,N__20057}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__20938,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__20745,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__25019),
            .RE(N__17560),
            .WCLKE(N__23209),
            .WCLK(N__25020),
            .WE(N__17591));
    defparam \this_sprites_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,\this_sprites_ram.mem_out_bus4_3 ,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,\this_sprites_ram.mem_out_bus4_2 ,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__18161,N__16427,N__23600,N__19682,N__10142,N__10424,N__10286,N__10916,N__9995,N__10781,N__11057}),
            .WADDR({N__19004,N__19133,N__19259,N__18845,N__21320,N__21452,N__20312,N__18389,N__18521,N__19910,N__20051}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__23076,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__24248,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__25022),
            .RE(N__17559),
            .WCLKE(N__23213),
            .WCLK(N__25023),
            .WE(N__17549));
    defparam \this_sprites_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,\this_sprites_ram.mem_out_bus5_1 ,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,\this_sprites_ram.mem_out_bus5_0 ,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__18155,N__16421,N__23594,N__19676,N__10136,N__10418,N__10280,N__10910,N__9989,N__10775,N__11051}),
            .WADDR({N__18998,N__19127,N__19253,N__18839,N__21314,N__21446,N__20306,N__18383,N__18515,N__19904,N__20045}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__20939,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__20744,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__25024),
            .RE(N__17503),
            .WCLKE(N__24226),
            .WCLK(N__25025),
            .WE(N__17540));
    defparam \this_sprites_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,\this_sprites_ram.mem_out_bus5_3 ,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,\this_sprites_ram.mem_out_bus5_2 ,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__18149,N__16415,N__23588,N__19670,N__10130,N__10412,N__10274,N__10904,N__9983,N__10769,N__11045}),
            .WADDR({N__18992,N__19121,N__19247,N__18833,N__21308,N__21440,N__20300,N__18377,N__18509,N__19898,N__20039}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__23092,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__24281,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__25026),
            .RE(N__17502),
            .WCLKE(N__24230),
            .WCLK(N__25027),
            .WE(N__17458));
    defparam \this_sprites_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,\this_sprites_ram.mem_out_bus6_1 ,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,\this_sprites_ram.mem_out_bus6_0 ,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__18143,N__16409,N__23582,N__19664,N__10124,N__10406,N__10268,N__10898,N__9977,N__10763,N__11039}),
            .WADDR({N__18986,N__19115,N__19241,N__18827,N__21302,N__21434,N__20294,N__18371,N__18503,N__19892,N__20033}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__20956,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__20763,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__25028),
            .RE(N__17522),
            .WCLKE(N__23878),
            .WCLK(N__25029),
            .WE(N__17533));
    defparam \this_sprites_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,\this_sprites_ram.mem_out_bus6_3 ,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,\this_sprites_ram.mem_out_bus6_2 ,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__18137,N__16403,N__23576,N__19658,N__10118,N__10400,N__10262,N__10892,N__9971,N__10757,N__11033}),
            .WADDR({N__18980,N__19109,N__19235,N__18821,N__21296,N__21428,N__20288,N__18365,N__18497,N__19886,N__20027}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__23103,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__24298,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__25030),
            .RE(N__17523),
            .WCLKE(N__23882),
            .WCLK(N__25031),
            .WE(N__17589));
    defparam \this_sprites_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,\this_sprites_ram.mem_out_bus7_1 ,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,\this_sprites_ram.mem_out_bus7_0 ,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__18131,N__16397,N__23570,N__19652,N__10112,N__10394,N__10256,N__10886,N__9965,N__10751,N__11027}),
            .WADDR({N__18974,N__19103,N__19229,N__18815,N__21290,N__21422,N__20282,N__18359,N__18491,N__19880,N__20021}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__20967,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__20777,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__25032),
            .RE(N__17584),
            .WCLKE(N__21886),
            .WCLK(N__25033),
            .WE(N__17590));
    defparam \this_sprites_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_sprites_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_sprites_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,\this_sprites_ram.mem_out_bus7_3 ,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,\this_sprites_ram.mem_out_bus7_2 ,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__18125,N__16391,N__23564,N__19646,N__10106,N__10388,N__10250,N__10879,N__9959,N__10745,N__11021}),
            .WADDR({N__18968,N__19097,N__19223,N__18809,N__21284,N__21416,N__20276,N__18353,N__18485,N__19874,N__20015}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__23108,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__24309,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__25036),
            .RE(N__17585),
            .WCLKE(N__21890),
            .WCLK(N__25037),
            .WE(N__17630));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_716,dangling_wire_717,dangling_wire_718,N__12761,N__9050,N__9002,N__9491,N__8987,N__9011,N__11156,N__17309}),
            .WADDR({dangling_wire_719,dangling_wire_720,dangling_wire_721,N__14597,N__10099,N__10381,N__10246,N__10882,N__9952,N__10738,N__11017}),
            .MASK({dangling_wire_722,dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737}),
            .WDATA({dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,N__22322,N__21836,N__20240,N__10682}),
            .RCLKE(),
            .RCLK(N__24976),
            .RE(N__17635),
            .WCLKE(N__9116),
            .WCLK(N__24975),
            .WE(N__17598));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__25731),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__25733),
            .DIN(N__25732),
            .DOUT(N__25731),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__25733),
            .PADOUT(N__25732),
            .PADIN(N__25731),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__25722),
            .DIN(N__25721),
            .DOUT(N__25720),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__25722),
            .PADOUT(N__25721),
            .PADIN(N__25720),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__25713),
            .DIN(N__25712),
            .DOUT(N__25711),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__25713),
            .PADOUT(N__25712),
            .PADIN(N__25711),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__25704),
            .DIN(N__25703),
            .DOUT(N__25702),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__25704),
            .PADOUT(N__25703),
            .PADIN(N__25702),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__9464),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__25695),
            .DIN(N__25694),
            .DOUT(N__25693),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__25695),
            .PADOUT(N__25694),
            .PADIN(N__25693),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13829),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__25686),
            .DIN(N__25685),
            .DOUT(N__25684),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__25686),
            .PADOUT(N__25685),
            .PADIN(N__25684),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__23363),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18673));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__25677),
            .DIN(N__25676),
            .DOUT(N__25675),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__25677),
            .PADOUT(N__25676),
            .PADIN(N__25675),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__23336),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18749));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__25668),
            .DIN(N__25667),
            .DOUT(N__25666),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__25668),
            .PADOUT(N__25667),
            .PADIN(N__25666),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__23315),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18729));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__25659),
            .DIN(N__25658),
            .DOUT(N__25657),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__25659),
            .PADOUT(N__25658),
            .PADIN(N__25657),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__23285),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18758));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__25650),
            .DIN(N__25649),
            .DOUT(N__25648),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__25650),
            .PADOUT(N__25649),
            .PADIN(N__25648),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__23261),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18642));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__25641),
            .DIN(N__25640),
            .DOUT(N__25639),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__25641),
            .PADOUT(N__25640),
            .PADIN(N__25639),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__24563),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18715));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__25632),
            .DIN(N__25631),
            .DOUT(N__25630),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__25632),
            .PADOUT(N__25631),
            .PADIN(N__25630),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__24542),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18740));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__25623),
            .DIN(N__25622),
            .DOUT(N__25621),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__25623),
            .PADOUT(N__25622),
            .PADIN(N__25621),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__24521),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18767));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__25614),
            .DIN(N__25613),
            .DOUT(N__25612),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__25614),
            .PADOUT(N__25613),
            .PADIN(N__25612),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24434),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18653));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__25605),
            .DIN(N__25604),
            .DOUT(N__25603),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__25605),
            .PADOUT(N__25604),
            .PADIN(N__25603),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24404),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18759));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__25596),
            .DIN(N__25595),
            .DOUT(N__25594),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__25596),
            .PADOUT(N__25595),
            .PADIN(N__25594),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24377),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18714));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__25587),
            .DIN(N__25586),
            .DOUT(N__25585),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__25587),
            .PADOUT(N__25586),
            .PADIN(N__25585),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__25325),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18716));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__25578),
            .DIN(N__25577),
            .DOUT(N__25576),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__25578),
            .PADOUT(N__25577),
            .PADIN(N__25576),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__25301),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18741));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__25569),
            .DIN(N__25568),
            .DOUT(N__25567),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__25569),
            .PADOUT(N__25568),
            .PADIN(N__25567),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__25061),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18766));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__25560),
            .DIN(N__25559),
            .DOUT(N__25558),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__25560),
            .PADOUT(N__25559),
            .PADIN(N__25558),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24494),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18638));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__25551),
            .DIN(N__25550),
            .DOUT(N__25549),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__25551),
            .PADOUT(N__25550),
            .PADIN(N__25549),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__24464),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18748));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__25542),
            .DIN(N__25541),
            .DOUT(N__25540),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__25542),
            .PADOUT(N__25541),
            .PADIN(N__25540),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__25533),
            .DIN(N__25532),
            .DOUT(N__25531),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__25533),
            .PADOUT(N__25532),
            .PADIN(N__25531),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__25524),
            .DIN(N__25523),
            .DOUT(N__25522),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__25524),
            .PADOUT(N__25523),
            .PADIN(N__25522),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__25515),
            .DIN(N__25514),
            .DOUT(N__25513),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__25515),
            .PADOUT(N__25514),
            .PADIN(N__25513),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__25506),
            .DIN(N__25505),
            .DOUT(N__25504),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__25506),
            .PADOUT(N__25505),
            .PADIN(N__25504),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__25497),
            .DIN(N__25496),
            .DOUT(N__25495),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__25497),
            .PADOUT(N__25496),
            .PADIN(N__25495),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__25488),
            .DIN(N__25487),
            .DOUT(N__25486),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__25488),
            .PADOUT(N__25487),
            .PADIN(N__25486),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__25479),
            .DIN(N__25478),
            .DOUT(N__25477),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__25479),
            .PADOUT(N__25478),
            .PADIN(N__25477),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__25470),
            .DIN(N__25469),
            .DOUT(N__25468),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__25470),
            .PADOUT(N__25469),
            .PADIN(N__25468),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__25461),
            .DIN(N__25460),
            .DOUT(N__25459),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__25461),
            .PADOUT(N__25460),
            .PADIN(N__25459),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8609),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__25452),
            .DIN(N__25451),
            .DOUT(N__25450),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__25452),
            .PADOUT(N__25451),
            .PADIN(N__25450),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__20222),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__25443),
            .DIN(N__25442),
            .DOUT(N__25441),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__25443),
            .PADOUT(N__25442),
            .PADIN(N__25441),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__25434),
            .DIN(N__25433),
            .DOUT(N__25432),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__25434),
            .PADOUT(N__25433),
            .PADIN(N__25432),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8651),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__25425),
            .DIN(N__25424),
            .DOUT(N__25423),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__25425),
            .PADOUT(N__25424),
            .PADIN(N__25423),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__17602),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__18739));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__25416),
            .DIN(N__25415),
            .DOUT(N__25414),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b010101;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__25416),
            .PADOUT(N__25415),
            .PADIN(N__25414),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8603),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__15620),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__25407),
            .DIN(N__25406),
            .DOUT(N__25405),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b010101;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__25407),
            .PADOUT(N__25406),
            .PADIN(N__25405),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8585),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__15609),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__25398),
            .DIN(N__25397),
            .DOUT(N__25396),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b010101;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__25398),
            .PADOUT(N__25397),
            .PADIN(N__25396),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8927),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__15613),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__25389),
            .DIN(N__25388),
            .DOUT(N__25387),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b010101;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__25389),
            .PADOUT(N__25388),
            .PADIN(N__25387),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8969),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__15622),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__25380),
            .DIN(N__25379),
            .DOUT(N__25378),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b010101;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__25380),
            .PADOUT(N__25379),
            .PADIN(N__25378),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8945),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__15621),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__25371),
            .DIN(N__25370),
            .DOUT(N__25369),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b010101;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__25371),
            .PADOUT(N__25370),
            .PADIN(N__25369),
            .CLOCKENABLE(VCCG0),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8672),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(N__15623),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__25362),
            .DIN(N__25361),
            .DOUT(N__25360),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__25362),
            .PADOUT(N__25361),
            .PADIN(N__25360),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__25353),
            .DIN(N__25352),
            .DOUT(N__25351),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__25353),
            .PADOUT(N__25352),
            .PADIN(N__25351),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8636),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__25344),
            .DIN(N__25343),
            .DOUT(N__25342),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__25344),
            .PADOUT(N__25343),
            .PADIN(N__25342),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__10646),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IoInMux I__6214 (
            .O(N__25325),
            .I(N__25322));
    LocalMux I__6213 (
            .O(N__25322),
            .I(N__25319));
    IoSpan4Mux I__6212 (
            .O(N__25319),
            .I(N__25316));
    Span4Mux_s1_h I__6211 (
            .O(N__25316),
            .I(N__25312));
    InMux I__6210 (
            .O(N__25315),
            .I(N__25309));
    Odrv4 I__6209 (
            .O(N__25312),
            .I(M_this_external_address_qZ0Z_13));
    LocalMux I__6208 (
            .O(N__25309),
            .I(M_this_external_address_qZ0Z_13));
    InMux I__6207 (
            .O(N__25304),
            .I(un1_M_this_external_address_q_cry_12));
    IoInMux I__6206 (
            .O(N__25301),
            .I(N__25298));
    LocalMux I__6205 (
            .O(N__25298),
            .I(N__25295));
    Span4Mux_s1_h I__6204 (
            .O(N__25295),
            .I(N__25292));
    Sp12to4 I__6203 (
            .O(N__25292),
            .I(N__25288));
    InMux I__6202 (
            .O(N__25291),
            .I(N__25285));
    Odrv12 I__6201 (
            .O(N__25288),
            .I(M_this_external_address_qZ0Z_14));
    LocalMux I__6200 (
            .O(N__25285),
            .I(M_this_external_address_qZ0Z_14));
    InMux I__6199 (
            .O(N__25280),
            .I(un1_M_this_external_address_q_cry_13));
    InMux I__6198 (
            .O(N__25277),
            .I(N__25265));
    InMux I__6197 (
            .O(N__25276),
            .I(N__25265));
    InMux I__6196 (
            .O(N__25275),
            .I(N__25265));
    InMux I__6195 (
            .O(N__25274),
            .I(N__25265));
    LocalMux I__6194 (
            .O(N__25265),
            .I(N__25248));
    InMux I__6193 (
            .O(N__25264),
            .I(N__25239));
    InMux I__6192 (
            .O(N__25263),
            .I(N__25239));
    InMux I__6191 (
            .O(N__25262),
            .I(N__25239));
    InMux I__6190 (
            .O(N__25261),
            .I(N__25239));
    InMux I__6189 (
            .O(N__25260),
            .I(N__25230));
    InMux I__6188 (
            .O(N__25259),
            .I(N__25230));
    InMux I__6187 (
            .O(N__25258),
            .I(N__25230));
    InMux I__6186 (
            .O(N__25257),
            .I(N__25230));
    InMux I__6185 (
            .O(N__25256),
            .I(N__25221));
    InMux I__6184 (
            .O(N__25255),
            .I(N__25221));
    InMux I__6183 (
            .O(N__25254),
            .I(N__25221));
    InMux I__6182 (
            .O(N__25253),
            .I(N__25221));
    CascadeMux I__6181 (
            .O(N__25252),
            .I(N__25216));
    InMux I__6180 (
            .O(N__25251),
            .I(N__25209));
    Span4Mux_h I__6179 (
            .O(N__25248),
            .I(N__25204));
    LocalMux I__6178 (
            .O(N__25239),
            .I(N__25204));
    LocalMux I__6177 (
            .O(N__25230),
            .I(N__25201));
    LocalMux I__6176 (
            .O(N__25221),
            .I(N__25198));
    InMux I__6175 (
            .O(N__25220),
            .I(N__25193));
    InMux I__6174 (
            .O(N__25219),
            .I(N__25190));
    InMux I__6173 (
            .O(N__25216),
            .I(N__25187));
    InMux I__6172 (
            .O(N__25215),
            .I(N__25182));
    InMux I__6171 (
            .O(N__25214),
            .I(N__25182));
    InMux I__6170 (
            .O(N__25213),
            .I(N__25179));
    InMux I__6169 (
            .O(N__25212),
            .I(N__25176));
    LocalMux I__6168 (
            .O(N__25209),
            .I(N__25173));
    Span4Mux_v I__6167 (
            .O(N__25204),
            .I(N__25170));
    Span4Mux_v I__6166 (
            .O(N__25201),
            .I(N__25165));
    Span4Mux_v I__6165 (
            .O(N__25198),
            .I(N__25165));
    InMux I__6164 (
            .O(N__25197),
            .I(N__25162));
    CascadeMux I__6163 (
            .O(N__25196),
            .I(N__25156));
    LocalMux I__6162 (
            .O(N__25193),
            .I(N__25147));
    LocalMux I__6161 (
            .O(N__25190),
            .I(N__25147));
    LocalMux I__6160 (
            .O(N__25187),
            .I(N__25144));
    LocalMux I__6159 (
            .O(N__25182),
            .I(N__25135));
    LocalMux I__6158 (
            .O(N__25179),
            .I(N__25135));
    LocalMux I__6157 (
            .O(N__25176),
            .I(N__25135));
    Span4Mux_v I__6156 (
            .O(N__25173),
            .I(N__25135));
    Span4Mux_h I__6155 (
            .O(N__25170),
            .I(N__25132));
    Sp12to4 I__6154 (
            .O(N__25165),
            .I(N__25129));
    LocalMux I__6153 (
            .O(N__25162),
            .I(N__25126));
    InMux I__6152 (
            .O(N__25161),
            .I(N__25121));
    InMux I__6151 (
            .O(N__25160),
            .I(N__25121));
    InMux I__6150 (
            .O(N__25159),
            .I(N__25118));
    InMux I__6149 (
            .O(N__25156),
            .I(N__25115));
    InMux I__6148 (
            .O(N__25155),
            .I(N__25110));
    InMux I__6147 (
            .O(N__25154),
            .I(N__25110));
    InMux I__6146 (
            .O(N__25153),
            .I(N__25107));
    InMux I__6145 (
            .O(N__25152),
            .I(N__25104));
    Span4Mux_v I__6144 (
            .O(N__25147),
            .I(N__25097));
    Span4Mux_v I__6143 (
            .O(N__25144),
            .I(N__25097));
    Span4Mux_v I__6142 (
            .O(N__25135),
            .I(N__25097));
    Sp12to4 I__6141 (
            .O(N__25132),
            .I(N__25092));
    Span12Mux_s3_h I__6140 (
            .O(N__25129),
            .I(N__25092));
    Span4Mux_h I__6139 (
            .O(N__25126),
            .I(N__25089));
    LocalMux I__6138 (
            .O(N__25121),
            .I(N__25082));
    LocalMux I__6137 (
            .O(N__25118),
            .I(N__25082));
    LocalMux I__6136 (
            .O(N__25115),
            .I(N__25082));
    LocalMux I__6135 (
            .O(N__25110),
            .I(N__25079));
    LocalMux I__6134 (
            .O(N__25107),
            .I(M_this_state_qZ0Z_0));
    LocalMux I__6133 (
            .O(N__25104),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__6132 (
            .O(N__25097),
            .I(M_this_state_qZ0Z_0));
    Odrv12 I__6131 (
            .O(N__25092),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__6130 (
            .O(N__25089),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__6129 (
            .O(N__25082),
            .I(M_this_state_qZ0Z_0));
    Odrv4 I__6128 (
            .O(N__25079),
            .I(M_this_state_qZ0Z_0));
    InMux I__6127 (
            .O(N__25064),
            .I(un1_M_this_external_address_q_cry_14));
    IoInMux I__6126 (
            .O(N__25061),
            .I(N__25058));
    LocalMux I__6125 (
            .O(N__25058),
            .I(N__25055));
    Span4Mux_s1_h I__6124 (
            .O(N__25055),
            .I(N__25052));
    Sp12to4 I__6123 (
            .O(N__25052),
            .I(N__25049));
    Span12Mux_v I__6122 (
            .O(N__25049),
            .I(N__25045));
    InMux I__6121 (
            .O(N__25048),
            .I(N__25042));
    Odrv12 I__6120 (
            .O(N__25045),
            .I(M_this_external_address_qZ0Z_15));
    LocalMux I__6119 (
            .O(N__25042),
            .I(M_this_external_address_qZ0Z_15));
    ClkMux I__6118 (
            .O(N__25037),
            .I(N__24806));
    ClkMux I__6117 (
            .O(N__25036),
            .I(N__24806));
    ClkMux I__6116 (
            .O(N__25035),
            .I(N__24806));
    ClkMux I__6115 (
            .O(N__25034),
            .I(N__24806));
    ClkMux I__6114 (
            .O(N__25033),
            .I(N__24806));
    ClkMux I__6113 (
            .O(N__25032),
            .I(N__24806));
    ClkMux I__6112 (
            .O(N__25031),
            .I(N__24806));
    ClkMux I__6111 (
            .O(N__25030),
            .I(N__24806));
    ClkMux I__6110 (
            .O(N__25029),
            .I(N__24806));
    ClkMux I__6109 (
            .O(N__25028),
            .I(N__24806));
    ClkMux I__6108 (
            .O(N__25027),
            .I(N__24806));
    ClkMux I__6107 (
            .O(N__25026),
            .I(N__24806));
    ClkMux I__6106 (
            .O(N__25025),
            .I(N__24806));
    ClkMux I__6105 (
            .O(N__25024),
            .I(N__24806));
    ClkMux I__6104 (
            .O(N__25023),
            .I(N__24806));
    ClkMux I__6103 (
            .O(N__25022),
            .I(N__24806));
    ClkMux I__6102 (
            .O(N__25021),
            .I(N__24806));
    ClkMux I__6101 (
            .O(N__25020),
            .I(N__24806));
    ClkMux I__6100 (
            .O(N__25019),
            .I(N__24806));
    ClkMux I__6099 (
            .O(N__25018),
            .I(N__24806));
    ClkMux I__6098 (
            .O(N__25017),
            .I(N__24806));
    ClkMux I__6097 (
            .O(N__25016),
            .I(N__24806));
    ClkMux I__6096 (
            .O(N__25015),
            .I(N__24806));
    ClkMux I__6095 (
            .O(N__25014),
            .I(N__24806));
    ClkMux I__6094 (
            .O(N__25013),
            .I(N__24806));
    ClkMux I__6093 (
            .O(N__25012),
            .I(N__24806));
    ClkMux I__6092 (
            .O(N__25011),
            .I(N__24806));
    ClkMux I__6091 (
            .O(N__25010),
            .I(N__24806));
    ClkMux I__6090 (
            .O(N__25009),
            .I(N__24806));
    ClkMux I__6089 (
            .O(N__25008),
            .I(N__24806));
    ClkMux I__6088 (
            .O(N__25007),
            .I(N__24806));
    ClkMux I__6087 (
            .O(N__25006),
            .I(N__24806));
    ClkMux I__6086 (
            .O(N__25005),
            .I(N__24806));
    ClkMux I__6085 (
            .O(N__25004),
            .I(N__24806));
    ClkMux I__6084 (
            .O(N__25003),
            .I(N__24806));
    ClkMux I__6083 (
            .O(N__25002),
            .I(N__24806));
    ClkMux I__6082 (
            .O(N__25001),
            .I(N__24806));
    ClkMux I__6081 (
            .O(N__25000),
            .I(N__24806));
    ClkMux I__6080 (
            .O(N__24999),
            .I(N__24806));
    ClkMux I__6079 (
            .O(N__24998),
            .I(N__24806));
    ClkMux I__6078 (
            .O(N__24997),
            .I(N__24806));
    ClkMux I__6077 (
            .O(N__24996),
            .I(N__24806));
    ClkMux I__6076 (
            .O(N__24995),
            .I(N__24806));
    ClkMux I__6075 (
            .O(N__24994),
            .I(N__24806));
    ClkMux I__6074 (
            .O(N__24993),
            .I(N__24806));
    ClkMux I__6073 (
            .O(N__24992),
            .I(N__24806));
    ClkMux I__6072 (
            .O(N__24991),
            .I(N__24806));
    ClkMux I__6071 (
            .O(N__24990),
            .I(N__24806));
    ClkMux I__6070 (
            .O(N__24989),
            .I(N__24806));
    ClkMux I__6069 (
            .O(N__24988),
            .I(N__24806));
    ClkMux I__6068 (
            .O(N__24987),
            .I(N__24806));
    ClkMux I__6067 (
            .O(N__24986),
            .I(N__24806));
    ClkMux I__6066 (
            .O(N__24985),
            .I(N__24806));
    ClkMux I__6065 (
            .O(N__24984),
            .I(N__24806));
    ClkMux I__6064 (
            .O(N__24983),
            .I(N__24806));
    ClkMux I__6063 (
            .O(N__24982),
            .I(N__24806));
    ClkMux I__6062 (
            .O(N__24981),
            .I(N__24806));
    ClkMux I__6061 (
            .O(N__24980),
            .I(N__24806));
    ClkMux I__6060 (
            .O(N__24979),
            .I(N__24806));
    ClkMux I__6059 (
            .O(N__24978),
            .I(N__24806));
    ClkMux I__6058 (
            .O(N__24977),
            .I(N__24806));
    ClkMux I__6057 (
            .O(N__24976),
            .I(N__24806));
    ClkMux I__6056 (
            .O(N__24975),
            .I(N__24806));
    ClkMux I__6055 (
            .O(N__24974),
            .I(N__24806));
    ClkMux I__6054 (
            .O(N__24973),
            .I(N__24806));
    ClkMux I__6053 (
            .O(N__24972),
            .I(N__24806));
    ClkMux I__6052 (
            .O(N__24971),
            .I(N__24806));
    ClkMux I__6051 (
            .O(N__24970),
            .I(N__24806));
    ClkMux I__6050 (
            .O(N__24969),
            .I(N__24806));
    ClkMux I__6049 (
            .O(N__24968),
            .I(N__24806));
    ClkMux I__6048 (
            .O(N__24967),
            .I(N__24806));
    ClkMux I__6047 (
            .O(N__24966),
            .I(N__24806));
    ClkMux I__6046 (
            .O(N__24965),
            .I(N__24806));
    ClkMux I__6045 (
            .O(N__24964),
            .I(N__24806));
    ClkMux I__6044 (
            .O(N__24963),
            .I(N__24806));
    ClkMux I__6043 (
            .O(N__24962),
            .I(N__24806));
    ClkMux I__6042 (
            .O(N__24961),
            .I(N__24806));
    GlobalMux I__6041 (
            .O(N__24806),
            .I(N__24803));
    gio2CtrlBuf I__6040 (
            .O(N__24803),
            .I(clk_0_c_g));
    CascadeMux I__6039 (
            .O(N__24800),
            .I(N__24795));
    InMux I__6038 (
            .O(N__24799),
            .I(N__24781));
    InMux I__6037 (
            .O(N__24798),
            .I(N__24778));
    InMux I__6036 (
            .O(N__24795),
            .I(N__24775));
    InMux I__6035 (
            .O(N__24794),
            .I(N__24770));
    InMux I__6034 (
            .O(N__24793),
            .I(N__24770));
    InMux I__6033 (
            .O(N__24792),
            .I(N__24765));
    InMux I__6032 (
            .O(N__24791),
            .I(N__24765));
    InMux I__6031 (
            .O(N__24790),
            .I(N__24762));
    InMux I__6030 (
            .O(N__24789),
            .I(N__24757));
    InMux I__6029 (
            .O(N__24788),
            .I(N__24757));
    InMux I__6028 (
            .O(N__24787),
            .I(N__24754));
    InMux I__6027 (
            .O(N__24786),
            .I(N__24751));
    InMux I__6026 (
            .O(N__24785),
            .I(N__24746));
    InMux I__6025 (
            .O(N__24784),
            .I(N__24746));
    LocalMux I__6024 (
            .O(N__24781),
            .I(N__24728));
    LocalMux I__6023 (
            .O(N__24778),
            .I(N__24725));
    LocalMux I__6022 (
            .O(N__24775),
            .I(N__24722));
    LocalMux I__6021 (
            .O(N__24770),
            .I(N__24719));
    LocalMux I__6020 (
            .O(N__24765),
            .I(N__24716));
    LocalMux I__6019 (
            .O(N__24762),
            .I(N__24713));
    LocalMux I__6018 (
            .O(N__24757),
            .I(N__24710));
    LocalMux I__6017 (
            .O(N__24754),
            .I(N__24707));
    LocalMux I__6016 (
            .O(N__24751),
            .I(N__24704));
    LocalMux I__6015 (
            .O(N__24746),
            .I(N__24701));
    SRMux I__6014 (
            .O(N__24745),
            .I(N__24650));
    SRMux I__6013 (
            .O(N__24744),
            .I(N__24650));
    SRMux I__6012 (
            .O(N__24743),
            .I(N__24650));
    SRMux I__6011 (
            .O(N__24742),
            .I(N__24650));
    SRMux I__6010 (
            .O(N__24741),
            .I(N__24650));
    SRMux I__6009 (
            .O(N__24740),
            .I(N__24650));
    SRMux I__6008 (
            .O(N__24739),
            .I(N__24650));
    SRMux I__6007 (
            .O(N__24738),
            .I(N__24650));
    SRMux I__6006 (
            .O(N__24737),
            .I(N__24650));
    SRMux I__6005 (
            .O(N__24736),
            .I(N__24650));
    SRMux I__6004 (
            .O(N__24735),
            .I(N__24650));
    SRMux I__6003 (
            .O(N__24734),
            .I(N__24650));
    SRMux I__6002 (
            .O(N__24733),
            .I(N__24650));
    SRMux I__6001 (
            .O(N__24732),
            .I(N__24650));
    SRMux I__6000 (
            .O(N__24731),
            .I(N__24650));
    Glb2LocalMux I__5999 (
            .O(N__24728),
            .I(N__24650));
    Glb2LocalMux I__5998 (
            .O(N__24725),
            .I(N__24650));
    Glb2LocalMux I__5997 (
            .O(N__24722),
            .I(N__24650));
    Glb2LocalMux I__5996 (
            .O(N__24719),
            .I(N__24650));
    Glb2LocalMux I__5995 (
            .O(N__24716),
            .I(N__24650));
    Glb2LocalMux I__5994 (
            .O(N__24713),
            .I(N__24650));
    Glb2LocalMux I__5993 (
            .O(N__24710),
            .I(N__24650));
    Glb2LocalMux I__5992 (
            .O(N__24707),
            .I(N__24650));
    Glb2LocalMux I__5991 (
            .O(N__24704),
            .I(N__24650));
    Glb2LocalMux I__5990 (
            .O(N__24701),
            .I(N__24650));
    GlobalMux I__5989 (
            .O(N__24650),
            .I(N__24647));
    gio2CtrlBuf I__5988 (
            .O(N__24647),
            .I(M_this_state_q_nss_g_0));
    InMux I__5987 (
            .O(N__24644),
            .I(N__24641));
    LocalMux I__5986 (
            .O(N__24641),
            .I(N__24638));
    Span12Mux_s10_h I__5985 (
            .O(N__24638),
            .I(N__24635));
    Odrv12 I__5984 (
            .O(N__24635),
            .I(port_address_in_2));
    InMux I__5983 (
            .O(N__24632),
            .I(N__24629));
    LocalMux I__5982 (
            .O(N__24629),
            .I(N__24626));
    Span12Mux_v I__5981 (
            .O(N__24626),
            .I(N__24623));
    Odrv12 I__5980 (
            .O(N__24623),
            .I(port_address_in_3));
    CascadeMux I__5979 (
            .O(N__24620),
            .I(N__24617));
    InMux I__5978 (
            .O(N__24617),
            .I(N__24614));
    LocalMux I__5977 (
            .O(N__24614),
            .I(port_address_in_4));
    InMux I__5976 (
            .O(N__24611),
            .I(N__24608));
    LocalMux I__5975 (
            .O(N__24608),
            .I(N__24605));
    Span4Mux_v I__5974 (
            .O(N__24605),
            .I(N__24602));
    Odrv4 I__5973 (
            .O(N__24602),
            .I(port_address_in_5));
    InMux I__5972 (
            .O(N__24599),
            .I(N__24596));
    LocalMux I__5971 (
            .O(N__24596),
            .I(N__24592));
    InMux I__5970 (
            .O(N__24595),
            .I(N__24589));
    Span4Mux_h I__5969 (
            .O(N__24592),
            .I(N__24586));
    LocalMux I__5968 (
            .O(N__24589),
            .I(N__24583));
    Sp12to4 I__5967 (
            .O(N__24586),
            .I(N__24580));
    Span4Mux_v I__5966 (
            .O(N__24583),
            .I(N__24577));
    Span12Mux_v I__5965 (
            .O(N__24580),
            .I(N__24572));
    Sp12to4 I__5964 (
            .O(N__24577),
            .I(N__24572));
    Span12Mux_h I__5963 (
            .O(N__24572),
            .I(N__24569));
    Odrv12 I__5962 (
            .O(N__24569),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_o4_5Z0Z_4 ));
    InMux I__5961 (
            .O(N__24566),
            .I(un1_M_this_external_address_q_cry_3));
    IoInMux I__5960 (
            .O(N__24563),
            .I(N__24560));
    LocalMux I__5959 (
            .O(N__24560),
            .I(N__24557));
    Span4Mux_s1_h I__5958 (
            .O(N__24557),
            .I(N__24553));
    InMux I__5957 (
            .O(N__24556),
            .I(N__24550));
    Odrv4 I__5956 (
            .O(N__24553),
            .I(M_this_external_address_qZ0Z_5));
    LocalMux I__5955 (
            .O(N__24550),
            .I(M_this_external_address_qZ0Z_5));
    InMux I__5954 (
            .O(N__24545),
            .I(un1_M_this_external_address_q_cry_4));
    IoInMux I__5953 (
            .O(N__24542),
            .I(N__24539));
    LocalMux I__5952 (
            .O(N__24539),
            .I(N__24536));
    Span12Mux_s1_h I__5951 (
            .O(N__24536),
            .I(N__24532));
    InMux I__5950 (
            .O(N__24535),
            .I(N__24529));
    Odrv12 I__5949 (
            .O(N__24532),
            .I(M_this_external_address_qZ0Z_6));
    LocalMux I__5948 (
            .O(N__24529),
            .I(M_this_external_address_qZ0Z_6));
    InMux I__5947 (
            .O(N__24524),
            .I(un1_M_this_external_address_q_cry_5));
    IoInMux I__5946 (
            .O(N__24521),
            .I(N__24518));
    LocalMux I__5945 (
            .O(N__24518),
            .I(N__24515));
    Span4Mux_s1_h I__5944 (
            .O(N__24515),
            .I(N__24512));
    Sp12to4 I__5943 (
            .O(N__24512),
            .I(N__24509));
    Span12Mux_v I__5942 (
            .O(N__24509),
            .I(N__24505));
    InMux I__5941 (
            .O(N__24508),
            .I(N__24502));
    Odrv12 I__5940 (
            .O(N__24505),
            .I(M_this_external_address_qZ0Z_7));
    LocalMux I__5939 (
            .O(N__24502),
            .I(M_this_external_address_qZ0Z_7));
    InMux I__5938 (
            .O(N__24497),
            .I(un1_M_this_external_address_q_cry_6));
    IoInMux I__5937 (
            .O(N__24494),
            .I(N__24491));
    LocalMux I__5936 (
            .O(N__24491),
            .I(N__24488));
    Span4Mux_s0_v I__5935 (
            .O(N__24488),
            .I(N__24485));
    Span4Mux_h I__5934 (
            .O(N__24485),
            .I(N__24482));
    Sp12to4 I__5933 (
            .O(N__24482),
            .I(N__24479));
    Span12Mux_h I__5932 (
            .O(N__24479),
            .I(N__24475));
    InMux I__5931 (
            .O(N__24478),
            .I(N__24472));
    Odrv12 I__5930 (
            .O(N__24475),
            .I(M_this_external_address_qZ0Z_8));
    LocalMux I__5929 (
            .O(N__24472),
            .I(M_this_external_address_qZ0Z_8));
    InMux I__5928 (
            .O(N__24467),
            .I(bfn_31_24_0_));
    IoInMux I__5927 (
            .O(N__24464),
            .I(N__24461));
    LocalMux I__5926 (
            .O(N__24461),
            .I(N__24458));
    IoSpan4Mux I__5925 (
            .O(N__24458),
            .I(N__24455));
    IoSpan4Mux I__5924 (
            .O(N__24455),
            .I(N__24452));
    IoSpan4Mux I__5923 (
            .O(N__24452),
            .I(N__24449));
    IoSpan4Mux I__5922 (
            .O(N__24449),
            .I(N__24445));
    InMux I__5921 (
            .O(N__24448),
            .I(N__24442));
    Odrv4 I__5920 (
            .O(N__24445),
            .I(M_this_external_address_qZ0Z_9));
    LocalMux I__5919 (
            .O(N__24442),
            .I(M_this_external_address_qZ0Z_9));
    InMux I__5918 (
            .O(N__24437),
            .I(un1_M_this_external_address_q_cry_8));
    IoInMux I__5917 (
            .O(N__24434),
            .I(N__24431));
    LocalMux I__5916 (
            .O(N__24431),
            .I(N__24428));
    Span4Mux_s2_v I__5915 (
            .O(N__24428),
            .I(N__24425));
    Span4Mux_v I__5914 (
            .O(N__24425),
            .I(N__24422));
    Sp12to4 I__5913 (
            .O(N__24422),
            .I(N__24419));
    Span12Mux_h I__5912 (
            .O(N__24419),
            .I(N__24415));
    InMux I__5911 (
            .O(N__24418),
            .I(N__24412));
    Odrv12 I__5910 (
            .O(N__24415),
            .I(M_this_external_address_qZ0Z_10));
    LocalMux I__5909 (
            .O(N__24412),
            .I(M_this_external_address_qZ0Z_10));
    InMux I__5908 (
            .O(N__24407),
            .I(un1_M_this_external_address_q_cry_9));
    IoInMux I__5907 (
            .O(N__24404),
            .I(N__24401));
    LocalMux I__5906 (
            .O(N__24401),
            .I(N__24398));
    Span4Mux_s0_v I__5905 (
            .O(N__24398),
            .I(N__24395));
    Span4Mux_v I__5904 (
            .O(N__24395),
            .I(N__24392));
    Span4Mux_v I__5903 (
            .O(N__24392),
            .I(N__24388));
    InMux I__5902 (
            .O(N__24391),
            .I(N__24385));
    Odrv4 I__5901 (
            .O(N__24388),
            .I(M_this_external_address_qZ0Z_11));
    LocalMux I__5900 (
            .O(N__24385),
            .I(M_this_external_address_qZ0Z_11));
    InMux I__5899 (
            .O(N__24380),
            .I(un1_M_this_external_address_q_cry_10));
    IoInMux I__5898 (
            .O(N__24377),
            .I(N__24374));
    LocalMux I__5897 (
            .O(N__24374),
            .I(N__24370));
    InMux I__5896 (
            .O(N__24373),
            .I(N__24367));
    Odrv12 I__5895 (
            .O(N__24370),
            .I(M_this_external_address_qZ0Z_12));
    LocalMux I__5894 (
            .O(N__24367),
            .I(M_this_external_address_qZ0Z_12));
    InMux I__5893 (
            .O(N__24362),
            .I(un1_M_this_external_address_q_cry_11));
    InMux I__5892 (
            .O(N__24359),
            .I(N__24355));
    InMux I__5891 (
            .O(N__24358),
            .I(N__24351));
    LocalMux I__5890 (
            .O(N__24355),
            .I(N__24348));
    InMux I__5889 (
            .O(N__24354),
            .I(N__24345));
    LocalMux I__5888 (
            .O(N__24351),
            .I(N__24341));
    Span4Mux_h I__5887 (
            .O(N__24348),
            .I(N__24338));
    LocalMux I__5886 (
            .O(N__24345),
            .I(N__24335));
    InMux I__5885 (
            .O(N__24344),
            .I(N__24332));
    Span12Mux_h I__5884 (
            .O(N__24341),
            .I(N__24329));
    Span4Mux_h I__5883 (
            .O(N__24338),
            .I(N__24326));
    Span4Mux_v I__5882 (
            .O(N__24335),
            .I(N__24321));
    LocalMux I__5881 (
            .O(N__24332),
            .I(N__24321));
    Odrv12 I__5880 (
            .O(N__24329),
            .I(\this_vga_signals.N_479 ));
    Odrv4 I__5879 (
            .O(N__24326),
            .I(\this_vga_signals.N_479 ));
    Odrv4 I__5878 (
            .O(N__24321),
            .I(\this_vga_signals.N_479 ));
    InMux I__5877 (
            .O(N__24314),
            .I(N__24311));
    LocalMux I__5876 (
            .O(N__24311),
            .I(N__24306));
    InMux I__5875 (
            .O(N__24310),
            .I(N__24303));
    InMux I__5874 (
            .O(N__24309),
            .I(N__24299));
    Span4Mux_h I__5873 (
            .O(N__24306),
            .I(N__24295));
    LocalMux I__5872 (
            .O(N__24303),
            .I(N__24292));
    InMux I__5871 (
            .O(N__24302),
            .I(N__24289));
    LocalMux I__5870 (
            .O(N__24299),
            .I(N__24285));
    InMux I__5869 (
            .O(N__24298),
            .I(N__24282));
    Span4Mux_v I__5868 (
            .O(N__24295),
            .I(N__24276));
    Span4Mux_h I__5867 (
            .O(N__24292),
            .I(N__24276));
    LocalMux I__5866 (
            .O(N__24289),
            .I(N__24273));
    InMux I__5865 (
            .O(N__24288),
            .I(N__24270));
    Span4Mux_v I__5864 (
            .O(N__24285),
            .I(N__24265));
    LocalMux I__5863 (
            .O(N__24282),
            .I(N__24265));
    InMux I__5862 (
            .O(N__24281),
            .I(N__24262));
    Span4Mux_v I__5861 (
            .O(N__24276),
            .I(N__24257));
    Span4Mux_h I__5860 (
            .O(N__24273),
            .I(N__24257));
    LocalMux I__5859 (
            .O(N__24270),
            .I(N__24254));
    Span4Mux_v I__5858 (
            .O(N__24265),
            .I(N__24249));
    LocalMux I__5857 (
            .O(N__24262),
            .I(N__24249));
    Span4Mux_v I__5856 (
            .O(N__24257),
            .I(N__24243));
    Span4Mux_h I__5855 (
            .O(N__24254),
            .I(N__24243));
    Span4Mux_v I__5854 (
            .O(N__24249),
            .I(N__24240));
    InMux I__5853 (
            .O(N__24248),
            .I(N__24237));
    Odrv4 I__5852 (
            .O(N__24243),
            .I(M_this_sprites_ram_write_data_2));
    Odrv4 I__5851 (
            .O(N__24240),
            .I(M_this_sprites_ram_write_data_2));
    LocalMux I__5850 (
            .O(N__24237),
            .I(M_this_sprites_ram_write_data_2));
    CEMux I__5849 (
            .O(N__24230),
            .I(N__24227));
    LocalMux I__5848 (
            .O(N__24227),
            .I(N__24223));
    CEMux I__5847 (
            .O(N__24226),
            .I(N__24220));
    Span4Mux_h I__5846 (
            .O(N__24223),
            .I(N__24217));
    LocalMux I__5845 (
            .O(N__24220),
            .I(N__24214));
    Odrv4 I__5844 (
            .O(N__24217),
            .I(\this_sprites_ram.mem_WE_4 ));
    Odrv12 I__5843 (
            .O(N__24214),
            .I(\this_sprites_ram.mem_WE_4 ));
    InMux I__5842 (
            .O(N__24209),
            .I(N__24203));
    InMux I__5841 (
            .O(N__24208),
            .I(N__24198));
    InMux I__5840 (
            .O(N__24207),
            .I(N__24198));
    InMux I__5839 (
            .O(N__24206),
            .I(N__24195));
    LocalMux I__5838 (
            .O(N__24203),
            .I(N__24191));
    LocalMux I__5837 (
            .O(N__24198),
            .I(N__24186));
    LocalMux I__5836 (
            .O(N__24195),
            .I(N__24186));
    InMux I__5835 (
            .O(N__24194),
            .I(N__24183));
    Span4Mux_v I__5834 (
            .O(N__24191),
            .I(N__24176));
    Span4Mux_v I__5833 (
            .O(N__24186),
            .I(N__24176));
    LocalMux I__5832 (
            .O(N__24183),
            .I(N__24176));
    Span4Mux_v I__5831 (
            .O(N__24176),
            .I(N__24170));
    InMux I__5830 (
            .O(N__24175),
            .I(N__24164));
    InMux I__5829 (
            .O(N__24174),
            .I(N__24164));
    InMux I__5828 (
            .O(N__24173),
            .I(N__24161));
    Span4Mux_v I__5827 (
            .O(N__24170),
            .I(N__24157));
    InMux I__5826 (
            .O(N__24169),
            .I(N__24154));
    LocalMux I__5825 (
            .O(N__24164),
            .I(N__24149));
    LocalMux I__5824 (
            .O(N__24161),
            .I(N__24149));
    InMux I__5823 (
            .O(N__24160),
            .I(N__24146));
    Span4Mux_h I__5822 (
            .O(N__24157),
            .I(N__24141));
    LocalMux I__5821 (
            .O(N__24154),
            .I(N__24141));
    Odrv12 I__5820 (
            .O(N__24149),
            .I(M_this_internal_address_qZ0Z_12));
    LocalMux I__5819 (
            .O(N__24146),
            .I(M_this_internal_address_qZ0Z_12));
    Odrv4 I__5818 (
            .O(N__24141),
            .I(M_this_internal_address_qZ0Z_12));
    CascadeMux I__5817 (
            .O(N__24134),
            .I(N__24131));
    InMux I__5816 (
            .O(N__24131),
            .I(N__24124));
    InMux I__5815 (
            .O(N__24130),
            .I(N__24124));
    InMux I__5814 (
            .O(N__24129),
            .I(N__24121));
    LocalMux I__5813 (
            .O(N__24124),
            .I(N__24115));
    LocalMux I__5812 (
            .O(N__24121),
            .I(N__24115));
    InMux I__5811 (
            .O(N__24120),
            .I(N__24112));
    Span4Mux_v I__5810 (
            .O(N__24115),
            .I(N__24107));
    LocalMux I__5809 (
            .O(N__24112),
            .I(N__24107));
    Span4Mux_h I__5808 (
            .O(N__24107),
            .I(N__24104));
    Span4Mux_v I__5807 (
            .O(N__24104),
            .I(N__24100));
    InMux I__5806 (
            .O(N__24103),
            .I(N__24097));
    Sp12to4 I__5805 (
            .O(N__24100),
            .I(N__24089));
    LocalMux I__5804 (
            .O(N__24097),
            .I(N__24089));
    InMux I__5803 (
            .O(N__24096),
            .I(N__24084));
    InMux I__5802 (
            .O(N__24095),
            .I(N__24084));
    InMux I__5801 (
            .O(N__24094),
            .I(N__24081));
    Span12Mux_h I__5800 (
            .O(N__24089),
            .I(N__24076));
    LocalMux I__5799 (
            .O(N__24084),
            .I(N__24071));
    LocalMux I__5798 (
            .O(N__24081),
            .I(N__24071));
    InMux I__5797 (
            .O(N__24080),
            .I(N__24068));
    InMux I__5796 (
            .O(N__24079),
            .I(N__24065));
    Odrv12 I__5795 (
            .O(N__24076),
            .I(M_this_internal_address_qZ0Z_11));
    Odrv12 I__5794 (
            .O(N__24071),
            .I(M_this_internal_address_qZ0Z_11));
    LocalMux I__5793 (
            .O(N__24068),
            .I(M_this_internal_address_qZ0Z_11));
    LocalMux I__5792 (
            .O(N__24065),
            .I(M_this_internal_address_qZ0Z_11));
    CascadeMux I__5791 (
            .O(N__24056),
            .I(N__24048));
    CascadeMux I__5790 (
            .O(N__24055),
            .I(N__24045));
    CascadeMux I__5789 (
            .O(N__24054),
            .I(N__24042));
    CascadeMux I__5788 (
            .O(N__24053),
            .I(N__24038));
    CascadeMux I__5787 (
            .O(N__24052),
            .I(N__24035));
    CascadeMux I__5786 (
            .O(N__24051),
            .I(N__24031));
    InMux I__5785 (
            .O(N__24048),
            .I(N__24027));
    InMux I__5784 (
            .O(N__24045),
            .I(N__24022));
    InMux I__5783 (
            .O(N__24042),
            .I(N__24022));
    CascadeMux I__5782 (
            .O(N__24041),
            .I(N__24019));
    InMux I__5781 (
            .O(N__24038),
            .I(N__24016));
    InMux I__5780 (
            .O(N__24035),
            .I(N__24013));
    InMux I__5779 (
            .O(N__24034),
            .I(N__24008));
    InMux I__5778 (
            .O(N__24031),
            .I(N__24008));
    InMux I__5777 (
            .O(N__24030),
            .I(N__24005));
    LocalMux I__5776 (
            .O(N__24027),
            .I(N__24002));
    LocalMux I__5775 (
            .O(N__24022),
            .I(N__23999));
    InMux I__5774 (
            .O(N__24019),
            .I(N__23996));
    LocalMux I__5773 (
            .O(N__24016),
            .I(N__23989));
    LocalMux I__5772 (
            .O(N__24013),
            .I(N__23989));
    LocalMux I__5771 (
            .O(N__24008),
            .I(N__23989));
    LocalMux I__5770 (
            .O(N__24005),
            .I(N__23985));
    Span4Mux_h I__5769 (
            .O(N__24002),
            .I(N__23982));
    Span4Mux_v I__5768 (
            .O(N__23999),
            .I(N__23979));
    LocalMux I__5767 (
            .O(N__23996),
            .I(N__23976));
    Span4Mux_v I__5766 (
            .O(N__23989),
            .I(N__23973));
    InMux I__5765 (
            .O(N__23988),
            .I(N__23970));
    Span4Mux_v I__5764 (
            .O(N__23985),
            .I(N__23963));
    Span4Mux_v I__5763 (
            .O(N__23982),
            .I(N__23963));
    Span4Mux_h I__5762 (
            .O(N__23979),
            .I(N__23963));
    Span4Mux_v I__5761 (
            .O(N__23976),
            .I(N__23960));
    Sp12to4 I__5760 (
            .O(N__23973),
            .I(N__23957));
    LocalMux I__5759 (
            .O(N__23970),
            .I(N__23950));
    Sp12to4 I__5758 (
            .O(N__23963),
            .I(N__23950));
    Sp12to4 I__5757 (
            .O(N__23960),
            .I(N__23950));
    Span12Mux_h I__5756 (
            .O(N__23957),
            .I(N__23947));
    Odrv12 I__5755 (
            .O(N__23950),
            .I(M_this_internal_address_qZ0Z_13));
    Odrv12 I__5754 (
            .O(N__23947),
            .I(M_this_internal_address_qZ0Z_13));
    InMux I__5753 (
            .O(N__23942),
            .I(N__23935));
    InMux I__5752 (
            .O(N__23941),
            .I(N__23935));
    InMux I__5751 (
            .O(N__23940),
            .I(N__23932));
    LocalMux I__5750 (
            .O(N__23935),
            .I(N__23926));
    LocalMux I__5749 (
            .O(N__23932),
            .I(N__23923));
    InMux I__5748 (
            .O(N__23931),
            .I(N__23920));
    InMux I__5747 (
            .O(N__23930),
            .I(N__23913));
    InMux I__5746 (
            .O(N__23929),
            .I(N__23913));
    Span4Mux_v I__5745 (
            .O(N__23926),
            .I(N__23906));
    Span4Mux_h I__5744 (
            .O(N__23923),
            .I(N__23906));
    LocalMux I__5743 (
            .O(N__23920),
            .I(N__23906));
    InMux I__5742 (
            .O(N__23919),
            .I(N__23903));
    InMux I__5741 (
            .O(N__23918),
            .I(N__23900));
    LocalMux I__5740 (
            .O(N__23913),
            .I(N__23897));
    Span4Mux_v I__5739 (
            .O(N__23906),
            .I(N__23892));
    LocalMux I__5738 (
            .O(N__23903),
            .I(N__23892));
    LocalMux I__5737 (
            .O(N__23900),
            .I(N__23889));
    Odrv4 I__5736 (
            .O(N__23897),
            .I(N_24_0));
    Odrv4 I__5735 (
            .O(N__23892),
            .I(N_24_0));
    Odrv4 I__5734 (
            .O(N__23889),
            .I(N_24_0));
    CEMux I__5733 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__5732 (
            .O(N__23879),
            .I(N__23875));
    CEMux I__5731 (
            .O(N__23878),
            .I(N__23872));
    Span4Mux_v I__5730 (
            .O(N__23875),
            .I(N__23867));
    LocalMux I__5729 (
            .O(N__23872),
            .I(N__23867));
    Span4Mux_v I__5728 (
            .O(N__23867),
            .I(N__23864));
    Odrv4 I__5727 (
            .O(N__23864),
            .I(\this_sprites_ram.mem_WE_2 ));
    CascadeMux I__5726 (
            .O(N__23861),
            .I(N__23847));
    InMux I__5725 (
            .O(N__23860),
            .I(N__23844));
    InMux I__5724 (
            .O(N__23859),
            .I(N__23839));
    InMux I__5723 (
            .O(N__23858),
            .I(N__23834));
    InMux I__5722 (
            .O(N__23857),
            .I(N__23834));
    CascadeMux I__5721 (
            .O(N__23856),
            .I(N__23831));
    InMux I__5720 (
            .O(N__23855),
            .I(N__23827));
    InMux I__5719 (
            .O(N__23854),
            .I(N__23824));
    InMux I__5718 (
            .O(N__23853),
            .I(N__23818));
    InMux I__5717 (
            .O(N__23852),
            .I(N__23818));
    InMux I__5716 (
            .O(N__23851),
            .I(N__23815));
    InMux I__5715 (
            .O(N__23850),
            .I(N__23812));
    InMux I__5714 (
            .O(N__23847),
            .I(N__23809));
    LocalMux I__5713 (
            .O(N__23844),
            .I(N__23806));
    CascadeMux I__5712 (
            .O(N__23843),
            .I(N__23803));
    InMux I__5711 (
            .O(N__23842),
            .I(N__23800));
    LocalMux I__5710 (
            .O(N__23839),
            .I(N__23797));
    LocalMux I__5709 (
            .O(N__23834),
            .I(N__23794));
    InMux I__5708 (
            .O(N__23831),
            .I(N__23789));
    InMux I__5707 (
            .O(N__23830),
            .I(N__23789));
    LocalMux I__5706 (
            .O(N__23827),
            .I(N__23786));
    LocalMux I__5705 (
            .O(N__23824),
            .I(N__23783));
    InMux I__5704 (
            .O(N__23823),
            .I(N__23780));
    LocalMux I__5703 (
            .O(N__23818),
            .I(N__23777));
    LocalMux I__5702 (
            .O(N__23815),
            .I(N__23772));
    LocalMux I__5701 (
            .O(N__23812),
            .I(N__23772));
    LocalMux I__5700 (
            .O(N__23809),
            .I(N__23769));
    Span4Mux_v I__5699 (
            .O(N__23806),
            .I(N__23766));
    InMux I__5698 (
            .O(N__23803),
            .I(N__23763));
    LocalMux I__5697 (
            .O(N__23800),
            .I(N__23760));
    Span4Mux_v I__5696 (
            .O(N__23797),
            .I(N__23753));
    Span4Mux_v I__5695 (
            .O(N__23794),
            .I(N__23753));
    LocalMux I__5694 (
            .O(N__23789),
            .I(N__23753));
    Span12Mux_s7_v I__5693 (
            .O(N__23786),
            .I(N__23750));
    Sp12to4 I__5692 (
            .O(N__23783),
            .I(N__23747));
    LocalMux I__5691 (
            .O(N__23780),
            .I(N__23744));
    Span4Mux_v I__5690 (
            .O(N__23777),
            .I(N__23739));
    Span4Mux_v I__5689 (
            .O(N__23772),
            .I(N__23739));
    Span4Mux_v I__5688 (
            .O(N__23769),
            .I(N__23736));
    Span4Mux_h I__5687 (
            .O(N__23766),
            .I(N__23731));
    LocalMux I__5686 (
            .O(N__23763),
            .I(N__23731));
    Span4Mux_v I__5685 (
            .O(N__23760),
            .I(N__23728));
    Span4Mux_h I__5684 (
            .O(N__23753),
            .I(N__23725));
    Span12Mux_h I__5683 (
            .O(N__23750),
            .I(N__23718));
    Span12Mux_v I__5682 (
            .O(N__23747),
            .I(N__23718));
    Span12Mux_s11_h I__5681 (
            .O(N__23744),
            .I(N__23718));
    Span4Mux_v I__5680 (
            .O(N__23739),
            .I(N__23709));
    Span4Mux_h I__5679 (
            .O(N__23736),
            .I(N__23709));
    Span4Mux_v I__5678 (
            .O(N__23731),
            .I(N__23709));
    Span4Mux_h I__5677 (
            .O(N__23728),
            .I(N__23709));
    Odrv4 I__5676 (
            .O(N__23725),
            .I(N_192_0));
    Odrv12 I__5675 (
            .O(N__23718),
            .I(N_192_0));
    Odrv4 I__5674 (
            .O(N__23709),
            .I(N_192_0));
    InMux I__5673 (
            .O(N__23702),
            .I(N__23699));
    LocalMux I__5672 (
            .O(N__23699),
            .I(N__23696));
    Span12Mux_h I__5671 (
            .O(N__23696),
            .I(N__23693));
    Span12Mux_v I__5670 (
            .O(N__23693),
            .I(N__23687));
    InMux I__5669 (
            .O(N__23692),
            .I(N__23684));
    InMux I__5668 (
            .O(N__23691),
            .I(N__23681));
    InMux I__5667 (
            .O(N__23690),
            .I(N__23678));
    Odrv12 I__5666 (
            .O(N__23687),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2));
    LocalMux I__5665 (
            .O(N__23684),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2));
    LocalMux I__5664 (
            .O(N__23681),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2));
    LocalMux I__5663 (
            .O(N__23678),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2));
    InMux I__5662 (
            .O(N__23669),
            .I(N__23666));
    LocalMux I__5661 (
            .O(N__23666),
            .I(N__23663));
    Span12Mux_h I__5660 (
            .O(N__23663),
            .I(N__23660));
    Span12Mux_v I__5659 (
            .O(N__23660),
            .I(N__23657));
    Odrv12 I__5658 (
            .O(N__23657),
            .I(\this_ppu.sprites_N_6 ));
    CascadeMux I__5657 (
            .O(N__23654),
            .I(N__23651));
    CascadeBuf I__5656 (
            .O(N__23651),
            .I(N__23648));
    CascadeMux I__5655 (
            .O(N__23648),
            .I(N__23645));
    CascadeBuf I__5654 (
            .O(N__23645),
            .I(N__23642));
    CascadeMux I__5653 (
            .O(N__23642),
            .I(N__23639));
    CascadeBuf I__5652 (
            .O(N__23639),
            .I(N__23636));
    CascadeMux I__5651 (
            .O(N__23636),
            .I(N__23633));
    CascadeBuf I__5650 (
            .O(N__23633),
            .I(N__23630));
    CascadeMux I__5649 (
            .O(N__23630),
            .I(N__23627));
    CascadeBuf I__5648 (
            .O(N__23627),
            .I(N__23624));
    CascadeMux I__5647 (
            .O(N__23624),
            .I(N__23621));
    CascadeBuf I__5646 (
            .O(N__23621),
            .I(N__23618));
    CascadeMux I__5645 (
            .O(N__23618),
            .I(N__23615));
    CascadeBuf I__5644 (
            .O(N__23615),
            .I(N__23612));
    CascadeMux I__5643 (
            .O(N__23612),
            .I(N__23609));
    CascadeBuf I__5642 (
            .O(N__23609),
            .I(N__23606));
    CascadeMux I__5641 (
            .O(N__23606),
            .I(N__23603));
    CascadeBuf I__5640 (
            .O(N__23603),
            .I(N__23600));
    CascadeMux I__5639 (
            .O(N__23600),
            .I(N__23597));
    CascadeBuf I__5638 (
            .O(N__23597),
            .I(N__23594));
    CascadeMux I__5637 (
            .O(N__23594),
            .I(N__23591));
    CascadeBuf I__5636 (
            .O(N__23591),
            .I(N__23588));
    CascadeMux I__5635 (
            .O(N__23588),
            .I(N__23585));
    CascadeBuf I__5634 (
            .O(N__23585),
            .I(N__23582));
    CascadeMux I__5633 (
            .O(N__23582),
            .I(N__23579));
    CascadeBuf I__5632 (
            .O(N__23579),
            .I(N__23576));
    CascadeMux I__5631 (
            .O(N__23576),
            .I(N__23573));
    CascadeBuf I__5630 (
            .O(N__23573),
            .I(N__23570));
    CascadeMux I__5629 (
            .O(N__23570),
            .I(N__23567));
    CascadeBuf I__5628 (
            .O(N__23567),
            .I(N__23564));
    CascadeMux I__5627 (
            .O(N__23564),
            .I(N__23561));
    InMux I__5626 (
            .O(N__23561),
            .I(N__23558));
    LocalMux I__5625 (
            .O(N__23558),
            .I(N__23555));
    Odrv4 I__5624 (
            .O(N__23555),
            .I(sprites_m7));
    InMux I__5623 (
            .O(N__23552),
            .I(N__23549));
    LocalMux I__5622 (
            .O(N__23549),
            .I(N__23537));
    CascadeMux I__5621 (
            .O(N__23548),
            .I(N__23531));
    CascadeMux I__5620 (
            .O(N__23547),
            .I(N__23527));
    CascadeMux I__5619 (
            .O(N__23546),
            .I(N__23523));
    CascadeMux I__5618 (
            .O(N__23545),
            .I(N__23519));
    CascadeMux I__5617 (
            .O(N__23544),
            .I(N__23516));
    InMux I__5616 (
            .O(N__23543),
            .I(N__23513));
    CascadeMux I__5615 (
            .O(N__23542),
            .I(N__23510));
    CascadeMux I__5614 (
            .O(N__23541),
            .I(N__23506));
    CascadeMux I__5613 (
            .O(N__23540),
            .I(N__23502));
    Span4Mux_h I__5612 (
            .O(N__23537),
            .I(N__23497));
    InMux I__5611 (
            .O(N__23536),
            .I(N__23494));
    InMux I__5610 (
            .O(N__23535),
            .I(N__23491));
    InMux I__5609 (
            .O(N__23534),
            .I(N__23474));
    InMux I__5608 (
            .O(N__23531),
            .I(N__23474));
    InMux I__5607 (
            .O(N__23530),
            .I(N__23474));
    InMux I__5606 (
            .O(N__23527),
            .I(N__23474));
    InMux I__5605 (
            .O(N__23526),
            .I(N__23474));
    InMux I__5604 (
            .O(N__23523),
            .I(N__23474));
    InMux I__5603 (
            .O(N__23522),
            .I(N__23474));
    InMux I__5602 (
            .O(N__23519),
            .I(N__23474));
    InMux I__5601 (
            .O(N__23516),
            .I(N__23471));
    LocalMux I__5600 (
            .O(N__23513),
            .I(N__23467));
    InMux I__5599 (
            .O(N__23510),
            .I(N__23456));
    InMux I__5598 (
            .O(N__23509),
            .I(N__23456));
    InMux I__5597 (
            .O(N__23506),
            .I(N__23456));
    InMux I__5596 (
            .O(N__23505),
            .I(N__23456));
    InMux I__5595 (
            .O(N__23502),
            .I(N__23456));
    InMux I__5594 (
            .O(N__23501),
            .I(N__23453));
    InMux I__5593 (
            .O(N__23500),
            .I(N__23450));
    Span4Mux_h I__5592 (
            .O(N__23497),
            .I(N__23447));
    LocalMux I__5591 (
            .O(N__23494),
            .I(N__23444));
    LocalMux I__5590 (
            .O(N__23491),
            .I(N__23441));
    LocalMux I__5589 (
            .O(N__23474),
            .I(N__23438));
    LocalMux I__5588 (
            .O(N__23471),
            .I(N__23435));
    InMux I__5587 (
            .O(N__23470),
            .I(N__23432));
    Span4Mux_v I__5586 (
            .O(N__23467),
            .I(N__23425));
    LocalMux I__5585 (
            .O(N__23456),
            .I(N__23425));
    LocalMux I__5584 (
            .O(N__23453),
            .I(N__23422));
    LocalMux I__5583 (
            .O(N__23450),
            .I(N__23415));
    Span4Mux_h I__5582 (
            .O(N__23447),
            .I(N__23415));
    Span4Mux_h I__5581 (
            .O(N__23444),
            .I(N__23415));
    Sp12to4 I__5580 (
            .O(N__23441),
            .I(N__23408));
    Span12Mux_h I__5579 (
            .O(N__23438),
            .I(N__23408));
    Span12Mux_s2_h I__5578 (
            .O(N__23435),
            .I(N__23408));
    LocalMux I__5577 (
            .O(N__23432),
            .I(N__23404));
    InMux I__5576 (
            .O(N__23431),
            .I(N__23401));
    InMux I__5575 (
            .O(N__23430),
            .I(N__23398));
    Span4Mux_v I__5574 (
            .O(N__23425),
            .I(N__23395));
    Span12Mux_h I__5573 (
            .O(N__23422),
            .I(N__23392));
    Span4Mux_v I__5572 (
            .O(N__23415),
            .I(N__23389));
    Span12Mux_h I__5571 (
            .O(N__23408),
            .I(N__23386));
    InMux I__5570 (
            .O(N__23407),
            .I(N__23383));
    Span12Mux_v I__5569 (
            .O(N__23404),
            .I(N__23380));
    LocalMux I__5568 (
            .O(N__23401),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__5567 (
            .O(N__23398),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__5566 (
            .O(N__23395),
            .I(M_this_state_qZ0Z_3));
    Odrv12 I__5565 (
            .O(N__23392),
            .I(M_this_state_qZ0Z_3));
    Odrv4 I__5564 (
            .O(N__23389),
            .I(M_this_state_qZ0Z_3));
    Odrv12 I__5563 (
            .O(N__23386),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__5562 (
            .O(N__23383),
            .I(M_this_state_qZ0Z_3));
    Odrv12 I__5561 (
            .O(N__23380),
            .I(M_this_state_qZ0Z_3));
    IoInMux I__5560 (
            .O(N__23363),
            .I(N__23360));
    LocalMux I__5559 (
            .O(N__23360),
            .I(N__23357));
    IoSpan4Mux I__5558 (
            .O(N__23357),
            .I(N__23354));
    Span4Mux_s1_v I__5557 (
            .O(N__23354),
            .I(N__23351));
    Sp12to4 I__5556 (
            .O(N__23351),
            .I(N__23348));
    Span12Mux_h I__5555 (
            .O(N__23348),
            .I(N__23344));
    InMux I__5554 (
            .O(N__23347),
            .I(N__23341));
    Odrv12 I__5553 (
            .O(N__23344),
            .I(M_this_external_address_qZ0Z_0));
    LocalMux I__5552 (
            .O(N__23341),
            .I(M_this_external_address_qZ0Z_0));
    IoInMux I__5551 (
            .O(N__23336),
            .I(N__23333));
    LocalMux I__5550 (
            .O(N__23333),
            .I(N__23330));
    Span12Mux_s9_v I__5549 (
            .O(N__23330),
            .I(N__23326));
    InMux I__5548 (
            .O(N__23329),
            .I(N__23323));
    Odrv12 I__5547 (
            .O(N__23326),
            .I(M_this_external_address_qZ0Z_1));
    LocalMux I__5546 (
            .O(N__23323),
            .I(M_this_external_address_qZ0Z_1));
    InMux I__5545 (
            .O(N__23318),
            .I(un1_M_this_external_address_q_cry_0));
    IoInMux I__5544 (
            .O(N__23315),
            .I(N__23312));
    LocalMux I__5543 (
            .O(N__23312),
            .I(N__23309));
    Span4Mux_s3_v I__5542 (
            .O(N__23309),
            .I(N__23306));
    Span4Mux_v I__5541 (
            .O(N__23306),
            .I(N__23303));
    Sp12to4 I__5540 (
            .O(N__23303),
            .I(N__23300));
    Span12Mux_h I__5539 (
            .O(N__23300),
            .I(N__23296));
    InMux I__5538 (
            .O(N__23299),
            .I(N__23293));
    Odrv12 I__5537 (
            .O(N__23296),
            .I(M_this_external_address_qZ0Z_2));
    LocalMux I__5536 (
            .O(N__23293),
            .I(M_this_external_address_qZ0Z_2));
    InMux I__5535 (
            .O(N__23288),
            .I(un1_M_this_external_address_q_cry_1));
    IoInMux I__5534 (
            .O(N__23285),
            .I(N__23282));
    LocalMux I__5533 (
            .O(N__23282),
            .I(N__23279));
    Span4Mux_s1_h I__5532 (
            .O(N__23279),
            .I(N__23276));
    Span4Mux_v I__5531 (
            .O(N__23276),
            .I(N__23272));
    InMux I__5530 (
            .O(N__23275),
            .I(N__23269));
    Odrv4 I__5529 (
            .O(N__23272),
            .I(M_this_external_address_qZ0Z_3));
    LocalMux I__5528 (
            .O(N__23269),
            .I(M_this_external_address_qZ0Z_3));
    InMux I__5527 (
            .O(N__23264),
            .I(un1_M_this_external_address_q_cry_2));
    IoInMux I__5526 (
            .O(N__23261),
            .I(N__23258));
    LocalMux I__5525 (
            .O(N__23258),
            .I(N__23254));
    InMux I__5524 (
            .O(N__23257),
            .I(N__23251));
    Odrv4 I__5523 (
            .O(N__23254),
            .I(M_this_external_address_qZ0Z_4));
    LocalMux I__5522 (
            .O(N__23251),
            .I(M_this_external_address_qZ0Z_4));
    InMux I__5521 (
            .O(N__23246),
            .I(N__23243));
    LocalMux I__5520 (
            .O(N__23243),
            .I(N__23240));
    Span4Mux_v I__5519 (
            .O(N__23240),
            .I(N__23237));
    Span4Mux_v I__5518 (
            .O(N__23237),
            .I(N__23234));
    Span4Mux_v I__5517 (
            .O(N__23234),
            .I(N__23231));
    Odrv4 I__5516 (
            .O(N__23231),
            .I(\this_sprites_ram.mem_out_bus7_3 ));
    InMux I__5515 (
            .O(N__23228),
            .I(N__23225));
    LocalMux I__5514 (
            .O(N__23225),
            .I(N__23222));
    Odrv4 I__5513 (
            .O(N__23222),
            .I(\this_sprites_ram.mem_out_bus3_3 ));
    InMux I__5512 (
            .O(N__23219),
            .I(N__23216));
    LocalMux I__5511 (
            .O(N__23216),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ));
    CEMux I__5510 (
            .O(N__23213),
            .I(N__23210));
    LocalMux I__5509 (
            .O(N__23210),
            .I(N__23206));
    CEMux I__5508 (
            .O(N__23209),
            .I(N__23203));
    Odrv4 I__5507 (
            .O(N__23206),
            .I(\this_sprites_ram.mem_WE_6 ));
    LocalMux I__5506 (
            .O(N__23203),
            .I(\this_sprites_ram.mem_WE_6 ));
    CascadeMux I__5505 (
            .O(N__23198),
            .I(N__23195));
    InMux I__5504 (
            .O(N__23195),
            .I(N__23189));
    CascadeMux I__5503 (
            .O(N__23194),
            .I(N__23186));
    InMux I__5502 (
            .O(N__23193),
            .I(N__23183));
    InMux I__5501 (
            .O(N__23192),
            .I(N__23180));
    LocalMux I__5500 (
            .O(N__23189),
            .I(N__23177));
    InMux I__5499 (
            .O(N__23186),
            .I(N__23174));
    LocalMux I__5498 (
            .O(N__23183),
            .I(N__23171));
    LocalMux I__5497 (
            .O(N__23180),
            .I(N__23168));
    Span4Mux_h I__5496 (
            .O(N__23177),
            .I(N__23163));
    LocalMux I__5495 (
            .O(N__23174),
            .I(N__23163));
    Span4Mux_h I__5494 (
            .O(N__23171),
            .I(N__23160));
    Span4Mux_v I__5493 (
            .O(N__23168),
            .I(N__23157));
    Sp12to4 I__5492 (
            .O(N__23163),
            .I(N__23154));
    Span4Mux_h I__5491 (
            .O(N__23160),
            .I(N__23151));
    Span4Mux_h I__5490 (
            .O(N__23157),
            .I(N__23148));
    Span12Mux_v I__5489 (
            .O(N__23154),
            .I(N__23145));
    Sp12to4 I__5488 (
            .O(N__23151),
            .I(N__23140));
    Sp12to4 I__5487 (
            .O(N__23148),
            .I(N__23140));
    Span12Mux_h I__5486 (
            .O(N__23145),
            .I(N__23137));
    Span12Mux_v I__5485 (
            .O(N__23140),
            .I(N__23134));
    Odrv12 I__5484 (
            .O(N__23137),
            .I(port_data_c_3));
    Odrv12 I__5483 (
            .O(N__23134),
            .I(port_data_c_3));
    CascadeMux I__5482 (
            .O(N__23129),
            .I(N__23126));
    InMux I__5481 (
            .O(N__23126),
            .I(N__23123));
    LocalMux I__5480 (
            .O(N__23123),
            .I(N__23120));
    Span4Mux_v I__5479 (
            .O(N__23120),
            .I(N__23117));
    Span4Mux_h I__5478 (
            .O(N__23117),
            .I(N__23114));
    IoSpan4Mux I__5477 (
            .O(N__23114),
            .I(N__23111));
    Odrv4 I__5476 (
            .O(N__23111),
            .I(port_data_c_7));
    InMux I__5475 (
            .O(N__23108),
            .I(N__23104));
    InMux I__5474 (
            .O(N__23107),
            .I(N__23100));
    LocalMux I__5473 (
            .O(N__23104),
            .I(N__23096));
    InMux I__5472 (
            .O(N__23103),
            .I(N__23093));
    LocalMux I__5471 (
            .O(N__23100),
            .I(N__23089));
    InMux I__5470 (
            .O(N__23099),
            .I(N__23086));
    Span4Mux_v I__5469 (
            .O(N__23096),
            .I(N__23080));
    LocalMux I__5468 (
            .O(N__23093),
            .I(N__23080));
    InMux I__5467 (
            .O(N__23092),
            .I(N__23077));
    Span4Mux_v I__5466 (
            .O(N__23089),
            .I(N__23071));
    LocalMux I__5465 (
            .O(N__23086),
            .I(N__23071));
    InMux I__5464 (
            .O(N__23085),
            .I(N__23068));
    Span4Mux_v I__5463 (
            .O(N__23080),
            .I(N__23062));
    LocalMux I__5462 (
            .O(N__23077),
            .I(N__23062));
    InMux I__5461 (
            .O(N__23076),
            .I(N__23059));
    Span4Mux_v I__5460 (
            .O(N__23071),
            .I(N__23054));
    LocalMux I__5459 (
            .O(N__23068),
            .I(N__23054));
    InMux I__5458 (
            .O(N__23067),
            .I(N__23051));
    Span4Mux_v I__5457 (
            .O(N__23062),
            .I(N__23046));
    LocalMux I__5456 (
            .O(N__23059),
            .I(N__23046));
    Span4Mux_v I__5455 (
            .O(N__23054),
            .I(N__23041));
    LocalMux I__5454 (
            .O(N__23051),
            .I(N__23041));
    Odrv4 I__5453 (
            .O(N__23046),
            .I(M_this_sprites_ram_write_data_3));
    Odrv4 I__5452 (
            .O(N__23041),
            .I(M_this_sprites_ram_write_data_3));
    InMux I__5451 (
            .O(N__23036),
            .I(N__23033));
    LocalMux I__5450 (
            .O(N__23033),
            .I(N__23030));
    Span4Mux_v I__5449 (
            .O(N__23030),
            .I(N__23027));
    Odrv4 I__5448 (
            .O(N__23027),
            .I(\this_sprites_ram.mem_out_bus5_3 ));
    InMux I__5447 (
            .O(N__23024),
            .I(N__23021));
    LocalMux I__5446 (
            .O(N__23021),
            .I(N__23018));
    Span4Mux_v I__5445 (
            .O(N__23018),
            .I(N__23015));
    Span4Mux_v I__5444 (
            .O(N__23015),
            .I(N__23012));
    Odrv4 I__5443 (
            .O(N__23012),
            .I(\this_sprites_ram.mem_out_bus1_3 ));
    InMux I__5442 (
            .O(N__23009),
            .I(N__23006));
    LocalMux I__5441 (
            .O(N__23006),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ));
    InMux I__5440 (
            .O(N__23003),
            .I(N__23000));
    LocalMux I__5439 (
            .O(N__23000),
            .I(N__22997));
    Sp12to4 I__5438 (
            .O(N__22997),
            .I(N__22994));
    Span12Mux_v I__5437 (
            .O(N__22994),
            .I(N__22991));
    Odrv12 I__5436 (
            .O(N__22991),
            .I(\this_sprites_ram.mem_out_bus0_3 ));
    InMux I__5435 (
            .O(N__22988),
            .I(N__22985));
    LocalMux I__5434 (
            .O(N__22985),
            .I(\this_sprites_ram.mem_out_bus4_3 ));
    InMux I__5433 (
            .O(N__22982),
            .I(N__22979));
    LocalMux I__5432 (
            .O(N__22979),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ));
    InMux I__5431 (
            .O(N__22976),
            .I(N__22973));
    LocalMux I__5430 (
            .O(N__22973),
            .I(N__22970));
    Sp12to4 I__5429 (
            .O(N__22970),
            .I(N__22967));
    Odrv12 I__5428 (
            .O(N__22967),
            .I(\this_sprites_ram.mem_out_bus6_3 ));
    InMux I__5427 (
            .O(N__22964),
            .I(N__22961));
    LocalMux I__5426 (
            .O(N__22961),
            .I(N__22958));
    Span4Mux_v I__5425 (
            .O(N__22958),
            .I(N__22955));
    Span4Mux_v I__5424 (
            .O(N__22955),
            .I(N__22952));
    Odrv4 I__5423 (
            .O(N__22952),
            .I(\this_sprites_ram.mem_out_bus2_3 ));
    InMux I__5422 (
            .O(N__22949),
            .I(N__22946));
    LocalMux I__5421 (
            .O(N__22946),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ));
    InMux I__5420 (
            .O(N__22943),
            .I(N__22940));
    LocalMux I__5419 (
            .O(N__22940),
            .I(N__22937));
    Span4Mux_v I__5418 (
            .O(N__22937),
            .I(N__22934));
    Span4Mux_v I__5417 (
            .O(N__22934),
            .I(N__22931));
    Odrv4 I__5416 (
            .O(N__22931),
            .I(\this_sprites_ram.mem_out_bus7_0 ));
    InMux I__5415 (
            .O(N__22928),
            .I(N__22925));
    LocalMux I__5414 (
            .O(N__22925),
            .I(N__22922));
    Span4Mux_v I__5413 (
            .O(N__22922),
            .I(N__22919));
    Odrv4 I__5412 (
            .O(N__22919),
            .I(\this_sprites_ram.mem_out_bus3_0 ));
    InMux I__5411 (
            .O(N__22916),
            .I(N__22911));
    InMux I__5410 (
            .O(N__22915),
            .I(N__22899));
    InMux I__5409 (
            .O(N__22914),
            .I(N__22899));
    LocalMux I__5408 (
            .O(N__22911),
            .I(N__22891));
    InMux I__5407 (
            .O(N__22910),
            .I(N__22888));
    InMux I__5406 (
            .O(N__22909),
            .I(N__22883));
    InMux I__5405 (
            .O(N__22908),
            .I(N__22883));
    InMux I__5404 (
            .O(N__22907),
            .I(N__22880));
    InMux I__5403 (
            .O(N__22906),
            .I(N__22873));
    InMux I__5402 (
            .O(N__22905),
            .I(N__22873));
    InMux I__5401 (
            .O(N__22904),
            .I(N__22873));
    LocalMux I__5400 (
            .O(N__22899),
            .I(N__22870));
    InMux I__5399 (
            .O(N__22898),
            .I(N__22867));
    InMux I__5398 (
            .O(N__22897),
            .I(N__22862));
    InMux I__5397 (
            .O(N__22896),
            .I(N__22862));
    InMux I__5396 (
            .O(N__22895),
            .I(N__22859));
    InMux I__5395 (
            .O(N__22894),
            .I(N__22856));
    Span4Mux_v I__5394 (
            .O(N__22891),
            .I(N__22850));
    LocalMux I__5393 (
            .O(N__22888),
            .I(N__22850));
    LocalMux I__5392 (
            .O(N__22883),
            .I(N__22841));
    LocalMux I__5391 (
            .O(N__22880),
            .I(N__22841));
    LocalMux I__5390 (
            .O(N__22873),
            .I(N__22841));
    Span4Mux_h I__5389 (
            .O(N__22870),
            .I(N__22841));
    LocalMux I__5388 (
            .O(N__22867),
            .I(N__22832));
    LocalMux I__5387 (
            .O(N__22862),
            .I(N__22832));
    LocalMux I__5386 (
            .O(N__22859),
            .I(N__22832));
    LocalMux I__5385 (
            .O(N__22856),
            .I(N__22832));
    InMux I__5384 (
            .O(N__22855),
            .I(N__22829));
    Span4Mux_h I__5383 (
            .O(N__22850),
            .I(N__22826));
    Span4Mux_v I__5382 (
            .O(N__22841),
            .I(N__22819));
    Span4Mux_v I__5381 (
            .O(N__22832),
            .I(N__22819));
    LocalMux I__5380 (
            .O(N__22829),
            .I(N__22819));
    Span4Mux_v I__5379 (
            .O(N__22826),
            .I(N__22814));
    Span4Mux_h I__5378 (
            .O(N__22819),
            .I(N__22814));
    Odrv4 I__5377 (
            .O(N__22814),
            .I(\this_sprites_ram.mem_radregZ0Z_13 ));
    InMux I__5376 (
            .O(N__22811),
            .I(N__22808));
    LocalMux I__5375 (
            .O(N__22808),
            .I(N__22805));
    Span12Mux_h I__5374 (
            .O(N__22805),
            .I(N__22802));
    Odrv12 I__5373 (
            .O(N__22802),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ));
    InMux I__5372 (
            .O(N__22799),
            .I(N__22796));
    LocalMux I__5371 (
            .O(N__22796),
            .I(N__22792));
    InMux I__5370 (
            .O(N__22795),
            .I(N__22789));
    Span4Mux_v I__5369 (
            .O(N__22792),
            .I(N__22783));
    LocalMux I__5368 (
            .O(N__22789),
            .I(N__22783));
    InMux I__5367 (
            .O(N__22788),
            .I(N__22780));
    Span4Mux_h I__5366 (
            .O(N__22783),
            .I(N__22774));
    LocalMux I__5365 (
            .O(N__22780),
            .I(N__22774));
    InMux I__5364 (
            .O(N__22779),
            .I(N__22771));
    Odrv4 I__5363 (
            .O(N__22774),
            .I(\this_vga_signals.N_481 ));
    LocalMux I__5362 (
            .O(N__22771),
            .I(\this_vga_signals.N_481 ));
    CascadeMux I__5361 (
            .O(N__22766),
            .I(N__22763));
    InMux I__5360 (
            .O(N__22763),
            .I(N__22760));
    LocalMux I__5359 (
            .O(N__22760),
            .I(N__22756));
    CascadeMux I__5358 (
            .O(N__22759),
            .I(N__22751));
    Span4Mux_h I__5357 (
            .O(N__22756),
            .I(N__22748));
    InMux I__5356 (
            .O(N__22755),
            .I(N__22745));
    InMux I__5355 (
            .O(N__22754),
            .I(N__22740));
    InMux I__5354 (
            .O(N__22751),
            .I(N__22740));
    Span4Mux_v I__5353 (
            .O(N__22748),
            .I(N__22735));
    LocalMux I__5352 (
            .O(N__22745),
            .I(N__22735));
    LocalMux I__5351 (
            .O(N__22740),
            .I(N__22732));
    Span4Mux_v I__5350 (
            .O(N__22735),
            .I(N__22729));
    Span12Mux_v I__5349 (
            .O(N__22732),
            .I(N__22726));
    Sp12to4 I__5348 (
            .O(N__22729),
            .I(N__22723));
    Span12Mux_h I__5347 (
            .O(N__22726),
            .I(N__22720));
    Span12Mux_h I__5346 (
            .O(N__22723),
            .I(N__22717));
    Odrv12 I__5345 (
            .O(N__22720),
            .I(port_data_c_2));
    Odrv12 I__5344 (
            .O(N__22717),
            .I(port_data_c_2));
    CascadeMux I__5343 (
            .O(N__22712),
            .I(N__22708));
    InMux I__5342 (
            .O(N__22711),
            .I(N__22703));
    InMux I__5341 (
            .O(N__22708),
            .I(N__22703));
    LocalMux I__5340 (
            .O(N__22703),
            .I(N__22700));
    Span4Mux_v I__5339 (
            .O(N__22700),
            .I(N__22696));
    CascadeMux I__5338 (
            .O(N__22699),
            .I(N__22693));
    Span4Mux_h I__5337 (
            .O(N__22696),
            .I(N__22690));
    InMux I__5336 (
            .O(N__22693),
            .I(N__22687));
    Sp12to4 I__5335 (
            .O(N__22690),
            .I(N__22682));
    LocalMux I__5334 (
            .O(N__22687),
            .I(N__22682));
    Span12Mux_v I__5333 (
            .O(N__22682),
            .I(N__22679));
    Odrv12 I__5332 (
            .O(N__22679),
            .I(port_data_c_6));
    CEMux I__5331 (
            .O(N__22676),
            .I(N__22672));
    CEMux I__5330 (
            .O(N__22675),
            .I(N__22669));
    LocalMux I__5329 (
            .O(N__22672),
            .I(N__22664));
    LocalMux I__5328 (
            .O(N__22669),
            .I(N__22664));
    Odrv4 I__5327 (
            .O(N__22664),
            .I(\this_sprites_ram.mem_WE_10 ));
    CEMux I__5326 (
            .O(N__22661),
            .I(N__22657));
    CEMux I__5325 (
            .O(N__22660),
            .I(N__22654));
    LocalMux I__5324 (
            .O(N__22657),
            .I(N__22651));
    LocalMux I__5323 (
            .O(N__22654),
            .I(N__22648));
    Span4Mux_v I__5322 (
            .O(N__22651),
            .I(N__22645));
    Span4Mux_h I__5321 (
            .O(N__22648),
            .I(N__22642));
    Odrv4 I__5320 (
            .O(N__22645),
            .I(\this_sprites_ram.mem_WE_12 ));
    Odrv4 I__5319 (
            .O(N__22642),
            .I(\this_sprites_ram.mem_WE_12 ));
    InMux I__5318 (
            .O(N__22637),
            .I(N__22634));
    LocalMux I__5317 (
            .O(N__22634),
            .I(N__22631));
    Span4Mux_v I__5316 (
            .O(N__22631),
            .I(N__22628));
    Sp12to4 I__5315 (
            .O(N__22628),
            .I(N__22625));
    Odrv12 I__5314 (
            .O(N__22625),
            .I(\this_sprites_ram.mem_out_bus5_2 ));
    InMux I__5313 (
            .O(N__22622),
            .I(N__22619));
    LocalMux I__5312 (
            .O(N__22619),
            .I(N__22616));
    Span4Mux_v I__5311 (
            .O(N__22616),
            .I(N__22613));
    Odrv4 I__5310 (
            .O(N__22613),
            .I(\this_sprites_ram.mem_out_bus1_2 ));
    InMux I__5309 (
            .O(N__22610),
            .I(N__22607));
    LocalMux I__5308 (
            .O(N__22607),
            .I(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ));
    InMux I__5307 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__5306 (
            .O(N__22601),
            .I(N__22598));
    Span4Mux_h I__5305 (
            .O(N__22598),
            .I(N__22595));
    Odrv4 I__5304 (
            .O(N__22595),
            .I(\this_sprites_ram.mem_out_bus4_1 ));
    InMux I__5303 (
            .O(N__22592),
            .I(N__22589));
    LocalMux I__5302 (
            .O(N__22589),
            .I(N__22586));
    Sp12to4 I__5301 (
            .O(N__22586),
            .I(N__22583));
    Span12Mux_v I__5300 (
            .O(N__22583),
            .I(N__22580));
    Odrv12 I__5299 (
            .O(N__22580),
            .I(\this_sprites_ram.mem_out_bus0_1 ));
    InMux I__5298 (
            .O(N__22577),
            .I(N__22574));
    LocalMux I__5297 (
            .O(N__22574),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ));
    InMux I__5296 (
            .O(N__22571),
            .I(N__22568));
    LocalMux I__5295 (
            .O(N__22568),
            .I(N__22565));
    Span4Mux_v I__5294 (
            .O(N__22565),
            .I(N__22562));
    Odrv4 I__5293 (
            .O(N__22562),
            .I(\this_sprites_ram.mem_out_bus4_2 ));
    InMux I__5292 (
            .O(N__22559),
            .I(N__22556));
    LocalMux I__5291 (
            .O(N__22556),
            .I(N__22553));
    Span4Mux_v I__5290 (
            .O(N__22553),
            .I(N__22550));
    Span4Mux_v I__5289 (
            .O(N__22550),
            .I(N__22547));
    Odrv4 I__5288 (
            .O(N__22547),
            .I(\this_sprites_ram.mem_out_bus0_2 ));
    InMux I__5287 (
            .O(N__22544),
            .I(N__22541));
    LocalMux I__5286 (
            .O(N__22541),
            .I(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0 ));
    CEMux I__5285 (
            .O(N__22538),
            .I(N__22534));
    CEMux I__5284 (
            .O(N__22537),
            .I(N__22531));
    LocalMux I__5283 (
            .O(N__22534),
            .I(N__22528));
    LocalMux I__5282 (
            .O(N__22531),
            .I(N__22525));
    Span4Mux_v I__5281 (
            .O(N__22528),
            .I(N__22522));
    Span4Mux_h I__5280 (
            .O(N__22525),
            .I(N__22519));
    Odrv4 I__5279 (
            .O(N__22522),
            .I(\this_sprites_ram.mem_WE_8 ));
    Odrv4 I__5278 (
            .O(N__22519),
            .I(\this_sprites_ram.mem_WE_8 ));
    InMux I__5277 (
            .O(N__22514),
            .I(N__22511));
    LocalMux I__5276 (
            .O(N__22511),
            .I(N__22508));
    Sp12to4 I__5275 (
            .O(N__22508),
            .I(N__22505));
    Span12Mux_v I__5274 (
            .O(N__22505),
            .I(N__22502));
    Span12Mux_v I__5273 (
            .O(N__22502),
            .I(N__22499));
    Odrv12 I__5272 (
            .O(N__22499),
            .I(\this_sprites_ram.mem_out_bus7_2 ));
    InMux I__5271 (
            .O(N__22496),
            .I(N__22493));
    LocalMux I__5270 (
            .O(N__22493),
            .I(N__22490));
    Span4Mux_h I__5269 (
            .O(N__22490),
            .I(N__22487));
    Odrv4 I__5268 (
            .O(N__22487),
            .I(\this_sprites_ram.mem_out_bus3_2 ));
    InMux I__5267 (
            .O(N__22484),
            .I(N__22481));
    LocalMux I__5266 (
            .O(N__22481),
            .I(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ));
    InMux I__5265 (
            .O(N__22478),
            .I(N__22475));
    LocalMux I__5264 (
            .O(N__22475),
            .I(N__22472));
    Span4Mux_v I__5263 (
            .O(N__22472),
            .I(N__22469));
    Span4Mux_v I__5262 (
            .O(N__22469),
            .I(N__22466));
    Span4Mux_v I__5261 (
            .O(N__22466),
            .I(N__22463));
    Odrv4 I__5260 (
            .O(N__22463),
            .I(\this_sprites_ram.mem_out_bus7_1 ));
    InMux I__5259 (
            .O(N__22460),
            .I(N__22457));
    LocalMux I__5258 (
            .O(N__22457),
            .I(\this_sprites_ram.mem_out_bus3_1 ));
    InMux I__5257 (
            .O(N__22454),
            .I(N__22451));
    LocalMux I__5256 (
            .O(N__22451),
            .I(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ));
    InMux I__5255 (
            .O(N__22448),
            .I(N__22445));
    LocalMux I__5254 (
            .O(N__22445),
            .I(N__22442));
    Span4Mux_v I__5253 (
            .O(N__22442),
            .I(N__22439));
    Span4Mux_v I__5252 (
            .O(N__22439),
            .I(N__22436));
    Odrv4 I__5251 (
            .O(N__22436),
            .I(\this_sprites_ram.mem_out_bus6_1 ));
    InMux I__5250 (
            .O(N__22433),
            .I(N__22430));
    LocalMux I__5249 (
            .O(N__22430),
            .I(N__22427));
    Span4Mux_v I__5248 (
            .O(N__22427),
            .I(N__22424));
    Odrv4 I__5247 (
            .O(N__22424),
            .I(\this_sprites_ram.mem_out_bus2_1 ));
    InMux I__5246 (
            .O(N__22421),
            .I(N__22418));
    LocalMux I__5245 (
            .O(N__22418),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ));
    CascadeMux I__5244 (
            .O(N__22415),
            .I(M_this_sprites_ram_read_data_3_cascade_));
    InMux I__5243 (
            .O(N__22412),
            .I(N__22408));
    InMux I__5242 (
            .O(N__22411),
            .I(N__22405));
    LocalMux I__5241 (
            .O(N__22408),
            .I(N__22401));
    LocalMux I__5240 (
            .O(N__22405),
            .I(N__22398));
    InMux I__5239 (
            .O(N__22404),
            .I(N__22395));
    Span4Mux_h I__5238 (
            .O(N__22401),
            .I(N__22392));
    Span4Mux_h I__5237 (
            .O(N__22398),
            .I(N__22387));
    LocalMux I__5236 (
            .O(N__22395),
            .I(N__22387));
    Span4Mux_h I__5235 (
            .O(N__22392),
            .I(N__22379));
    Span4Mux_v I__5234 (
            .O(N__22387),
            .I(N__22379));
    InMux I__5233 (
            .O(N__22386),
            .I(N__22375));
    InMux I__5232 (
            .O(N__22385),
            .I(N__22372));
    InMux I__5231 (
            .O(N__22384),
            .I(N__22369));
    Span4Mux_h I__5230 (
            .O(N__22379),
            .I(N__22366));
    CascadeMux I__5229 (
            .O(N__22378),
            .I(N__22360));
    LocalMux I__5228 (
            .O(N__22375),
            .I(N__22357));
    LocalMux I__5227 (
            .O(N__22372),
            .I(N__22354));
    LocalMux I__5226 (
            .O(N__22369),
            .I(N__22351));
    Span4Mux_h I__5225 (
            .O(N__22366),
            .I(N__22348));
    InMux I__5224 (
            .O(N__22365),
            .I(N__22341));
    InMux I__5223 (
            .O(N__22364),
            .I(N__22341));
    InMux I__5222 (
            .O(N__22363),
            .I(N__22341));
    InMux I__5221 (
            .O(N__22360),
            .I(N__22338));
    Span4Mux_h I__5220 (
            .O(N__22357),
            .I(N__22331));
    Span4Mux_v I__5219 (
            .O(N__22354),
            .I(N__22331));
    Span4Mux_h I__5218 (
            .O(N__22351),
            .I(N__22331));
    Odrv4 I__5217 (
            .O(N__22348),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__5216 (
            .O(N__22341),
            .I(M_this_ppu_vram_en_0));
    LocalMux I__5215 (
            .O(N__22338),
            .I(M_this_ppu_vram_en_0));
    Odrv4 I__5214 (
            .O(N__22331),
            .I(M_this_ppu_vram_en_0));
    InMux I__5213 (
            .O(N__22322),
            .I(N__22319));
    LocalMux I__5212 (
            .O(N__22319),
            .I(N__22316));
    Span4Mux_v I__5211 (
            .O(N__22316),
            .I(N__22313));
    Span4Mux_h I__5210 (
            .O(N__22313),
            .I(N__22310));
    Sp12to4 I__5209 (
            .O(N__22310),
            .I(N__22307));
    Span12Mux_h I__5208 (
            .O(N__22307),
            .I(N__22304));
    Odrv12 I__5207 (
            .O(N__22304),
            .I(M_this_vram_write_data_3));
    CascadeMux I__5206 (
            .O(N__22301),
            .I(N__22295));
    CascadeMux I__5205 (
            .O(N__22300),
            .I(N__22292));
    InMux I__5204 (
            .O(N__22299),
            .I(N__22289));
    InMux I__5203 (
            .O(N__22298),
            .I(N__22286));
    InMux I__5202 (
            .O(N__22295),
            .I(N__22282));
    InMux I__5201 (
            .O(N__22292),
            .I(N__22279));
    LocalMux I__5200 (
            .O(N__22289),
            .I(N__22274));
    LocalMux I__5199 (
            .O(N__22286),
            .I(N__22274));
    InMux I__5198 (
            .O(N__22285),
            .I(N__22271));
    LocalMux I__5197 (
            .O(N__22282),
            .I(N__22265));
    LocalMux I__5196 (
            .O(N__22279),
            .I(N__22260));
    Span4Mux_h I__5195 (
            .O(N__22274),
            .I(N__22260));
    LocalMux I__5194 (
            .O(N__22271),
            .I(N__22257));
    InMux I__5193 (
            .O(N__22270),
            .I(N__22254));
    InMux I__5192 (
            .O(N__22269),
            .I(N__22251));
    InMux I__5191 (
            .O(N__22268),
            .I(N__22248));
    Span4Mux_v I__5190 (
            .O(N__22265),
            .I(N__22245));
    Span4Mux_v I__5189 (
            .O(N__22260),
            .I(N__22238));
    Span4Mux_h I__5188 (
            .O(N__22257),
            .I(N__22238));
    LocalMux I__5187 (
            .O(N__22254),
            .I(N__22238));
    LocalMux I__5186 (
            .O(N__22251),
            .I(N__22233));
    LocalMux I__5185 (
            .O(N__22248),
            .I(N__22233));
    Span4Mux_h I__5184 (
            .O(N__22245),
            .I(N__22228));
    Span4Mux_h I__5183 (
            .O(N__22238),
            .I(N__22228));
    Span12Mux_h I__5182 (
            .O(N__22233),
            .I(N__22225));
    Span4Mux_h I__5181 (
            .O(N__22228),
            .I(N__22222));
    Odrv12 I__5180 (
            .O(N__22225),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    Odrv4 I__5179 (
            .O(N__22222),
            .I(\this_sprites_ram.mem_radregZ0Z_11 ));
    CascadeMux I__5178 (
            .O(N__22217),
            .I(N__22214));
    InMux I__5177 (
            .O(N__22214),
            .I(N__22208));
    CascadeMux I__5176 (
            .O(N__22213),
            .I(N__22205));
    CascadeMux I__5175 (
            .O(N__22212),
            .I(N__22202));
    InMux I__5174 (
            .O(N__22211),
            .I(N__22199));
    LocalMux I__5173 (
            .O(N__22208),
            .I(N__22196));
    InMux I__5172 (
            .O(N__22205),
            .I(N__22193));
    InMux I__5171 (
            .O(N__22202),
            .I(N__22190));
    LocalMux I__5170 (
            .O(N__22199),
            .I(N__22187));
    Span4Mux_v I__5169 (
            .O(N__22196),
            .I(N__22182));
    LocalMux I__5168 (
            .O(N__22193),
            .I(N__22182));
    LocalMux I__5167 (
            .O(N__22190),
            .I(N__22179));
    Span4Mux_h I__5166 (
            .O(N__22187),
            .I(N__22176));
    Span4Mux_v I__5165 (
            .O(N__22182),
            .I(N__22173));
    Span4Mux_v I__5164 (
            .O(N__22179),
            .I(N__22170));
    Span4Mux_v I__5163 (
            .O(N__22176),
            .I(N__22165));
    Span4Mux_h I__5162 (
            .O(N__22173),
            .I(N__22165));
    Span4Mux_h I__5161 (
            .O(N__22170),
            .I(N__22162));
    Odrv4 I__5160 (
            .O(N__22165),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    Odrv4 I__5159 (
            .O(N__22162),
            .I(\this_sprites_ram.mem_radregZ0Z_12 ));
    InMux I__5158 (
            .O(N__22157),
            .I(N__22154));
    LocalMux I__5157 (
            .O(N__22154),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3 ));
    InMux I__5156 (
            .O(N__22151),
            .I(N__22148));
    LocalMux I__5155 (
            .O(N__22148),
            .I(N__22145));
    Span12Mux_h I__5154 (
            .O(N__22145),
            .I(N__22142));
    Odrv12 I__5153 (
            .O(N__22142),
            .I(\this_sprites_ram.mem_out_bus6_0 ));
    InMux I__5152 (
            .O(N__22139),
            .I(N__22136));
    LocalMux I__5151 (
            .O(N__22136),
            .I(N__22133));
    Span4Mux_v I__5150 (
            .O(N__22133),
            .I(N__22130));
    Span4Mux_v I__5149 (
            .O(N__22130),
            .I(N__22127));
    Odrv4 I__5148 (
            .O(N__22127),
            .I(\this_sprites_ram.mem_out_bus2_0 ));
    InMux I__5147 (
            .O(N__22124),
            .I(N__22121));
    LocalMux I__5146 (
            .O(N__22121),
            .I(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ));
    InMux I__5145 (
            .O(N__22118),
            .I(N__22115));
    LocalMux I__5144 (
            .O(N__22115),
            .I(N__22112));
    Span4Mux_v I__5143 (
            .O(N__22112),
            .I(N__22109));
    Odrv4 I__5142 (
            .O(N__22109),
            .I(\this_sprites_ram.mem_out_bus5_0 ));
    InMux I__5141 (
            .O(N__22106),
            .I(N__22103));
    LocalMux I__5140 (
            .O(N__22103),
            .I(N__22100));
    Span4Mux_v I__5139 (
            .O(N__22100),
            .I(N__22097));
    Span4Mux_v I__5138 (
            .O(N__22097),
            .I(N__22094));
    Span4Mux_v I__5137 (
            .O(N__22094),
            .I(N__22091));
    Span4Mux_v I__5136 (
            .O(N__22091),
            .I(N__22088));
    Odrv4 I__5135 (
            .O(N__22088),
            .I(\this_sprites_ram.mem_out_bus1_0 ));
    InMux I__5134 (
            .O(N__22085),
            .I(N__22082));
    LocalMux I__5133 (
            .O(N__22082),
            .I(N__22079));
    Span12Mux_h I__5132 (
            .O(N__22079),
            .I(N__22076));
    Odrv12 I__5131 (
            .O(N__22076),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ));
    InMux I__5130 (
            .O(N__22073),
            .I(N__22069));
    InMux I__5129 (
            .O(N__22072),
            .I(N__22066));
    LocalMux I__5128 (
            .O(N__22069),
            .I(N__22063));
    LocalMux I__5127 (
            .O(N__22066),
            .I(N__22060));
    Odrv12 I__5126 (
            .O(N__22063),
            .I(\this_vga_signals.N_483 ));
    Odrv4 I__5125 (
            .O(N__22060),
            .I(\this_vga_signals.N_483 ));
    InMux I__5124 (
            .O(N__22055),
            .I(N__22049));
    InMux I__5123 (
            .O(N__22054),
            .I(N__22046));
    InMux I__5122 (
            .O(N__22053),
            .I(N__22037));
    InMux I__5121 (
            .O(N__22052),
            .I(N__22032));
    LocalMux I__5120 (
            .O(N__22049),
            .I(N__22023));
    LocalMux I__5119 (
            .O(N__22046),
            .I(N__22018));
    InMux I__5118 (
            .O(N__22045),
            .I(N__22011));
    InMux I__5117 (
            .O(N__22044),
            .I(N__22011));
    InMux I__5116 (
            .O(N__22043),
            .I(N__22011));
    InMux I__5115 (
            .O(N__22042),
            .I(N__22004));
    InMux I__5114 (
            .O(N__22041),
            .I(N__22004));
    InMux I__5113 (
            .O(N__22040),
            .I(N__22004));
    LocalMux I__5112 (
            .O(N__22037),
            .I(N__22000));
    InMux I__5111 (
            .O(N__22036),
            .I(N__21995));
    InMux I__5110 (
            .O(N__22035),
            .I(N__21995));
    LocalMux I__5109 (
            .O(N__22032),
            .I(N__21992));
    InMux I__5108 (
            .O(N__22031),
            .I(N__21989));
    InMux I__5107 (
            .O(N__22030),
            .I(N__21986));
    InMux I__5106 (
            .O(N__22029),
            .I(N__21983));
    InMux I__5105 (
            .O(N__22028),
            .I(N__21978));
    InMux I__5104 (
            .O(N__22027),
            .I(N__21978));
    InMux I__5103 (
            .O(N__22026),
            .I(N__21972));
    Span4Mux_v I__5102 (
            .O(N__22023),
            .I(N__21969));
    InMux I__5101 (
            .O(N__22022),
            .I(N__21966));
    InMux I__5100 (
            .O(N__22021),
            .I(N__21963));
    Span4Mux_v I__5099 (
            .O(N__22018),
            .I(N__21956));
    LocalMux I__5098 (
            .O(N__22011),
            .I(N__21956));
    LocalMux I__5097 (
            .O(N__22004),
            .I(N__21956));
    InMux I__5096 (
            .O(N__22003),
            .I(N__21953));
    Sp12to4 I__5095 (
            .O(N__22000),
            .I(N__21948));
    LocalMux I__5094 (
            .O(N__21995),
            .I(N__21948));
    Span4Mux_v I__5093 (
            .O(N__21992),
            .I(N__21939));
    LocalMux I__5092 (
            .O(N__21989),
            .I(N__21939));
    LocalMux I__5091 (
            .O(N__21986),
            .I(N__21939));
    LocalMux I__5090 (
            .O(N__21983),
            .I(N__21939));
    LocalMux I__5089 (
            .O(N__21978),
            .I(N__21936));
    InMux I__5088 (
            .O(N__21977),
            .I(N__21929));
    InMux I__5087 (
            .O(N__21976),
            .I(N__21929));
    InMux I__5086 (
            .O(N__21975),
            .I(N__21929));
    LocalMux I__5085 (
            .O(N__21972),
            .I(N__21922));
    Sp12to4 I__5084 (
            .O(N__21969),
            .I(N__21922));
    LocalMux I__5083 (
            .O(N__21966),
            .I(N__21922));
    LocalMux I__5082 (
            .O(N__21963),
            .I(N__21917));
    Span4Mux_h I__5081 (
            .O(N__21956),
            .I(N__21917));
    LocalMux I__5080 (
            .O(N__21953),
            .I(N__21912));
    Span12Mux_v I__5079 (
            .O(N__21948),
            .I(N__21912));
    Span4Mux_h I__5078 (
            .O(N__21939),
            .I(N__21905));
    Span4Mux_v I__5077 (
            .O(N__21936),
            .I(N__21905));
    LocalMux I__5076 (
            .O(N__21929),
            .I(N__21905));
    Span12Mux_h I__5075 (
            .O(N__21922),
            .I(N__21902));
    Span4Mux_h I__5074 (
            .O(N__21917),
            .I(N__21899));
    Odrv12 I__5073 (
            .O(N__21912),
            .I(N_175_0));
    Odrv4 I__5072 (
            .O(N__21905),
            .I(N_175_0));
    Odrv12 I__5071 (
            .O(N__21902),
            .I(N_175_0));
    Odrv4 I__5070 (
            .O(N__21899),
            .I(N_175_0));
    CEMux I__5069 (
            .O(N__21890),
            .I(N__21887));
    LocalMux I__5068 (
            .O(N__21887),
            .I(N__21883));
    CEMux I__5067 (
            .O(N__21886),
            .I(N__21880));
    Span4Mux_s2_v I__5066 (
            .O(N__21883),
            .I(N__21875));
    LocalMux I__5065 (
            .O(N__21880),
            .I(N__21875));
    Span4Mux_v I__5064 (
            .O(N__21875),
            .I(N__21872));
    Span4Mux_v I__5063 (
            .O(N__21872),
            .I(N__21869));
    Odrv4 I__5062 (
            .O(N__21869),
            .I(\this_sprites_ram.mem_WE_0 ));
    CEMux I__5061 (
            .O(N__21866),
            .I(N__21862));
    CEMux I__5060 (
            .O(N__21865),
            .I(N__21859));
    LocalMux I__5059 (
            .O(N__21862),
            .I(N__21856));
    LocalMux I__5058 (
            .O(N__21859),
            .I(N__21853));
    Span4Mux_s3_v I__5057 (
            .O(N__21856),
            .I(N__21850));
    Span4Mux_h I__5056 (
            .O(N__21853),
            .I(N__21847));
    Span4Mux_v I__5055 (
            .O(N__21850),
            .I(N__21844));
    Span4Mux_v I__5054 (
            .O(N__21847),
            .I(N__21841));
    Odrv4 I__5053 (
            .O(N__21844),
            .I(\this_sprites_ram.mem_WE_14 ));
    Odrv4 I__5052 (
            .O(N__21841),
            .I(\this_sprites_ram.mem_WE_14 ));
    InMux I__5051 (
            .O(N__21836),
            .I(N__21833));
    LocalMux I__5050 (
            .O(N__21833),
            .I(N__21830));
    Span4Mux_v I__5049 (
            .O(N__21830),
            .I(N__21827));
    Span4Mux_h I__5048 (
            .O(N__21827),
            .I(N__21824));
    Sp12to4 I__5047 (
            .O(N__21824),
            .I(N__21821));
    Odrv12 I__5046 (
            .O(N__21821),
            .I(M_this_vram_write_data_2));
    InMux I__5045 (
            .O(N__21818),
            .I(N__21815));
    LocalMux I__5044 (
            .O(N__21815),
            .I(N__21812));
    Span4Mux_v I__5043 (
            .O(N__21812),
            .I(N__21809));
    Span4Mux_h I__5042 (
            .O(N__21809),
            .I(N__21806));
    Span4Mux_h I__5041 (
            .O(N__21806),
            .I(N__21803));
    Odrv4 I__5040 (
            .O(N__21803),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ));
    InMux I__5039 (
            .O(N__21800),
            .I(N__21797));
    LocalMux I__5038 (
            .O(N__21797),
            .I(N__21794));
    Span4Mux_v I__5037 (
            .O(N__21794),
            .I(N__21791));
    Span4Mux_v I__5036 (
            .O(N__21791),
            .I(N__21788));
    Span4Mux_v I__5035 (
            .O(N__21788),
            .I(N__21785));
    Span4Mux_v I__5034 (
            .O(N__21785),
            .I(N__21782));
    Odrv4 I__5033 (
            .O(N__21782),
            .I(\this_sprites_ram.mem_out_bus6_2 ));
    InMux I__5032 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__5031 (
            .O(N__21776),
            .I(N__21773));
    Span4Mux_v I__5030 (
            .O(N__21773),
            .I(N__21770));
    Odrv4 I__5029 (
            .O(N__21770),
            .I(\this_sprites_ram.mem_out_bus2_2 ));
    CascadeMux I__5028 (
            .O(N__21767),
            .I(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_ ));
    CascadeMux I__5027 (
            .O(N__21764),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ));
    InMux I__5026 (
            .O(N__21761),
            .I(N__21758));
    LocalMux I__5025 (
            .O(N__21758),
            .I(M_this_sprites_ram_read_data_2));
    CascadeMux I__5024 (
            .O(N__21755),
            .I(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ));
    InMux I__5023 (
            .O(N__21752),
            .I(N__21749));
    LocalMux I__5022 (
            .O(N__21749),
            .I(N__21746));
    Odrv12 I__5021 (
            .O(N__21746),
            .I(M_this_sprites_ram_read_data_1));
    InMux I__5020 (
            .O(N__21743),
            .I(N__21740));
    LocalMux I__5019 (
            .O(N__21740),
            .I(N__21737));
    Span4Mux_v I__5018 (
            .O(N__21737),
            .I(N__21734));
    Span4Mux_v I__5017 (
            .O(N__21734),
            .I(N__21731));
    Odrv4 I__5016 (
            .O(N__21731),
            .I(\this_sprites_ram.mem_out_bus5_1 ));
    InMux I__5015 (
            .O(N__21728),
            .I(N__21725));
    LocalMux I__5014 (
            .O(N__21725),
            .I(N__21722));
    Span4Mux_v I__5013 (
            .O(N__21722),
            .I(N__21719));
    Span4Mux_v I__5012 (
            .O(N__21719),
            .I(N__21716));
    Span4Mux_v I__5011 (
            .O(N__21716),
            .I(N__21713));
    Odrv4 I__5010 (
            .O(N__21713),
            .I(\this_sprites_ram.mem_out_bus1_1 ));
    InMux I__5009 (
            .O(N__21710),
            .I(N__21707));
    LocalMux I__5008 (
            .O(N__21707),
            .I(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ));
    InMux I__5007 (
            .O(N__21704),
            .I(N__21701));
    LocalMux I__5006 (
            .O(N__21701),
            .I(N__21698));
    Span4Mux_h I__5005 (
            .O(N__21698),
            .I(N__21695));
    Odrv4 I__5004 (
            .O(N__21695),
            .I(\this_sprites_ram.mem_out_bus4_0 ));
    InMux I__5003 (
            .O(N__21692),
            .I(N__21689));
    LocalMux I__5002 (
            .O(N__21689),
            .I(N__21686));
    Span4Mux_h I__5001 (
            .O(N__21686),
            .I(N__21683));
    Span4Mux_v I__5000 (
            .O(N__21683),
            .I(N__21680));
    Span4Mux_v I__4999 (
            .O(N__21680),
            .I(N__21677));
    Span4Mux_v I__4998 (
            .O(N__21677),
            .I(N__21674));
    Odrv4 I__4997 (
            .O(N__21674),
            .I(\this_sprites_ram.mem_out_bus0_0 ));
    InMux I__4996 (
            .O(N__21671),
            .I(N__21668));
    LocalMux I__4995 (
            .O(N__21668),
            .I(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ));
    CascadeMux I__4994 (
            .O(N__21665),
            .I(N__21662));
    InMux I__4993 (
            .O(N__21662),
            .I(N__21653));
    InMux I__4992 (
            .O(N__21661),
            .I(N__21653));
    InMux I__4991 (
            .O(N__21660),
            .I(N__21653));
    LocalMux I__4990 (
            .O(N__21653),
            .I(M_this_state_qZ0Z_5));
    InMux I__4989 (
            .O(N__21650),
            .I(N__21646));
    InMux I__4988 (
            .O(N__21649),
            .I(N__21643));
    LocalMux I__4987 (
            .O(N__21646),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__4986 (
            .O(N__21643),
            .I(M_this_state_qZ0Z_6));
    CascadeMux I__4985 (
            .O(N__21638),
            .I(N__21630));
    CascadeMux I__4984 (
            .O(N__21637),
            .I(N__21627));
    CascadeMux I__4983 (
            .O(N__21636),
            .I(N__21622));
    CascadeMux I__4982 (
            .O(N__21635),
            .I(N__21619));
    CascadeMux I__4981 (
            .O(N__21634),
            .I(N__21616));
    CascadeMux I__4980 (
            .O(N__21633),
            .I(N__21613));
    InMux I__4979 (
            .O(N__21630),
            .I(N__21609));
    InMux I__4978 (
            .O(N__21627),
            .I(N__21606));
    CascadeMux I__4977 (
            .O(N__21626),
            .I(N__21603));
    CascadeMux I__4976 (
            .O(N__21625),
            .I(N__21598));
    InMux I__4975 (
            .O(N__21622),
            .I(N__21595));
    InMux I__4974 (
            .O(N__21619),
            .I(N__21592));
    InMux I__4973 (
            .O(N__21616),
            .I(N__21587));
    InMux I__4972 (
            .O(N__21613),
            .I(N__21587));
    CascadeMux I__4971 (
            .O(N__21612),
            .I(N__21584));
    LocalMux I__4970 (
            .O(N__21609),
            .I(N__21580));
    LocalMux I__4969 (
            .O(N__21606),
            .I(N__21577));
    InMux I__4968 (
            .O(N__21603),
            .I(N__21572));
    InMux I__4967 (
            .O(N__21602),
            .I(N__21572));
    InMux I__4966 (
            .O(N__21601),
            .I(N__21567));
    InMux I__4965 (
            .O(N__21598),
            .I(N__21567));
    LocalMux I__4964 (
            .O(N__21595),
            .I(N__21563));
    LocalMux I__4963 (
            .O(N__21592),
            .I(N__21560));
    LocalMux I__4962 (
            .O(N__21587),
            .I(N__21557));
    InMux I__4961 (
            .O(N__21584),
            .I(N__21554));
    InMux I__4960 (
            .O(N__21583),
            .I(N__21551));
    Span4Mux_v I__4959 (
            .O(N__21580),
            .I(N__21542));
    Span4Mux_h I__4958 (
            .O(N__21577),
            .I(N__21542));
    LocalMux I__4957 (
            .O(N__21572),
            .I(N__21542));
    LocalMux I__4956 (
            .O(N__21567),
            .I(N__21542));
    CascadeMux I__4955 (
            .O(N__21566),
            .I(N__21538));
    Span4Mux_h I__4954 (
            .O(N__21563),
            .I(N__21535));
    Span4Mux_v I__4953 (
            .O(N__21560),
            .I(N__21528));
    Span4Mux_h I__4952 (
            .O(N__21557),
            .I(N__21528));
    LocalMux I__4951 (
            .O(N__21554),
            .I(N__21528));
    LocalMux I__4950 (
            .O(N__21551),
            .I(N__21525));
    Span4Mux_h I__4949 (
            .O(N__21542),
            .I(N__21522));
    InMux I__4948 (
            .O(N__21541),
            .I(N__21517));
    InMux I__4947 (
            .O(N__21538),
            .I(N__21517));
    Odrv4 I__4946 (
            .O(N__21535),
            .I(N_14_0));
    Odrv4 I__4945 (
            .O(N__21528),
            .I(N_14_0));
    Odrv4 I__4944 (
            .O(N__21525),
            .I(N_14_0));
    Odrv4 I__4943 (
            .O(N__21522),
            .I(N_14_0));
    LocalMux I__4942 (
            .O(N__21517),
            .I(N_14_0));
    CascadeMux I__4941 (
            .O(N__21506),
            .I(N__21503));
    CascadeBuf I__4940 (
            .O(N__21503),
            .I(N__21500));
    CascadeMux I__4939 (
            .O(N__21500),
            .I(N__21497));
    CascadeBuf I__4938 (
            .O(N__21497),
            .I(N__21494));
    CascadeMux I__4937 (
            .O(N__21494),
            .I(N__21491));
    CascadeBuf I__4936 (
            .O(N__21491),
            .I(N__21488));
    CascadeMux I__4935 (
            .O(N__21488),
            .I(N__21485));
    CascadeBuf I__4934 (
            .O(N__21485),
            .I(N__21482));
    CascadeMux I__4933 (
            .O(N__21482),
            .I(N__21479));
    CascadeBuf I__4932 (
            .O(N__21479),
            .I(N__21476));
    CascadeMux I__4931 (
            .O(N__21476),
            .I(N__21473));
    CascadeBuf I__4930 (
            .O(N__21473),
            .I(N__21470));
    CascadeMux I__4929 (
            .O(N__21470),
            .I(N__21467));
    CascadeBuf I__4928 (
            .O(N__21467),
            .I(N__21464));
    CascadeMux I__4927 (
            .O(N__21464),
            .I(N__21461));
    CascadeBuf I__4926 (
            .O(N__21461),
            .I(N__21458));
    CascadeMux I__4925 (
            .O(N__21458),
            .I(N__21455));
    CascadeBuf I__4924 (
            .O(N__21455),
            .I(N__21452));
    CascadeMux I__4923 (
            .O(N__21452),
            .I(N__21449));
    CascadeBuf I__4922 (
            .O(N__21449),
            .I(N__21446));
    CascadeMux I__4921 (
            .O(N__21446),
            .I(N__21443));
    CascadeBuf I__4920 (
            .O(N__21443),
            .I(N__21440));
    CascadeMux I__4919 (
            .O(N__21440),
            .I(N__21437));
    CascadeBuf I__4918 (
            .O(N__21437),
            .I(N__21434));
    CascadeMux I__4917 (
            .O(N__21434),
            .I(N__21431));
    CascadeBuf I__4916 (
            .O(N__21431),
            .I(N__21428));
    CascadeMux I__4915 (
            .O(N__21428),
            .I(N__21425));
    CascadeBuf I__4914 (
            .O(N__21425),
            .I(N__21422));
    CascadeMux I__4913 (
            .O(N__21422),
            .I(N__21419));
    CascadeBuf I__4912 (
            .O(N__21419),
            .I(N__21416));
    CascadeMux I__4911 (
            .O(N__21416),
            .I(N__21413));
    InMux I__4910 (
            .O(N__21413),
            .I(N__21410));
    LocalMux I__4909 (
            .O(N__21410),
            .I(N__21407));
    Span4Mux_s1_v I__4908 (
            .O(N__21407),
            .I(N__21403));
    InMux I__4907 (
            .O(N__21406),
            .I(N__21400));
    Sp12to4 I__4906 (
            .O(N__21403),
            .I(N__21396));
    LocalMux I__4905 (
            .O(N__21400),
            .I(N__21393));
    InMux I__4904 (
            .O(N__21399),
            .I(N__21390));
    Span12Mux_h I__4903 (
            .O(N__21396),
            .I(N__21387));
    Odrv12 I__4902 (
            .O(N__21393),
            .I(M_this_internal_address_qZ0Z_5));
    LocalMux I__4901 (
            .O(N__21390),
            .I(M_this_internal_address_qZ0Z_5));
    Odrv12 I__4900 (
            .O(N__21387),
            .I(M_this_internal_address_qZ0Z_5));
    InMux I__4899 (
            .O(N__21380),
            .I(N__21377));
    LocalMux I__4898 (
            .O(N__21377),
            .I(M_this_internal_address_q_3_ns_1_5));
    CascadeMux I__4897 (
            .O(N__21374),
            .I(N__21371));
    CascadeBuf I__4896 (
            .O(N__21371),
            .I(N__21368));
    CascadeMux I__4895 (
            .O(N__21368),
            .I(N__21365));
    CascadeBuf I__4894 (
            .O(N__21365),
            .I(N__21362));
    CascadeMux I__4893 (
            .O(N__21362),
            .I(N__21359));
    CascadeBuf I__4892 (
            .O(N__21359),
            .I(N__21356));
    CascadeMux I__4891 (
            .O(N__21356),
            .I(N__21353));
    CascadeBuf I__4890 (
            .O(N__21353),
            .I(N__21350));
    CascadeMux I__4889 (
            .O(N__21350),
            .I(N__21347));
    CascadeBuf I__4888 (
            .O(N__21347),
            .I(N__21344));
    CascadeMux I__4887 (
            .O(N__21344),
            .I(N__21341));
    CascadeBuf I__4886 (
            .O(N__21341),
            .I(N__21338));
    CascadeMux I__4885 (
            .O(N__21338),
            .I(N__21335));
    CascadeBuf I__4884 (
            .O(N__21335),
            .I(N__21332));
    CascadeMux I__4883 (
            .O(N__21332),
            .I(N__21329));
    CascadeBuf I__4882 (
            .O(N__21329),
            .I(N__21326));
    CascadeMux I__4881 (
            .O(N__21326),
            .I(N__21323));
    CascadeBuf I__4880 (
            .O(N__21323),
            .I(N__21320));
    CascadeMux I__4879 (
            .O(N__21320),
            .I(N__21317));
    CascadeBuf I__4878 (
            .O(N__21317),
            .I(N__21314));
    CascadeMux I__4877 (
            .O(N__21314),
            .I(N__21311));
    CascadeBuf I__4876 (
            .O(N__21311),
            .I(N__21308));
    CascadeMux I__4875 (
            .O(N__21308),
            .I(N__21305));
    CascadeBuf I__4874 (
            .O(N__21305),
            .I(N__21302));
    CascadeMux I__4873 (
            .O(N__21302),
            .I(N__21299));
    CascadeBuf I__4872 (
            .O(N__21299),
            .I(N__21296));
    CascadeMux I__4871 (
            .O(N__21296),
            .I(N__21293));
    CascadeBuf I__4870 (
            .O(N__21293),
            .I(N__21290));
    CascadeMux I__4869 (
            .O(N__21290),
            .I(N__21287));
    CascadeBuf I__4868 (
            .O(N__21287),
            .I(N__21284));
    CascadeMux I__4867 (
            .O(N__21284),
            .I(N__21281));
    InMux I__4866 (
            .O(N__21281),
            .I(N__21276));
    CascadeMux I__4865 (
            .O(N__21280),
            .I(N__21273));
    InMux I__4864 (
            .O(N__21279),
            .I(N__21270));
    LocalMux I__4863 (
            .O(N__21276),
            .I(N__21267));
    InMux I__4862 (
            .O(N__21273),
            .I(N__21264));
    LocalMux I__4861 (
            .O(N__21270),
            .I(N__21261));
    Span12Mux_h I__4860 (
            .O(N__21267),
            .I(N__21258));
    LocalMux I__4859 (
            .O(N__21264),
            .I(M_this_internal_address_qZ0Z_6));
    Odrv4 I__4858 (
            .O(N__21261),
            .I(M_this_internal_address_qZ0Z_6));
    Odrv12 I__4857 (
            .O(N__21258),
            .I(M_this_internal_address_qZ0Z_6));
    CascadeMux I__4856 (
            .O(N__21251),
            .I(N__21248));
    InMux I__4855 (
            .O(N__21248),
            .I(N__21245));
    LocalMux I__4854 (
            .O(N__21245),
            .I(M_this_internal_address_q_3_ns_1_6));
    InMux I__4853 (
            .O(N__21242),
            .I(N__21239));
    LocalMux I__4852 (
            .O(N__21239),
            .I(N__21236));
    Odrv12 I__4851 (
            .O(N__21236),
            .I(M_this_internal_address_q_3_ns_1_13));
    InMux I__4850 (
            .O(N__21233),
            .I(N__21226));
    InMux I__4849 (
            .O(N__21232),
            .I(N__21226));
    CascadeMux I__4848 (
            .O(N__21231),
            .I(N__21220));
    LocalMux I__4847 (
            .O(N__21226),
            .I(N__21216));
    InMux I__4846 (
            .O(N__21225),
            .I(N__21207));
    InMux I__4845 (
            .O(N__21224),
            .I(N__21207));
    InMux I__4844 (
            .O(N__21223),
            .I(N__21204));
    InMux I__4843 (
            .O(N__21220),
            .I(N__21199));
    InMux I__4842 (
            .O(N__21219),
            .I(N__21199));
    Span4Mux_v I__4841 (
            .O(N__21216),
            .I(N__21193));
    InMux I__4840 (
            .O(N__21215),
            .I(N__21190));
    InMux I__4839 (
            .O(N__21214),
            .I(N__21183));
    InMux I__4838 (
            .O(N__21213),
            .I(N__21183));
    InMux I__4837 (
            .O(N__21212),
            .I(N__21183));
    LocalMux I__4836 (
            .O(N__21207),
            .I(N__21178));
    LocalMux I__4835 (
            .O(N__21204),
            .I(N__21178));
    LocalMux I__4834 (
            .O(N__21199),
            .I(N__21175));
    InMux I__4833 (
            .O(N__21198),
            .I(N__21172));
    InMux I__4832 (
            .O(N__21197),
            .I(N__21166));
    InMux I__4831 (
            .O(N__21196),
            .I(N__21163));
    Span4Mux_h I__4830 (
            .O(N__21193),
            .I(N__21160));
    LocalMux I__4829 (
            .O(N__21190),
            .I(N__21155));
    LocalMux I__4828 (
            .O(N__21183),
            .I(N__21155));
    Span4Mux_h I__4827 (
            .O(N__21178),
            .I(N__21152));
    Span4Mux_v I__4826 (
            .O(N__21175),
            .I(N__21147));
    LocalMux I__4825 (
            .O(N__21172),
            .I(N__21147));
    InMux I__4824 (
            .O(N__21171),
            .I(N__21142));
    InMux I__4823 (
            .O(N__21170),
            .I(N__21142));
    InMux I__4822 (
            .O(N__21169),
            .I(N__21139));
    LocalMux I__4821 (
            .O(N__21166),
            .I(N_355));
    LocalMux I__4820 (
            .O(N__21163),
            .I(N_355));
    Odrv4 I__4819 (
            .O(N__21160),
            .I(N_355));
    Odrv12 I__4818 (
            .O(N__21155),
            .I(N_355));
    Odrv4 I__4817 (
            .O(N__21152),
            .I(N_355));
    Odrv4 I__4816 (
            .O(N__21147),
            .I(N_355));
    LocalMux I__4815 (
            .O(N__21142),
            .I(N_355));
    LocalMux I__4814 (
            .O(N__21139),
            .I(N_355));
    InMux I__4813 (
            .O(N__21122),
            .I(N__21119));
    LocalMux I__4812 (
            .O(N__21119),
            .I(M_this_internal_address_q_3_ns_1_12));
    InMux I__4811 (
            .O(N__21116),
            .I(N__21110));
    InMux I__4810 (
            .O(N__21115),
            .I(N__21107));
    InMux I__4809 (
            .O(N__21114),
            .I(N__21104));
    InMux I__4808 (
            .O(N__21113),
            .I(N__21101));
    LocalMux I__4807 (
            .O(N__21110),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__4806 (
            .O(N__21107),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__4805 (
            .O(N__21104),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__4804 (
            .O(N__21101),
            .I(M_this_state_qZ0Z_7));
    CascadeMux I__4803 (
            .O(N__21092),
            .I(N__21088));
    CascadeMux I__4802 (
            .O(N__21091),
            .I(N__21085));
    InMux I__4801 (
            .O(N__21088),
            .I(N__21082));
    InMux I__4800 (
            .O(N__21085),
            .I(N__21079));
    LocalMux I__4799 (
            .O(N__21082),
            .I(N__21073));
    LocalMux I__4798 (
            .O(N__21079),
            .I(N__21073));
    InMux I__4797 (
            .O(N__21078),
            .I(N__21070));
    Span4Mux_v I__4796 (
            .O(N__21073),
            .I(N__21067));
    LocalMux I__4795 (
            .O(N__21070),
            .I(N__21064));
    Sp12to4 I__4794 (
            .O(N__21067),
            .I(N__21061));
    Span4Mux_v I__4793 (
            .O(N__21064),
            .I(N__21058));
    Span12Mux_h I__4792 (
            .O(N__21061),
            .I(N__21055));
    Sp12to4 I__4791 (
            .O(N__21058),
            .I(N__21052));
    Odrv12 I__4790 (
            .O(N__21055),
            .I(port_data_c_5));
    Odrv12 I__4789 (
            .O(N__21052),
            .I(port_data_c_5));
    CascadeMux I__4788 (
            .O(N__21047),
            .I(N__21044));
    InMux I__4787 (
            .O(N__21044),
            .I(N__21039));
    CascadeMux I__4786 (
            .O(N__21043),
            .I(N__21036));
    CascadeMux I__4785 (
            .O(N__21042),
            .I(N__21032));
    LocalMux I__4784 (
            .O(N__21039),
            .I(N__21029));
    InMux I__4783 (
            .O(N__21036),
            .I(N__21026));
    CascadeMux I__4782 (
            .O(N__21035),
            .I(N__21023));
    InMux I__4781 (
            .O(N__21032),
            .I(N__21020));
    Span4Mux_v I__4780 (
            .O(N__21029),
            .I(N__21017));
    LocalMux I__4779 (
            .O(N__21026),
            .I(N__21014));
    InMux I__4778 (
            .O(N__21023),
            .I(N__21011));
    LocalMux I__4777 (
            .O(N__21020),
            .I(N__21008));
    Span4Mux_h I__4776 (
            .O(N__21017),
            .I(N__21001));
    Span4Mux_v I__4775 (
            .O(N__21014),
            .I(N__21001));
    LocalMux I__4774 (
            .O(N__21011),
            .I(N__21001));
    Span4Mux_v I__4773 (
            .O(N__21008),
            .I(N__20998));
    Span4Mux_h I__4772 (
            .O(N__21001),
            .I(N__20995));
    Sp12to4 I__4771 (
            .O(N__20998),
            .I(N__20992));
    Span4Mux_v I__4770 (
            .O(N__20995),
            .I(N__20989));
    Span12Mux_h I__4769 (
            .O(N__20992),
            .I(N__20986));
    Span4Mux_v I__4768 (
            .O(N__20989),
            .I(N__20983));
    Span12Mux_v I__4767 (
            .O(N__20986),
            .I(N__20980));
    Span4Mux_v I__4766 (
            .O(N__20983),
            .I(N__20977));
    Odrv12 I__4765 (
            .O(N__20980),
            .I(port_data_c_1));
    Odrv4 I__4764 (
            .O(N__20977),
            .I(port_data_c_1));
    InMux I__4763 (
            .O(N__20972),
            .I(N__20969));
    LocalMux I__4762 (
            .O(N__20969),
            .I(N__20963));
    InMux I__4761 (
            .O(N__20968),
            .I(N__20960));
    InMux I__4760 (
            .O(N__20967),
            .I(N__20957));
    InMux I__4759 (
            .O(N__20966),
            .I(N__20953));
    Span4Mux_h I__4758 (
            .O(N__20963),
            .I(N__20949));
    LocalMux I__4757 (
            .O(N__20960),
            .I(N__20946));
    LocalMux I__4756 (
            .O(N__20957),
            .I(N__20943));
    InMux I__4755 (
            .O(N__20956),
            .I(N__20940));
    LocalMux I__4754 (
            .O(N__20953),
            .I(N__20935));
    InMux I__4753 (
            .O(N__20952),
            .I(N__20932));
    Span4Mux_v I__4752 (
            .O(N__20949),
            .I(N__20927));
    Span4Mux_h I__4751 (
            .O(N__20946),
            .I(N__20927));
    Span4Mux_v I__4750 (
            .O(N__20943),
            .I(N__20922));
    LocalMux I__4749 (
            .O(N__20940),
            .I(N__20922));
    InMux I__4748 (
            .O(N__20939),
            .I(N__20919));
    InMux I__4747 (
            .O(N__20938),
            .I(N__20916));
    Span12Mux_s11_h I__4746 (
            .O(N__20935),
            .I(N__20913));
    LocalMux I__4745 (
            .O(N__20932),
            .I(N__20910));
    Span4Mux_v I__4744 (
            .O(N__20927),
            .I(N__20907));
    Span4Mux_v I__4743 (
            .O(N__20922),
            .I(N__20902));
    LocalMux I__4742 (
            .O(N__20919),
            .I(N__20902));
    LocalMux I__4741 (
            .O(N__20916),
            .I(N__20899));
    Span12Mux_v I__4740 (
            .O(N__20913),
            .I(N__20894));
    Span12Mux_s11_h I__4739 (
            .O(N__20910),
            .I(N__20894));
    Span4Mux_v I__4738 (
            .O(N__20907),
            .I(N__20887));
    Span4Mux_h I__4737 (
            .O(N__20902),
            .I(N__20887));
    Span4Mux_h I__4736 (
            .O(N__20899),
            .I(N__20887));
    Odrv12 I__4735 (
            .O(N__20894),
            .I(M_this_sprites_ram_write_data_1));
    Odrv4 I__4734 (
            .O(N__20887),
            .I(M_this_sprites_ram_write_data_1));
    InMux I__4733 (
            .O(N__20882),
            .I(N__20878));
    InMux I__4732 (
            .O(N__20881),
            .I(N__20875));
    LocalMux I__4731 (
            .O(N__20878),
            .I(N__20870));
    LocalMux I__4730 (
            .O(N__20875),
            .I(N__20867));
    CascadeMux I__4729 (
            .O(N__20874),
            .I(N__20864));
    CascadeMux I__4728 (
            .O(N__20873),
            .I(N__20861));
    Span12Mux_h I__4727 (
            .O(N__20870),
            .I(N__20858));
    Span4Mux_v I__4726 (
            .O(N__20867),
            .I(N__20855));
    InMux I__4725 (
            .O(N__20864),
            .I(N__20850));
    InMux I__4724 (
            .O(N__20861),
            .I(N__20850));
    Span12Mux_v I__4723 (
            .O(N__20858),
            .I(N__20847));
    Sp12to4 I__4722 (
            .O(N__20855),
            .I(N__20842));
    LocalMux I__4721 (
            .O(N__20850),
            .I(N__20842));
    Span12Mux_h I__4720 (
            .O(N__20847),
            .I(N__20839));
    Span12Mux_h I__4719 (
            .O(N__20842),
            .I(N__20836));
    Odrv12 I__4718 (
            .O(N__20839),
            .I(port_data_c_0));
    Odrv12 I__4717 (
            .O(N__20836),
            .I(port_data_c_0));
    CascadeMux I__4716 (
            .O(N__20831),
            .I(N__20828));
    InMux I__4715 (
            .O(N__20828),
            .I(N__20824));
    CascadeMux I__4714 (
            .O(N__20827),
            .I(N__20820));
    LocalMux I__4713 (
            .O(N__20824),
            .I(N__20817));
    InMux I__4712 (
            .O(N__20823),
            .I(N__20812));
    InMux I__4711 (
            .O(N__20820),
            .I(N__20812));
    Span4Mux_v I__4710 (
            .O(N__20817),
            .I(N__20809));
    LocalMux I__4709 (
            .O(N__20812),
            .I(N__20806));
    Span4Mux_v I__4708 (
            .O(N__20809),
            .I(N__20803));
    Span12Mux_v I__4707 (
            .O(N__20806),
            .I(N__20800));
    Sp12to4 I__4706 (
            .O(N__20803),
            .I(N__20797));
    Span12Mux_h I__4705 (
            .O(N__20800),
            .I(N__20794));
    Odrv12 I__4704 (
            .O(N__20797),
            .I(port_data_c_4));
    Odrv12 I__4703 (
            .O(N__20794),
            .I(port_data_c_4));
    InMux I__4702 (
            .O(N__20789),
            .I(N__20786));
    LocalMux I__4701 (
            .O(N__20786),
            .I(N__20782));
    InMux I__4700 (
            .O(N__20785),
            .I(N__20779));
    Span4Mux_h I__4699 (
            .O(N__20782),
            .I(N__20774));
    LocalMux I__4698 (
            .O(N__20779),
            .I(N__20771));
    InMux I__4697 (
            .O(N__20778),
            .I(N__20768));
    InMux I__4696 (
            .O(N__20777),
            .I(N__20764));
    Span4Mux_v I__4695 (
            .O(N__20774),
            .I(N__20758));
    Span4Mux_h I__4694 (
            .O(N__20771),
            .I(N__20758));
    LocalMux I__4693 (
            .O(N__20768),
            .I(N__20755));
    InMux I__4692 (
            .O(N__20767),
            .I(N__20752));
    LocalMux I__4691 (
            .O(N__20764),
            .I(N__20749));
    InMux I__4690 (
            .O(N__20763),
            .I(N__20746));
    Span4Mux_v I__4689 (
            .O(N__20758),
            .I(N__20739));
    Span4Mux_h I__4688 (
            .O(N__20755),
            .I(N__20739));
    LocalMux I__4687 (
            .O(N__20752),
            .I(N__20736));
    Span4Mux_v I__4686 (
            .O(N__20749),
            .I(N__20731));
    LocalMux I__4685 (
            .O(N__20746),
            .I(N__20731));
    InMux I__4684 (
            .O(N__20745),
            .I(N__20728));
    InMux I__4683 (
            .O(N__20744),
            .I(N__20725));
    Span4Mux_v I__4682 (
            .O(N__20739),
            .I(N__20720));
    Span4Mux_h I__4681 (
            .O(N__20736),
            .I(N__20720));
    Span4Mux_h I__4680 (
            .O(N__20731),
            .I(N__20717));
    LocalMux I__4679 (
            .O(N__20728),
            .I(N__20714));
    LocalMux I__4678 (
            .O(N__20725),
            .I(N__20711));
    Span4Mux_v I__4677 (
            .O(N__20720),
            .I(N__20702));
    Span4Mux_v I__4676 (
            .O(N__20717),
            .I(N__20702));
    Span4Mux_h I__4675 (
            .O(N__20714),
            .I(N__20702));
    Span4Mux_h I__4674 (
            .O(N__20711),
            .I(N__20702));
    Odrv4 I__4673 (
            .O(N__20702),
            .I(M_this_sprites_ram_write_data_0));
    InMux I__4672 (
            .O(N__20699),
            .I(N__20696));
    LocalMux I__4671 (
            .O(N__20696),
            .I(N__20693));
    Span4Mux_v I__4670 (
            .O(N__20693),
            .I(N__20690));
    Sp12to4 I__4669 (
            .O(N__20690),
            .I(N__20687));
    Span12Mux_h I__4668 (
            .O(N__20687),
            .I(N__20684));
    Span12Mux_v I__4667 (
            .O(N__20684),
            .I(N__20681));
    Odrv12 I__4666 (
            .O(N__20681),
            .I(port_address_in_7));
    InMux I__4665 (
            .O(N__20678),
            .I(N__20675));
    LocalMux I__4664 (
            .O(N__20675),
            .I(N__20672));
    Sp12to4 I__4663 (
            .O(N__20672),
            .I(N__20669));
    Span12Mux_v I__4662 (
            .O(N__20669),
            .I(N__20666));
    Span12Mux_h I__4661 (
            .O(N__20666),
            .I(N__20663));
    Odrv12 I__4660 (
            .O(N__20663),
            .I(port_address_in_6));
    CascadeMux I__4659 (
            .O(N__20660),
            .I(N__20657));
    InMux I__4658 (
            .O(N__20657),
            .I(N__20654));
    LocalMux I__4657 (
            .O(N__20654),
            .I(N__20651));
    Span4Mux_v I__4656 (
            .O(N__20651),
            .I(N__20648));
    Span4Mux_v I__4655 (
            .O(N__20648),
            .I(N__20645));
    Sp12to4 I__4654 (
            .O(N__20645),
            .I(N__20642));
    Span12Mux_h I__4653 (
            .O(N__20642),
            .I(N__20638));
    InMux I__4652 (
            .O(N__20641),
            .I(N__20635));
    Odrv12 I__4651 (
            .O(N__20638),
            .I(port_rw_in));
    LocalMux I__4650 (
            .O(N__20635),
            .I(port_rw_in));
    CascadeMux I__4649 (
            .O(N__20630),
            .I(N__20627));
    InMux I__4648 (
            .O(N__20627),
            .I(N__20622));
    InMux I__4647 (
            .O(N__20626),
            .I(N__20619));
    InMux I__4646 (
            .O(N__20625),
            .I(N__20616));
    LocalMux I__4645 (
            .O(N__20622),
            .I(N__20611));
    LocalMux I__4644 (
            .O(N__20619),
            .I(N__20611));
    LocalMux I__4643 (
            .O(N__20616),
            .I(N__20608));
    Span4Mux_h I__4642 (
            .O(N__20611),
            .I(N__20603));
    Span4Mux_h I__4641 (
            .O(N__20608),
            .I(N__20603));
    Odrv4 I__4640 (
            .O(N__20603),
            .I(\this_vga_signals.N_185_0 ));
    InMux I__4639 (
            .O(N__20600),
            .I(N__20597));
    LocalMux I__4638 (
            .O(N__20597),
            .I(N__20594));
    Odrv4 I__4637 (
            .O(N__20594),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4 ));
    CascadeMux I__4636 (
            .O(N__20591),
            .I(N__20586));
    InMux I__4635 (
            .O(N__20590),
            .I(N__20583));
    CascadeMux I__4634 (
            .O(N__20589),
            .I(N__20580));
    InMux I__4633 (
            .O(N__20586),
            .I(N__20577));
    LocalMux I__4632 (
            .O(N__20583),
            .I(N__20574));
    InMux I__4631 (
            .O(N__20580),
            .I(N__20571));
    LocalMux I__4630 (
            .O(N__20577),
            .I(N__20568));
    Odrv4 I__4629 (
            .O(N__20574),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__4628 (
            .O(N__20571),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__4627 (
            .O(N__20568),
            .I(M_this_state_qZ0Z_4));
    CascadeMux I__4626 (
            .O(N__20561),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4_cascade_ ));
    CascadeMux I__4625 (
            .O(N__20558),
            .I(\this_vga_signals.N_490_cascade_ ));
    CascadeMux I__4624 (
            .O(N__20555),
            .I(\this_vga_signals.N_386_cascade_ ));
    CascadeMux I__4623 (
            .O(N__20552),
            .I(\this_vga_signals.N_387_cascade_ ));
    CascadeMux I__4622 (
            .O(N__20549),
            .I(N__20546));
    InMux I__4621 (
            .O(N__20546),
            .I(N__20540));
    InMux I__4620 (
            .O(N__20545),
            .I(N__20537));
    InMux I__4619 (
            .O(N__20544),
            .I(N__20532));
    InMux I__4618 (
            .O(N__20543),
            .I(N__20532));
    LocalMux I__4617 (
            .O(N__20540),
            .I(N__20529));
    LocalMux I__4616 (
            .O(N__20537),
            .I(N__20524));
    LocalMux I__4615 (
            .O(N__20532),
            .I(N__20524));
    Span4Mux_v I__4614 (
            .O(N__20529),
            .I(N__20521));
    Span4Mux_v I__4613 (
            .O(N__20524),
            .I(N__20518));
    Sp12to4 I__4612 (
            .O(N__20521),
            .I(N__20513));
    Sp12to4 I__4611 (
            .O(N__20518),
            .I(N__20513));
    Span12Mux_h I__4610 (
            .O(N__20513),
            .I(N__20510));
    Odrv12 I__4609 (
            .O(N__20510),
            .I(port_address_in_1));
    InMux I__4608 (
            .O(N__20507),
            .I(N__20502));
    InMux I__4607 (
            .O(N__20506),
            .I(N__20499));
    InMux I__4606 (
            .O(N__20505),
            .I(N__20496));
    LocalMux I__4605 (
            .O(N__20502),
            .I(N__20491));
    LocalMux I__4604 (
            .O(N__20499),
            .I(N__20491));
    LocalMux I__4603 (
            .O(N__20496),
            .I(N__20488));
    Span4Mux_v I__4602 (
            .O(N__20491),
            .I(N__20482));
    Span4Mux_v I__4601 (
            .O(N__20488),
            .I(N__20482));
    InMux I__4600 (
            .O(N__20487),
            .I(N__20479));
    Sp12to4 I__4599 (
            .O(N__20482),
            .I(N__20476));
    LocalMux I__4598 (
            .O(N__20479),
            .I(N__20473));
    Span12Mux_h I__4597 (
            .O(N__20476),
            .I(N__20470));
    Span12Mux_v I__4596 (
            .O(N__20473),
            .I(N__20467));
    Odrv12 I__4595 (
            .O(N__20470),
            .I(port_address_in_0));
    Odrv12 I__4594 (
            .O(N__20467),
            .I(port_address_in_0));
    CascadeMux I__4593 (
            .O(N__20462),
            .I(\this_vga_signals.N_391_cascade_ ));
    InMux I__4592 (
            .O(N__20459),
            .I(N__20453));
    InMux I__4591 (
            .O(N__20458),
            .I(N__20453));
    LocalMux I__4590 (
            .O(N__20453),
            .I(\this_vga_signals.N_490 ));
    InMux I__4589 (
            .O(N__20450),
            .I(N__20442));
    InMux I__4588 (
            .O(N__20449),
            .I(N__20439));
    InMux I__4587 (
            .O(N__20448),
            .I(N__20436));
    InMux I__4586 (
            .O(N__20447),
            .I(N__20433));
    InMux I__4585 (
            .O(N__20446),
            .I(N__20428));
    InMux I__4584 (
            .O(N__20445),
            .I(N__20428));
    LocalMux I__4583 (
            .O(N__20442),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__4582 (
            .O(N__20439),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__4581 (
            .O(N__20436),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__4580 (
            .O(N__20433),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__4579 (
            .O(N__20428),
            .I(M_this_state_qZ0Z_2));
    InMux I__4578 (
            .O(N__20417),
            .I(N__20414));
    LocalMux I__4577 (
            .O(N__20414),
            .I(N__20411));
    Odrv4 I__4576 (
            .O(N__20411),
            .I(M_this_internal_address_q_RNO_1Z0Z_5));
    InMux I__4575 (
            .O(N__20408),
            .I(N__20405));
    LocalMux I__4574 (
            .O(N__20405),
            .I(N__20402));
    Odrv4 I__4573 (
            .O(N__20402),
            .I(M_this_internal_address_q_RNO_1Z0Z_6));
    InMux I__4572 (
            .O(N__20399),
            .I(N__20396));
    LocalMux I__4571 (
            .O(N__20396),
            .I(N__20393));
    Odrv4 I__4570 (
            .O(N__20393),
            .I(M_this_internal_address_q_RNO_1Z0Z_12));
    InMux I__4569 (
            .O(N__20390),
            .I(N__20387));
    LocalMux I__4568 (
            .O(N__20387),
            .I(M_this_internal_address_q_3_ns_1_11));
    InMux I__4567 (
            .O(N__20384),
            .I(N__20381));
    LocalMux I__4566 (
            .O(N__20381),
            .I(M_this_internal_address_q_3_ns_1_4));
    InMux I__4565 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__4564 (
            .O(N__20375),
            .I(N__20372));
    Span4Mux_h I__4563 (
            .O(N__20372),
            .I(N__20369));
    Odrv4 I__4562 (
            .O(N__20369),
            .I(M_this_internal_address_q_RNO_1Z0Z_4));
    CascadeMux I__4561 (
            .O(N__20366),
            .I(N__20363));
    CascadeBuf I__4560 (
            .O(N__20363),
            .I(N__20360));
    CascadeMux I__4559 (
            .O(N__20360),
            .I(N__20357));
    CascadeBuf I__4558 (
            .O(N__20357),
            .I(N__20354));
    CascadeMux I__4557 (
            .O(N__20354),
            .I(N__20351));
    CascadeBuf I__4556 (
            .O(N__20351),
            .I(N__20348));
    CascadeMux I__4555 (
            .O(N__20348),
            .I(N__20345));
    CascadeBuf I__4554 (
            .O(N__20345),
            .I(N__20342));
    CascadeMux I__4553 (
            .O(N__20342),
            .I(N__20339));
    CascadeBuf I__4552 (
            .O(N__20339),
            .I(N__20336));
    CascadeMux I__4551 (
            .O(N__20336),
            .I(N__20333));
    CascadeBuf I__4550 (
            .O(N__20333),
            .I(N__20330));
    CascadeMux I__4549 (
            .O(N__20330),
            .I(N__20327));
    CascadeBuf I__4548 (
            .O(N__20327),
            .I(N__20324));
    CascadeMux I__4547 (
            .O(N__20324),
            .I(N__20321));
    CascadeBuf I__4546 (
            .O(N__20321),
            .I(N__20318));
    CascadeMux I__4545 (
            .O(N__20318),
            .I(N__20315));
    CascadeBuf I__4544 (
            .O(N__20315),
            .I(N__20312));
    CascadeMux I__4543 (
            .O(N__20312),
            .I(N__20309));
    CascadeBuf I__4542 (
            .O(N__20309),
            .I(N__20306));
    CascadeMux I__4541 (
            .O(N__20306),
            .I(N__20303));
    CascadeBuf I__4540 (
            .O(N__20303),
            .I(N__20300));
    CascadeMux I__4539 (
            .O(N__20300),
            .I(N__20297));
    CascadeBuf I__4538 (
            .O(N__20297),
            .I(N__20294));
    CascadeMux I__4537 (
            .O(N__20294),
            .I(N__20291));
    CascadeBuf I__4536 (
            .O(N__20291),
            .I(N__20288));
    CascadeMux I__4535 (
            .O(N__20288),
            .I(N__20285));
    CascadeBuf I__4534 (
            .O(N__20285),
            .I(N__20282));
    CascadeMux I__4533 (
            .O(N__20282),
            .I(N__20279));
    CascadeBuf I__4532 (
            .O(N__20279),
            .I(N__20276));
    CascadeMux I__4531 (
            .O(N__20276),
            .I(N__20273));
    InMux I__4530 (
            .O(N__20273),
            .I(N__20270));
    LocalMux I__4529 (
            .O(N__20270),
            .I(N__20266));
    InMux I__4528 (
            .O(N__20269),
            .I(N__20263));
    Span4Mux_v I__4527 (
            .O(N__20266),
            .I(N__20260));
    LocalMux I__4526 (
            .O(N__20263),
            .I(N__20256));
    Span4Mux_h I__4525 (
            .O(N__20260),
            .I(N__20253));
    InMux I__4524 (
            .O(N__20259),
            .I(N__20250));
    Span4Mux_v I__4523 (
            .O(N__20256),
            .I(N__20245));
    Span4Mux_v I__4522 (
            .O(N__20253),
            .I(N__20245));
    LocalMux I__4521 (
            .O(N__20250),
            .I(M_this_internal_address_qZ0Z_4));
    Odrv4 I__4520 (
            .O(N__20245),
            .I(M_this_internal_address_qZ0Z_4));
    InMux I__4519 (
            .O(N__20240),
            .I(N__20237));
    LocalMux I__4518 (
            .O(N__20237),
            .I(N__20234));
    Span4Mux_h I__4517 (
            .O(N__20234),
            .I(N__20231));
    Span4Mux_h I__4516 (
            .O(N__20231),
            .I(N__20228));
    Span4Mux_h I__4515 (
            .O(N__20228),
            .I(N__20225));
    Odrv4 I__4514 (
            .O(N__20225),
            .I(M_this_vram_write_data_1));
    IoInMux I__4513 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__4512 (
            .O(N__20219),
            .I(N__20215));
    InMux I__4511 (
            .O(N__20218),
            .I(N__20211));
    Span4Mux_s3_h I__4510 (
            .O(N__20215),
            .I(N__20208));
    InMux I__4509 (
            .O(N__20214),
            .I(N__20205));
    LocalMux I__4508 (
            .O(N__20211),
            .I(N__20202));
    Span4Mux_v I__4507 (
            .O(N__20208),
            .I(N__20199));
    LocalMux I__4506 (
            .O(N__20205),
            .I(N__20196));
    Span4Mux_v I__4505 (
            .O(N__20202),
            .I(N__20193));
    Sp12to4 I__4504 (
            .O(N__20199),
            .I(N__20189));
    Span4Mux_v I__4503 (
            .O(N__20196),
            .I(N__20186));
    Span4Mux_v I__4502 (
            .O(N__20193),
            .I(N__20183));
    InMux I__4501 (
            .O(N__20192),
            .I(N__20180));
    Span12Mux_h I__4500 (
            .O(N__20189),
            .I(N__20177));
    Sp12to4 I__4499 (
            .O(N__20186),
            .I(N__20174));
    Span4Mux_h I__4498 (
            .O(N__20183),
            .I(N__20171));
    LocalMux I__4497 (
            .O(N__20180),
            .I(N__20168));
    Span12Mux_v I__4496 (
            .O(N__20177),
            .I(N__20162));
    Span12Mux_h I__4495 (
            .O(N__20174),
            .I(N__20162));
    Span4Mux_h I__4494 (
            .O(N__20171),
            .I(N__20157));
    Span4Mux_v I__4493 (
            .O(N__20168),
            .I(N__20157));
    InMux I__4492 (
            .O(N__20167),
            .I(N__20154));
    Odrv12 I__4491 (
            .O(N__20162),
            .I(N_235_0));
    Odrv4 I__4490 (
            .O(N__20157),
            .I(N_235_0));
    LocalMux I__4489 (
            .O(N__20154),
            .I(N_235_0));
    InMux I__4488 (
            .O(N__20147),
            .I(N__20144));
    LocalMux I__4487 (
            .O(N__20144),
            .I(\this_vga_signals.N_319 ));
    CascadeMux I__4486 (
            .O(N__20141),
            .I(N__20137));
    InMux I__4485 (
            .O(N__20140),
            .I(N__20134));
    InMux I__4484 (
            .O(N__20137),
            .I(N__20131));
    LocalMux I__4483 (
            .O(N__20134),
            .I(un19_i_i_i_a2));
    LocalMux I__4482 (
            .O(N__20131),
            .I(un19_i_i_i_a2));
    InMux I__4481 (
            .O(N__20126),
            .I(N__20123));
    LocalMux I__4480 (
            .O(N__20123),
            .I(M_this_internal_address_q_RNO_1Z0Z_11));
    InMux I__4479 (
            .O(N__20120),
            .I(N__20117));
    LocalMux I__4478 (
            .O(N__20117),
            .I(M_this_internal_address_q_3_ns_1_0));
    InMux I__4477 (
            .O(N__20114),
            .I(N__20111));
    LocalMux I__4476 (
            .O(N__20111),
            .I(N__20108));
    Odrv4 I__4475 (
            .O(N__20108),
            .I(M_this_internal_address_q_RNO_1Z0Z_0));
    CascadeMux I__4474 (
            .O(N__20105),
            .I(N__20102));
    CascadeBuf I__4473 (
            .O(N__20102),
            .I(N__20099));
    CascadeMux I__4472 (
            .O(N__20099),
            .I(N__20096));
    CascadeBuf I__4471 (
            .O(N__20096),
            .I(N__20093));
    CascadeMux I__4470 (
            .O(N__20093),
            .I(N__20090));
    CascadeBuf I__4469 (
            .O(N__20090),
            .I(N__20087));
    CascadeMux I__4468 (
            .O(N__20087),
            .I(N__20084));
    CascadeBuf I__4467 (
            .O(N__20084),
            .I(N__20081));
    CascadeMux I__4466 (
            .O(N__20081),
            .I(N__20078));
    CascadeBuf I__4465 (
            .O(N__20078),
            .I(N__20075));
    CascadeMux I__4464 (
            .O(N__20075),
            .I(N__20072));
    CascadeBuf I__4463 (
            .O(N__20072),
            .I(N__20069));
    CascadeMux I__4462 (
            .O(N__20069),
            .I(N__20066));
    CascadeBuf I__4461 (
            .O(N__20066),
            .I(N__20063));
    CascadeMux I__4460 (
            .O(N__20063),
            .I(N__20060));
    CascadeBuf I__4459 (
            .O(N__20060),
            .I(N__20057));
    CascadeMux I__4458 (
            .O(N__20057),
            .I(N__20054));
    CascadeBuf I__4457 (
            .O(N__20054),
            .I(N__20051));
    CascadeMux I__4456 (
            .O(N__20051),
            .I(N__20048));
    CascadeBuf I__4455 (
            .O(N__20048),
            .I(N__20045));
    CascadeMux I__4454 (
            .O(N__20045),
            .I(N__20042));
    CascadeBuf I__4453 (
            .O(N__20042),
            .I(N__20039));
    CascadeMux I__4452 (
            .O(N__20039),
            .I(N__20036));
    CascadeBuf I__4451 (
            .O(N__20036),
            .I(N__20033));
    CascadeMux I__4450 (
            .O(N__20033),
            .I(N__20030));
    CascadeBuf I__4449 (
            .O(N__20030),
            .I(N__20027));
    CascadeMux I__4448 (
            .O(N__20027),
            .I(N__20024));
    CascadeBuf I__4447 (
            .O(N__20024),
            .I(N__20021));
    CascadeMux I__4446 (
            .O(N__20021),
            .I(N__20018));
    CascadeBuf I__4445 (
            .O(N__20018),
            .I(N__20015));
    CascadeMux I__4444 (
            .O(N__20015),
            .I(N__20012));
    InMux I__4443 (
            .O(N__20012),
            .I(N__20008));
    InMux I__4442 (
            .O(N__20011),
            .I(N__20005));
    LocalMux I__4441 (
            .O(N__20008),
            .I(N__20001));
    LocalMux I__4440 (
            .O(N__20005),
            .I(N__19998));
    InMux I__4439 (
            .O(N__20004),
            .I(N__19995));
    Span12Mux_s9_v I__4438 (
            .O(N__20001),
            .I(N__19992));
    Odrv4 I__4437 (
            .O(N__19998),
            .I(M_this_internal_address_qZ0Z_0));
    LocalMux I__4436 (
            .O(N__19995),
            .I(M_this_internal_address_qZ0Z_0));
    Odrv12 I__4435 (
            .O(N__19992),
            .I(M_this_internal_address_qZ0Z_0));
    InMux I__4434 (
            .O(N__19985),
            .I(N__19982));
    LocalMux I__4433 (
            .O(N__19982),
            .I(N__19979));
    Odrv4 I__4432 (
            .O(N__19979),
            .I(M_this_internal_address_q_3_ns_1_1));
    InMux I__4431 (
            .O(N__19976),
            .I(N__19973));
    LocalMux I__4430 (
            .O(N__19973),
            .I(N__19970));
    Span4Mux_h I__4429 (
            .O(N__19970),
            .I(N__19967));
    Odrv4 I__4428 (
            .O(N__19967),
            .I(M_this_internal_address_q_RNO_1Z0Z_1));
    CascadeMux I__4427 (
            .O(N__19964),
            .I(N__19961));
    CascadeBuf I__4426 (
            .O(N__19961),
            .I(N__19958));
    CascadeMux I__4425 (
            .O(N__19958),
            .I(N__19955));
    CascadeBuf I__4424 (
            .O(N__19955),
            .I(N__19952));
    CascadeMux I__4423 (
            .O(N__19952),
            .I(N__19949));
    CascadeBuf I__4422 (
            .O(N__19949),
            .I(N__19946));
    CascadeMux I__4421 (
            .O(N__19946),
            .I(N__19943));
    CascadeBuf I__4420 (
            .O(N__19943),
            .I(N__19940));
    CascadeMux I__4419 (
            .O(N__19940),
            .I(N__19937));
    CascadeBuf I__4418 (
            .O(N__19937),
            .I(N__19934));
    CascadeMux I__4417 (
            .O(N__19934),
            .I(N__19931));
    CascadeBuf I__4416 (
            .O(N__19931),
            .I(N__19928));
    CascadeMux I__4415 (
            .O(N__19928),
            .I(N__19925));
    CascadeBuf I__4414 (
            .O(N__19925),
            .I(N__19922));
    CascadeMux I__4413 (
            .O(N__19922),
            .I(N__19919));
    CascadeBuf I__4412 (
            .O(N__19919),
            .I(N__19916));
    CascadeMux I__4411 (
            .O(N__19916),
            .I(N__19913));
    CascadeBuf I__4410 (
            .O(N__19913),
            .I(N__19910));
    CascadeMux I__4409 (
            .O(N__19910),
            .I(N__19907));
    CascadeBuf I__4408 (
            .O(N__19907),
            .I(N__19904));
    CascadeMux I__4407 (
            .O(N__19904),
            .I(N__19901));
    CascadeBuf I__4406 (
            .O(N__19901),
            .I(N__19898));
    CascadeMux I__4405 (
            .O(N__19898),
            .I(N__19895));
    CascadeBuf I__4404 (
            .O(N__19895),
            .I(N__19892));
    CascadeMux I__4403 (
            .O(N__19892),
            .I(N__19889));
    CascadeBuf I__4402 (
            .O(N__19889),
            .I(N__19886));
    CascadeMux I__4401 (
            .O(N__19886),
            .I(N__19883));
    CascadeBuf I__4400 (
            .O(N__19883),
            .I(N__19880));
    CascadeMux I__4399 (
            .O(N__19880),
            .I(N__19877));
    CascadeBuf I__4398 (
            .O(N__19877),
            .I(N__19874));
    CascadeMux I__4397 (
            .O(N__19874),
            .I(N__19871));
    InMux I__4396 (
            .O(N__19871),
            .I(N__19868));
    LocalMux I__4395 (
            .O(N__19868),
            .I(N__19865));
    Span4Mux_s2_v I__4394 (
            .O(N__19865),
            .I(N__19862));
    Span4Mux_h I__4393 (
            .O(N__19862),
            .I(N__19857));
    InMux I__4392 (
            .O(N__19861),
            .I(N__19854));
    InMux I__4391 (
            .O(N__19860),
            .I(N__19851));
    Span4Mux_h I__4390 (
            .O(N__19857),
            .I(N__19848));
    LocalMux I__4389 (
            .O(N__19854),
            .I(N__19843));
    LocalMux I__4388 (
            .O(N__19851),
            .I(N__19843));
    Span4Mux_v I__4387 (
            .O(N__19848),
            .I(N__19840));
    Odrv4 I__4386 (
            .O(N__19843),
            .I(M_this_internal_address_qZ0Z_1));
    Odrv4 I__4385 (
            .O(N__19840),
            .I(M_this_internal_address_qZ0Z_1));
    InMux I__4384 (
            .O(N__19835),
            .I(N__19832));
    LocalMux I__4383 (
            .O(N__19832),
            .I(N_476));
    InMux I__4382 (
            .O(N__19829),
            .I(N__19825));
    InMux I__4381 (
            .O(N__19828),
            .I(N__19822));
    LocalMux I__4380 (
            .O(N__19825),
            .I(N__19816));
    LocalMux I__4379 (
            .O(N__19822),
            .I(N__19816));
    InMux I__4378 (
            .O(N__19821),
            .I(N__19813));
    Span4Mux_h I__4377 (
            .O(N__19816),
            .I(N__19808));
    LocalMux I__4376 (
            .O(N__19813),
            .I(N__19808));
    Span4Mux_v I__4375 (
            .O(N__19808),
            .I(N__19805));
    Odrv4 I__4374 (
            .O(N__19805),
            .I(N_240));
    CascadeMux I__4373 (
            .O(N__19802),
            .I(N__19795));
    InMux I__4372 (
            .O(N__19801),
            .I(N__19789));
    InMux I__4371 (
            .O(N__19800),
            .I(N__19789));
    InMux I__4370 (
            .O(N__19799),
            .I(N__19786));
    InMux I__4369 (
            .O(N__19798),
            .I(N__19783));
    InMux I__4368 (
            .O(N__19795),
            .I(N__19778));
    InMux I__4367 (
            .O(N__19794),
            .I(N__19778));
    LocalMux I__4366 (
            .O(N__19789),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__4365 (
            .O(N__19786),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__4364 (
            .O(N__19783),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__4363 (
            .O(N__19778),
            .I(M_this_state_qZ0Z_1));
    CascadeMux I__4362 (
            .O(N__19769),
            .I(\this_vga_signals.N_343_cascade_ ));
    InMux I__4361 (
            .O(N__19766),
            .I(N__19763));
    LocalMux I__4360 (
            .O(N__19763),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0));
    InMux I__4359 (
            .O(N__19760),
            .I(N__19757));
    LocalMux I__4358 (
            .O(N__19757),
            .I(N__19751));
    InMux I__4357 (
            .O(N__19756),
            .I(N__19746));
    InMux I__4356 (
            .O(N__19755),
            .I(N__19746));
    InMux I__4355 (
            .O(N__19754),
            .I(N__19743));
    Odrv4 I__4354 (
            .O(N__19751),
            .I(this_ppu_sprites_N_2_1));
    LocalMux I__4353 (
            .O(N__19746),
            .I(this_ppu_sprites_N_2_1));
    LocalMux I__4352 (
            .O(N__19743),
            .I(this_ppu_sprites_N_2_1));
    CascadeMux I__4351 (
            .O(N__19736),
            .I(N__19733));
    CascadeBuf I__4350 (
            .O(N__19733),
            .I(N__19730));
    CascadeMux I__4349 (
            .O(N__19730),
            .I(N__19727));
    CascadeBuf I__4348 (
            .O(N__19727),
            .I(N__19724));
    CascadeMux I__4347 (
            .O(N__19724),
            .I(N__19721));
    CascadeBuf I__4346 (
            .O(N__19721),
            .I(N__19718));
    CascadeMux I__4345 (
            .O(N__19718),
            .I(N__19715));
    CascadeBuf I__4344 (
            .O(N__19715),
            .I(N__19712));
    CascadeMux I__4343 (
            .O(N__19712),
            .I(N__19709));
    CascadeBuf I__4342 (
            .O(N__19709),
            .I(N__19706));
    CascadeMux I__4341 (
            .O(N__19706),
            .I(N__19703));
    CascadeBuf I__4340 (
            .O(N__19703),
            .I(N__19700));
    CascadeMux I__4339 (
            .O(N__19700),
            .I(N__19697));
    CascadeBuf I__4338 (
            .O(N__19697),
            .I(N__19694));
    CascadeMux I__4337 (
            .O(N__19694),
            .I(N__19691));
    CascadeBuf I__4336 (
            .O(N__19691),
            .I(N__19688));
    CascadeMux I__4335 (
            .O(N__19688),
            .I(N__19685));
    CascadeBuf I__4334 (
            .O(N__19685),
            .I(N__19682));
    CascadeMux I__4333 (
            .O(N__19682),
            .I(N__19679));
    CascadeBuf I__4332 (
            .O(N__19679),
            .I(N__19676));
    CascadeMux I__4331 (
            .O(N__19676),
            .I(N__19673));
    CascadeBuf I__4330 (
            .O(N__19673),
            .I(N__19670));
    CascadeMux I__4329 (
            .O(N__19670),
            .I(N__19667));
    CascadeBuf I__4328 (
            .O(N__19667),
            .I(N__19664));
    CascadeMux I__4327 (
            .O(N__19664),
            .I(N__19661));
    CascadeBuf I__4326 (
            .O(N__19661),
            .I(N__19658));
    CascadeMux I__4325 (
            .O(N__19658),
            .I(N__19655));
    CascadeBuf I__4324 (
            .O(N__19655),
            .I(N__19652));
    CascadeMux I__4323 (
            .O(N__19652),
            .I(N__19649));
    CascadeBuf I__4322 (
            .O(N__19649),
            .I(N__19646));
    CascadeMux I__4321 (
            .O(N__19646),
            .I(N__19643));
    InMux I__4320 (
            .O(N__19643),
            .I(N__19640));
    LocalMux I__4319 (
            .O(N__19640),
            .I(N__19637));
    Span12Mux_s10_h I__4318 (
            .O(N__19637),
            .I(N__19634));
    Span12Mux_v I__4317 (
            .O(N__19634),
            .I(N__19631));
    Odrv12 I__4316 (
            .O(N__19631),
            .I(N_134_0));
    InMux I__4315 (
            .O(N__19628),
            .I(N__19625));
    LocalMux I__4314 (
            .O(N__19625),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4 ));
    CascadeMux I__4313 (
            .O(N__19622),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4_cascade_ ));
    InMux I__4312 (
            .O(N__19619),
            .I(N__19616));
    LocalMux I__4311 (
            .O(N__19616),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_1Z0Z_4 ));
    InMux I__4310 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__4309 (
            .O(N__19610),
            .I(\this_vga_signals.M_this_state_q_srsts_0_i_0Z0Z_4 ));
    CascadeMux I__4308 (
            .O(N__19607),
            .I(N__19604));
    InMux I__4307 (
            .O(N__19604),
            .I(N__19601));
    LocalMux I__4306 (
            .O(N__19601),
            .I(\this_vga_signals.N_224_0 ));
    InMux I__4305 (
            .O(N__19598),
            .I(N__19595));
    LocalMux I__4304 (
            .O(N__19595),
            .I(N__19591));
    IoInMux I__4303 (
            .O(N__19594),
            .I(N__19588));
    Span4Mux_v I__4302 (
            .O(N__19591),
            .I(N__19585));
    LocalMux I__4301 (
            .O(N__19588),
            .I(N__19582));
    Span4Mux_v I__4300 (
            .O(N__19585),
            .I(N__19579));
    Span12Mux_s11_v I__4299 (
            .O(N__19582),
            .I(N__19576));
    Odrv4 I__4298 (
            .O(N__19579),
            .I(M_this_state_q_nss_0));
    Odrv12 I__4297 (
            .O(N__19576),
            .I(M_this_state_q_nss_0));
    CascadeMux I__4296 (
            .O(N__19571),
            .I(N__19568));
    InMux I__4295 (
            .O(N__19568),
            .I(N__19564));
    InMux I__4294 (
            .O(N__19567),
            .I(N__19561));
    LocalMux I__4293 (
            .O(N__19564),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__4292 (
            .O(N__19561),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__4291 (
            .O(N__19556),
            .I(N__19552));
    InMux I__4290 (
            .O(N__19555),
            .I(N__19549));
    LocalMux I__4289 (
            .O(N__19552),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__4288 (
            .O(N__19549),
            .I(M_this_data_count_qZ0Z_0));
    CascadeMux I__4287 (
            .O(N__19544),
            .I(N__19541));
    InMux I__4286 (
            .O(N__19541),
            .I(N__19537));
    InMux I__4285 (
            .O(N__19540),
            .I(N__19534));
    LocalMux I__4284 (
            .O(N__19537),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__4283 (
            .O(N__19534),
            .I(M_this_data_count_qZ0Z_11));
    CascadeMux I__4282 (
            .O(N__19529),
            .I(N__19526));
    InMux I__4281 (
            .O(N__19526),
            .I(N__19522));
    InMux I__4280 (
            .O(N__19525),
            .I(N__19519));
    LocalMux I__4279 (
            .O(N__19522),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__4278 (
            .O(N__19519),
            .I(M_this_data_count_qZ0Z_9));
    CascadeMux I__4277 (
            .O(N__19514),
            .I(N__19510));
    InMux I__4276 (
            .O(N__19513),
            .I(N__19507));
    InMux I__4275 (
            .O(N__19510),
            .I(N__19504));
    LocalMux I__4274 (
            .O(N__19507),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__4273 (
            .O(N__19504),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__4272 (
            .O(N__19499),
            .I(N__19495));
    InMux I__4271 (
            .O(N__19498),
            .I(N__19492));
    LocalMux I__4270 (
            .O(N__19495),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__4269 (
            .O(N__19492),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__4268 (
            .O(N__19487),
            .I(N__19483));
    InMux I__4267 (
            .O(N__19486),
            .I(N__19480));
    LocalMux I__4266 (
            .O(N__19483),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__4265 (
            .O(N__19480),
            .I(M_this_data_count_qZ0Z_6));
    CascadeMux I__4264 (
            .O(N__19475),
            .I(N__19472));
    InMux I__4263 (
            .O(N__19472),
            .I(N__19468));
    InMux I__4262 (
            .O(N__19471),
            .I(N__19465));
    LocalMux I__4261 (
            .O(N__19468),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__4260 (
            .O(N__19465),
            .I(M_this_data_count_qZ0Z_5));
    CascadeMux I__4259 (
            .O(N__19460),
            .I(N__19456));
    CascadeMux I__4258 (
            .O(N__19459),
            .I(N__19453));
    InMux I__4257 (
            .O(N__19456),
            .I(N__19450));
    InMux I__4256 (
            .O(N__19453),
            .I(N__19447));
    LocalMux I__4255 (
            .O(N__19450),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__4254 (
            .O(N__19447),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__4253 (
            .O(N__19442),
            .I(N__19438));
    InMux I__4252 (
            .O(N__19441),
            .I(N__19435));
    LocalMux I__4251 (
            .O(N__19438),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__4250 (
            .O(N__19435),
            .I(M_this_data_count_qZ0Z_4));
    CascadeMux I__4249 (
            .O(N__19430),
            .I(N__19427));
    InMux I__4248 (
            .O(N__19427),
            .I(N__19423));
    InMux I__4247 (
            .O(N__19426),
            .I(N__19420));
    LocalMux I__4246 (
            .O(N__19423),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__4245 (
            .O(N__19420),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__4244 (
            .O(N__19415),
            .I(N__19411));
    InMux I__4243 (
            .O(N__19414),
            .I(N__19408));
    LocalMux I__4242 (
            .O(N__19411),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__4241 (
            .O(N__19408),
            .I(M_this_data_count_qZ0Z_2));
    CascadeMux I__4240 (
            .O(N__19403),
            .I(N__19399));
    InMux I__4239 (
            .O(N__19402),
            .I(N__19396));
    InMux I__4238 (
            .O(N__19399),
            .I(N__19393));
    LocalMux I__4237 (
            .O(N__19396),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__4236 (
            .O(N__19393),
            .I(M_this_data_count_qZ0Z_10));
    CascadeMux I__4235 (
            .O(N__19388),
            .I(N__19385));
    InMux I__4234 (
            .O(N__19385),
            .I(N__19381));
    InMux I__4233 (
            .O(N__19384),
            .I(N__19378));
    LocalMux I__4232 (
            .O(N__19381),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__4231 (
            .O(N__19378),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__4230 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__4229 (
            .O(N__19370),
            .I(M_this_state_q_srsts_0_a2_1_9_4));
    InMux I__4228 (
            .O(N__19367),
            .I(N__19364));
    LocalMux I__4227 (
            .O(N__19364),
            .I(M_this_state_q_srsts_0_a2_1_7_4));
    CascadeMux I__4226 (
            .O(N__19361),
            .I(M_this_state_q_srsts_0_a2_1_8_4_cascade_));
    InMux I__4225 (
            .O(N__19358),
            .I(N__19355));
    LocalMux I__4224 (
            .O(N__19355),
            .I(M_this_state_q_srsts_0_a2_1_6_4));
    InMux I__4223 (
            .O(N__19352),
            .I(N__19346));
    InMux I__4222 (
            .O(N__19351),
            .I(N__19346));
    LocalMux I__4221 (
            .O(N__19346),
            .I(N__19341));
    InMux I__4220 (
            .O(N__19345),
            .I(N__19336));
    InMux I__4219 (
            .O(N__19344),
            .I(N__19336));
    Sp12to4 I__4218 (
            .O(N__19341),
            .I(N__19331));
    LocalMux I__4217 (
            .O(N__19336),
            .I(N__19331));
    Span12Mux_v I__4216 (
            .O(N__19331),
            .I(N__19328));
    Odrv12 I__4215 (
            .O(N__19328),
            .I(rst_n_c));
    InMux I__4214 (
            .O(N__19325),
            .I(N__19322));
    LocalMux I__4213 (
            .O(N__19322),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__4212 (
            .O(N__19319),
            .I(N__19316));
    LocalMux I__4211 (
            .O(N__19316),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    CascadeMux I__4210 (
            .O(N__19313),
            .I(N__19310));
    CascadeBuf I__4209 (
            .O(N__19310),
            .I(N__19307));
    CascadeMux I__4208 (
            .O(N__19307),
            .I(N__19304));
    CascadeBuf I__4207 (
            .O(N__19304),
            .I(N__19301));
    CascadeMux I__4206 (
            .O(N__19301),
            .I(N__19298));
    CascadeBuf I__4205 (
            .O(N__19298),
            .I(N__19295));
    CascadeMux I__4204 (
            .O(N__19295),
            .I(N__19292));
    CascadeBuf I__4203 (
            .O(N__19292),
            .I(N__19289));
    CascadeMux I__4202 (
            .O(N__19289),
            .I(N__19286));
    CascadeBuf I__4201 (
            .O(N__19286),
            .I(N__19283));
    CascadeMux I__4200 (
            .O(N__19283),
            .I(N__19280));
    CascadeBuf I__4199 (
            .O(N__19280),
            .I(N__19277));
    CascadeMux I__4198 (
            .O(N__19277),
            .I(N__19274));
    CascadeBuf I__4197 (
            .O(N__19274),
            .I(N__19271));
    CascadeMux I__4196 (
            .O(N__19271),
            .I(N__19268));
    CascadeBuf I__4195 (
            .O(N__19268),
            .I(N__19265));
    CascadeMux I__4194 (
            .O(N__19265),
            .I(N__19262));
    CascadeBuf I__4193 (
            .O(N__19262),
            .I(N__19259));
    CascadeMux I__4192 (
            .O(N__19259),
            .I(N__19256));
    CascadeBuf I__4191 (
            .O(N__19256),
            .I(N__19253));
    CascadeMux I__4190 (
            .O(N__19253),
            .I(N__19250));
    CascadeBuf I__4189 (
            .O(N__19250),
            .I(N__19247));
    CascadeMux I__4188 (
            .O(N__19247),
            .I(N__19244));
    CascadeBuf I__4187 (
            .O(N__19244),
            .I(N__19241));
    CascadeMux I__4186 (
            .O(N__19241),
            .I(N__19238));
    CascadeBuf I__4185 (
            .O(N__19238),
            .I(N__19235));
    CascadeMux I__4184 (
            .O(N__19235),
            .I(N__19232));
    CascadeBuf I__4183 (
            .O(N__19232),
            .I(N__19229));
    CascadeMux I__4182 (
            .O(N__19229),
            .I(N__19226));
    CascadeBuf I__4181 (
            .O(N__19226),
            .I(N__19223));
    CascadeMux I__4180 (
            .O(N__19223),
            .I(N__19220));
    InMux I__4179 (
            .O(N__19220),
            .I(N__19217));
    LocalMux I__4178 (
            .O(N__19217),
            .I(N__19212));
    InMux I__4177 (
            .O(N__19216),
            .I(N__19209));
    InMux I__4176 (
            .O(N__19215),
            .I(N__19206));
    Span12Mux_s11_v I__4175 (
            .O(N__19212),
            .I(N__19203));
    LocalMux I__4174 (
            .O(N__19209),
            .I(M_this_internal_address_qZ0Z_8));
    LocalMux I__4173 (
            .O(N__19206),
            .I(M_this_internal_address_qZ0Z_8));
    Odrv12 I__4172 (
            .O(N__19203),
            .I(M_this_internal_address_qZ0Z_8));
    InMux I__4171 (
            .O(N__19196),
            .I(N__19193));
    LocalMux I__4170 (
            .O(N__19193),
            .I(M_this_internal_address_q_RNO_1Z0Z_8));
    InMux I__4169 (
            .O(N__19190),
            .I(bfn_16_22_0_));
    CascadeMux I__4168 (
            .O(N__19187),
            .I(N__19184));
    CascadeBuf I__4167 (
            .O(N__19184),
            .I(N__19181));
    CascadeMux I__4166 (
            .O(N__19181),
            .I(N__19178));
    CascadeBuf I__4165 (
            .O(N__19178),
            .I(N__19175));
    CascadeMux I__4164 (
            .O(N__19175),
            .I(N__19172));
    CascadeBuf I__4163 (
            .O(N__19172),
            .I(N__19169));
    CascadeMux I__4162 (
            .O(N__19169),
            .I(N__19166));
    CascadeBuf I__4161 (
            .O(N__19166),
            .I(N__19163));
    CascadeMux I__4160 (
            .O(N__19163),
            .I(N__19160));
    CascadeBuf I__4159 (
            .O(N__19160),
            .I(N__19157));
    CascadeMux I__4158 (
            .O(N__19157),
            .I(N__19154));
    CascadeBuf I__4157 (
            .O(N__19154),
            .I(N__19151));
    CascadeMux I__4156 (
            .O(N__19151),
            .I(N__19148));
    CascadeBuf I__4155 (
            .O(N__19148),
            .I(N__19145));
    CascadeMux I__4154 (
            .O(N__19145),
            .I(N__19142));
    CascadeBuf I__4153 (
            .O(N__19142),
            .I(N__19139));
    CascadeMux I__4152 (
            .O(N__19139),
            .I(N__19136));
    CascadeBuf I__4151 (
            .O(N__19136),
            .I(N__19133));
    CascadeMux I__4150 (
            .O(N__19133),
            .I(N__19130));
    CascadeBuf I__4149 (
            .O(N__19130),
            .I(N__19127));
    CascadeMux I__4148 (
            .O(N__19127),
            .I(N__19124));
    CascadeBuf I__4147 (
            .O(N__19124),
            .I(N__19121));
    CascadeMux I__4146 (
            .O(N__19121),
            .I(N__19118));
    CascadeBuf I__4145 (
            .O(N__19118),
            .I(N__19115));
    CascadeMux I__4144 (
            .O(N__19115),
            .I(N__19112));
    CascadeBuf I__4143 (
            .O(N__19112),
            .I(N__19109));
    CascadeMux I__4142 (
            .O(N__19109),
            .I(N__19106));
    CascadeBuf I__4141 (
            .O(N__19106),
            .I(N__19103));
    CascadeMux I__4140 (
            .O(N__19103),
            .I(N__19100));
    CascadeBuf I__4139 (
            .O(N__19100),
            .I(N__19097));
    CascadeMux I__4138 (
            .O(N__19097),
            .I(N__19094));
    InMux I__4137 (
            .O(N__19094),
            .I(N__19090));
    CascadeMux I__4136 (
            .O(N__19093),
            .I(N__19087));
    LocalMux I__4135 (
            .O(N__19090),
            .I(N__19083));
    InMux I__4134 (
            .O(N__19087),
            .I(N__19080));
    InMux I__4133 (
            .O(N__19086),
            .I(N__19077));
    Span12Mux_h I__4132 (
            .O(N__19083),
            .I(N__19074));
    LocalMux I__4131 (
            .O(N__19080),
            .I(M_this_internal_address_qZ0Z_9));
    LocalMux I__4130 (
            .O(N__19077),
            .I(M_this_internal_address_qZ0Z_9));
    Odrv12 I__4129 (
            .O(N__19074),
            .I(M_this_internal_address_qZ0Z_9));
    InMux I__4128 (
            .O(N__19067),
            .I(N__19064));
    LocalMux I__4127 (
            .O(N__19064),
            .I(M_this_internal_address_q_RNO_1Z0Z_9));
    InMux I__4126 (
            .O(N__19061),
            .I(un1_M_this_internal_address_q_cry_8));
    CascadeMux I__4125 (
            .O(N__19058),
            .I(N__19055));
    CascadeBuf I__4124 (
            .O(N__19055),
            .I(N__19052));
    CascadeMux I__4123 (
            .O(N__19052),
            .I(N__19049));
    CascadeBuf I__4122 (
            .O(N__19049),
            .I(N__19046));
    CascadeMux I__4121 (
            .O(N__19046),
            .I(N__19043));
    CascadeBuf I__4120 (
            .O(N__19043),
            .I(N__19040));
    CascadeMux I__4119 (
            .O(N__19040),
            .I(N__19037));
    CascadeBuf I__4118 (
            .O(N__19037),
            .I(N__19034));
    CascadeMux I__4117 (
            .O(N__19034),
            .I(N__19031));
    CascadeBuf I__4116 (
            .O(N__19031),
            .I(N__19028));
    CascadeMux I__4115 (
            .O(N__19028),
            .I(N__19025));
    CascadeBuf I__4114 (
            .O(N__19025),
            .I(N__19022));
    CascadeMux I__4113 (
            .O(N__19022),
            .I(N__19019));
    CascadeBuf I__4112 (
            .O(N__19019),
            .I(N__19016));
    CascadeMux I__4111 (
            .O(N__19016),
            .I(N__19013));
    CascadeBuf I__4110 (
            .O(N__19013),
            .I(N__19010));
    CascadeMux I__4109 (
            .O(N__19010),
            .I(N__19007));
    CascadeBuf I__4108 (
            .O(N__19007),
            .I(N__19004));
    CascadeMux I__4107 (
            .O(N__19004),
            .I(N__19001));
    CascadeBuf I__4106 (
            .O(N__19001),
            .I(N__18998));
    CascadeMux I__4105 (
            .O(N__18998),
            .I(N__18995));
    CascadeBuf I__4104 (
            .O(N__18995),
            .I(N__18992));
    CascadeMux I__4103 (
            .O(N__18992),
            .I(N__18989));
    CascadeBuf I__4102 (
            .O(N__18989),
            .I(N__18986));
    CascadeMux I__4101 (
            .O(N__18986),
            .I(N__18983));
    CascadeBuf I__4100 (
            .O(N__18983),
            .I(N__18980));
    CascadeMux I__4099 (
            .O(N__18980),
            .I(N__18977));
    CascadeBuf I__4098 (
            .O(N__18977),
            .I(N__18974));
    CascadeMux I__4097 (
            .O(N__18974),
            .I(N__18971));
    CascadeBuf I__4096 (
            .O(N__18971),
            .I(N__18968));
    CascadeMux I__4095 (
            .O(N__18968),
            .I(N__18965));
    InMux I__4094 (
            .O(N__18965),
            .I(N__18962));
    LocalMux I__4093 (
            .O(N__18962),
            .I(N__18959));
    Span4Mux_s3_v I__4092 (
            .O(N__18959),
            .I(N__18955));
    InMux I__4091 (
            .O(N__18958),
            .I(N__18952));
    Sp12to4 I__4090 (
            .O(N__18955),
            .I(N__18948));
    LocalMux I__4089 (
            .O(N__18952),
            .I(N__18945));
    InMux I__4088 (
            .O(N__18951),
            .I(N__18942));
    Span12Mux_h I__4087 (
            .O(N__18948),
            .I(N__18939));
    Odrv4 I__4086 (
            .O(N__18945),
            .I(M_this_internal_address_qZ0Z_10));
    LocalMux I__4085 (
            .O(N__18942),
            .I(M_this_internal_address_qZ0Z_10));
    Odrv12 I__4084 (
            .O(N__18939),
            .I(M_this_internal_address_qZ0Z_10));
    InMux I__4083 (
            .O(N__18932),
            .I(N__18929));
    LocalMux I__4082 (
            .O(N__18929),
            .I(N__18926));
    Odrv4 I__4081 (
            .O(N__18926),
            .I(M_this_internal_address_q_RNO_1Z0Z_10));
    InMux I__4080 (
            .O(N__18923),
            .I(un1_M_this_internal_address_q_cry_9));
    InMux I__4079 (
            .O(N__18920),
            .I(un1_M_this_internal_address_q_cry_10));
    InMux I__4078 (
            .O(N__18917),
            .I(un1_M_this_internal_address_q_cry_11));
    InMux I__4077 (
            .O(N__18914),
            .I(un1_M_this_internal_address_q_cry_12));
    InMux I__4076 (
            .O(N__18911),
            .I(N__18908));
    LocalMux I__4075 (
            .O(N__18908),
            .I(N__18905));
    Span4Mux_h I__4074 (
            .O(N__18905),
            .I(N__18902));
    Odrv4 I__4073 (
            .O(N__18902),
            .I(M_this_internal_address_q_RNO_1Z0Z_13));
    CascadeMux I__4072 (
            .O(N__18899),
            .I(N__18896));
    CascadeBuf I__4071 (
            .O(N__18896),
            .I(N__18893));
    CascadeMux I__4070 (
            .O(N__18893),
            .I(N__18890));
    CascadeBuf I__4069 (
            .O(N__18890),
            .I(N__18887));
    CascadeMux I__4068 (
            .O(N__18887),
            .I(N__18884));
    CascadeBuf I__4067 (
            .O(N__18884),
            .I(N__18881));
    CascadeMux I__4066 (
            .O(N__18881),
            .I(N__18878));
    CascadeBuf I__4065 (
            .O(N__18878),
            .I(N__18875));
    CascadeMux I__4064 (
            .O(N__18875),
            .I(N__18872));
    CascadeBuf I__4063 (
            .O(N__18872),
            .I(N__18869));
    CascadeMux I__4062 (
            .O(N__18869),
            .I(N__18866));
    CascadeBuf I__4061 (
            .O(N__18866),
            .I(N__18863));
    CascadeMux I__4060 (
            .O(N__18863),
            .I(N__18860));
    CascadeBuf I__4059 (
            .O(N__18860),
            .I(N__18857));
    CascadeMux I__4058 (
            .O(N__18857),
            .I(N__18854));
    CascadeBuf I__4057 (
            .O(N__18854),
            .I(N__18851));
    CascadeMux I__4056 (
            .O(N__18851),
            .I(N__18848));
    CascadeBuf I__4055 (
            .O(N__18848),
            .I(N__18845));
    CascadeMux I__4054 (
            .O(N__18845),
            .I(N__18842));
    CascadeBuf I__4053 (
            .O(N__18842),
            .I(N__18839));
    CascadeMux I__4052 (
            .O(N__18839),
            .I(N__18836));
    CascadeBuf I__4051 (
            .O(N__18836),
            .I(N__18833));
    CascadeMux I__4050 (
            .O(N__18833),
            .I(N__18830));
    CascadeBuf I__4049 (
            .O(N__18830),
            .I(N__18827));
    CascadeMux I__4048 (
            .O(N__18827),
            .I(N__18824));
    CascadeBuf I__4047 (
            .O(N__18824),
            .I(N__18821));
    CascadeMux I__4046 (
            .O(N__18821),
            .I(N__18818));
    CascadeBuf I__4045 (
            .O(N__18818),
            .I(N__18815));
    CascadeMux I__4044 (
            .O(N__18815),
            .I(N__18812));
    CascadeBuf I__4043 (
            .O(N__18812),
            .I(N__18809));
    CascadeMux I__4042 (
            .O(N__18809),
            .I(N__18805));
    InMux I__4041 (
            .O(N__18808),
            .I(N__18802));
    InMux I__4040 (
            .O(N__18805),
            .I(N__18798));
    LocalMux I__4039 (
            .O(N__18802),
            .I(N__18795));
    InMux I__4038 (
            .O(N__18801),
            .I(N__18792));
    LocalMux I__4037 (
            .O(N__18798),
            .I(N__18789));
    Span4Mux_v I__4036 (
            .O(N__18795),
            .I(N__18784));
    LocalMux I__4035 (
            .O(N__18792),
            .I(N__18784));
    Span12Mux_h I__4034 (
            .O(N__18789),
            .I(N__18781));
    Odrv4 I__4033 (
            .O(N__18784),
            .I(M_this_internal_address_qZ0Z_7));
    Odrv12 I__4032 (
            .O(N__18781),
            .I(M_this_internal_address_qZ0Z_7));
    InMux I__4031 (
            .O(N__18776),
            .I(N__18773));
    LocalMux I__4030 (
            .O(N__18773),
            .I(N__18770));
    Odrv4 I__4029 (
            .O(N__18770),
            .I(M_this_internal_address_q_3_ns_1_7));
    IoInMux I__4028 (
            .O(N__18767),
            .I(N__18763));
    IoInMux I__4027 (
            .O(N__18766),
            .I(N__18760));
    LocalMux I__4026 (
            .O(N__18763),
            .I(N__18753));
    LocalMux I__4025 (
            .O(N__18760),
            .I(N__18753));
    IoInMux I__4024 (
            .O(N__18759),
            .I(N__18750));
    IoInMux I__4023 (
            .O(N__18758),
            .I(N__18745));
    IoSpan4Mux I__4022 (
            .O(N__18753),
            .I(N__18742));
    LocalMux I__4021 (
            .O(N__18750),
            .I(N__18736));
    IoInMux I__4020 (
            .O(N__18749),
            .I(N__18733));
    IoInMux I__4019 (
            .O(N__18748),
            .I(N__18730));
    LocalMux I__4018 (
            .O(N__18745),
            .I(N__18726));
    IoSpan4Mux I__4017 (
            .O(N__18742),
            .I(N__18723));
    IoInMux I__4016 (
            .O(N__18741),
            .I(N__18720));
    IoInMux I__4015 (
            .O(N__18740),
            .I(N__18717));
    IoInMux I__4014 (
            .O(N__18739),
            .I(N__18711));
    IoSpan4Mux I__4013 (
            .O(N__18736),
            .I(N__18704));
    LocalMux I__4012 (
            .O(N__18733),
            .I(N__18704));
    LocalMux I__4011 (
            .O(N__18730),
            .I(N__18704));
    IoInMux I__4010 (
            .O(N__18729),
            .I(N__18701));
    IoSpan4Mux I__4009 (
            .O(N__18726),
            .I(N__18698));
    IoSpan4Mux I__4008 (
            .O(N__18723),
            .I(N__18691));
    LocalMux I__4007 (
            .O(N__18720),
            .I(N__18691));
    LocalMux I__4006 (
            .O(N__18717),
            .I(N__18691));
    IoInMux I__4005 (
            .O(N__18716),
            .I(N__18688));
    IoInMux I__4004 (
            .O(N__18715),
            .I(N__18685));
    IoInMux I__4003 (
            .O(N__18714),
            .I(N__18682));
    LocalMux I__4002 (
            .O(N__18711),
            .I(N__18679));
    IoSpan4Mux I__4001 (
            .O(N__18704),
            .I(N__18674));
    LocalMux I__4000 (
            .O(N__18701),
            .I(N__18674));
    Span4Mux_s3_h I__3999 (
            .O(N__18698),
            .I(N__18670));
    IoSpan4Mux I__3998 (
            .O(N__18691),
            .I(N__18663));
    LocalMux I__3997 (
            .O(N__18688),
            .I(N__18663));
    LocalMux I__3996 (
            .O(N__18685),
            .I(N__18663));
    LocalMux I__3995 (
            .O(N__18682),
            .I(N__18660));
    Span4Mux_s3_h I__3994 (
            .O(N__18679),
            .I(N__18657));
    IoSpan4Mux I__3993 (
            .O(N__18674),
            .I(N__18654));
    IoInMux I__3992 (
            .O(N__18673),
            .I(N__18650));
    Span4Mux_v I__3991 (
            .O(N__18670),
            .I(N__18643));
    IoSpan4Mux I__3990 (
            .O(N__18663),
            .I(N__18643));
    IoSpan4Mux I__3989 (
            .O(N__18660),
            .I(N__18643));
    Sp12to4 I__3988 (
            .O(N__18657),
            .I(N__18639));
    Span4Mux_s1_v I__3987 (
            .O(N__18654),
            .I(N__18635));
    IoInMux I__3986 (
            .O(N__18653),
            .I(N__18632));
    LocalMux I__3985 (
            .O(N__18650),
            .I(N__18629));
    Span4Mux_s3_h I__3984 (
            .O(N__18643),
            .I(N__18626));
    IoInMux I__3983 (
            .O(N__18642),
            .I(N__18623));
    Span12Mux_s9_v I__3982 (
            .O(N__18639),
            .I(N__18620));
    IoInMux I__3981 (
            .O(N__18638),
            .I(N__18617));
    Sp12to4 I__3980 (
            .O(N__18635),
            .I(N__18612));
    LocalMux I__3979 (
            .O(N__18632),
            .I(N__18612));
    Span4Mux_s2_v I__3978 (
            .O(N__18629),
            .I(N__18609));
    Span4Mux_h I__3977 (
            .O(N__18626),
            .I(N__18606));
    LocalMux I__3976 (
            .O(N__18623),
            .I(N__18603));
    Span12Mux_h I__3975 (
            .O(N__18620),
            .I(N__18598));
    LocalMux I__3974 (
            .O(N__18617),
            .I(N__18598));
    Span12Mux_s9_v I__3973 (
            .O(N__18612),
            .I(N__18595));
    Span4Mux_v I__3972 (
            .O(N__18609),
            .I(N__18592));
    Sp12to4 I__3971 (
            .O(N__18606),
            .I(N__18585));
    Span12Mux_s4_h I__3970 (
            .O(N__18603),
            .I(N__18585));
    Span12Mux_s9_v I__3969 (
            .O(N__18598),
            .I(N__18585));
    Odrv12 I__3968 (
            .O(N__18595),
            .I(N_235_0_i));
    Odrv4 I__3967 (
            .O(N__18592),
            .I(N_235_0_i));
    Odrv12 I__3966 (
            .O(N__18585),
            .I(N_235_0_i));
    InMux I__3965 (
            .O(N__18578),
            .I(un1_M_this_internal_address_q_cry_0));
    CascadeMux I__3964 (
            .O(N__18575),
            .I(N__18572));
    CascadeBuf I__3963 (
            .O(N__18572),
            .I(N__18569));
    CascadeMux I__3962 (
            .O(N__18569),
            .I(N__18566));
    CascadeBuf I__3961 (
            .O(N__18566),
            .I(N__18563));
    CascadeMux I__3960 (
            .O(N__18563),
            .I(N__18560));
    CascadeBuf I__3959 (
            .O(N__18560),
            .I(N__18557));
    CascadeMux I__3958 (
            .O(N__18557),
            .I(N__18554));
    CascadeBuf I__3957 (
            .O(N__18554),
            .I(N__18551));
    CascadeMux I__3956 (
            .O(N__18551),
            .I(N__18548));
    CascadeBuf I__3955 (
            .O(N__18548),
            .I(N__18545));
    CascadeMux I__3954 (
            .O(N__18545),
            .I(N__18542));
    CascadeBuf I__3953 (
            .O(N__18542),
            .I(N__18539));
    CascadeMux I__3952 (
            .O(N__18539),
            .I(N__18536));
    CascadeBuf I__3951 (
            .O(N__18536),
            .I(N__18533));
    CascadeMux I__3950 (
            .O(N__18533),
            .I(N__18530));
    CascadeBuf I__3949 (
            .O(N__18530),
            .I(N__18527));
    CascadeMux I__3948 (
            .O(N__18527),
            .I(N__18524));
    CascadeBuf I__3947 (
            .O(N__18524),
            .I(N__18521));
    CascadeMux I__3946 (
            .O(N__18521),
            .I(N__18518));
    CascadeBuf I__3945 (
            .O(N__18518),
            .I(N__18515));
    CascadeMux I__3944 (
            .O(N__18515),
            .I(N__18512));
    CascadeBuf I__3943 (
            .O(N__18512),
            .I(N__18509));
    CascadeMux I__3942 (
            .O(N__18509),
            .I(N__18506));
    CascadeBuf I__3941 (
            .O(N__18506),
            .I(N__18503));
    CascadeMux I__3940 (
            .O(N__18503),
            .I(N__18500));
    CascadeBuf I__3939 (
            .O(N__18500),
            .I(N__18497));
    CascadeMux I__3938 (
            .O(N__18497),
            .I(N__18494));
    CascadeBuf I__3937 (
            .O(N__18494),
            .I(N__18491));
    CascadeMux I__3936 (
            .O(N__18491),
            .I(N__18488));
    CascadeBuf I__3935 (
            .O(N__18488),
            .I(N__18485));
    CascadeMux I__3934 (
            .O(N__18485),
            .I(N__18482));
    InMux I__3933 (
            .O(N__18482),
            .I(N__18479));
    LocalMux I__3932 (
            .O(N__18479),
            .I(N__18476));
    Span4Mux_h I__3931 (
            .O(N__18476),
            .I(N__18473));
    Sp12to4 I__3930 (
            .O(N__18473),
            .I(N__18468));
    InMux I__3929 (
            .O(N__18472),
            .I(N__18465));
    InMux I__3928 (
            .O(N__18471),
            .I(N__18462));
    Span12Mux_s11_v I__3927 (
            .O(N__18468),
            .I(N__18459));
    LocalMux I__3926 (
            .O(N__18465),
            .I(M_this_internal_address_qZ0Z_2));
    LocalMux I__3925 (
            .O(N__18462),
            .I(M_this_internal_address_qZ0Z_2));
    Odrv12 I__3924 (
            .O(N__18459),
            .I(M_this_internal_address_qZ0Z_2));
    InMux I__3923 (
            .O(N__18452),
            .I(N__18449));
    LocalMux I__3922 (
            .O(N__18449),
            .I(M_this_internal_address_q_RNO_1Z0Z_2));
    InMux I__3921 (
            .O(N__18446),
            .I(un1_M_this_internal_address_q_cry_1));
    CascadeMux I__3920 (
            .O(N__18443),
            .I(N__18440));
    CascadeBuf I__3919 (
            .O(N__18440),
            .I(N__18437));
    CascadeMux I__3918 (
            .O(N__18437),
            .I(N__18434));
    CascadeBuf I__3917 (
            .O(N__18434),
            .I(N__18431));
    CascadeMux I__3916 (
            .O(N__18431),
            .I(N__18428));
    CascadeBuf I__3915 (
            .O(N__18428),
            .I(N__18425));
    CascadeMux I__3914 (
            .O(N__18425),
            .I(N__18422));
    CascadeBuf I__3913 (
            .O(N__18422),
            .I(N__18419));
    CascadeMux I__3912 (
            .O(N__18419),
            .I(N__18416));
    CascadeBuf I__3911 (
            .O(N__18416),
            .I(N__18413));
    CascadeMux I__3910 (
            .O(N__18413),
            .I(N__18410));
    CascadeBuf I__3909 (
            .O(N__18410),
            .I(N__18407));
    CascadeMux I__3908 (
            .O(N__18407),
            .I(N__18404));
    CascadeBuf I__3907 (
            .O(N__18404),
            .I(N__18401));
    CascadeMux I__3906 (
            .O(N__18401),
            .I(N__18398));
    CascadeBuf I__3905 (
            .O(N__18398),
            .I(N__18395));
    CascadeMux I__3904 (
            .O(N__18395),
            .I(N__18392));
    CascadeBuf I__3903 (
            .O(N__18392),
            .I(N__18389));
    CascadeMux I__3902 (
            .O(N__18389),
            .I(N__18386));
    CascadeBuf I__3901 (
            .O(N__18386),
            .I(N__18383));
    CascadeMux I__3900 (
            .O(N__18383),
            .I(N__18380));
    CascadeBuf I__3899 (
            .O(N__18380),
            .I(N__18377));
    CascadeMux I__3898 (
            .O(N__18377),
            .I(N__18374));
    CascadeBuf I__3897 (
            .O(N__18374),
            .I(N__18371));
    CascadeMux I__3896 (
            .O(N__18371),
            .I(N__18368));
    CascadeBuf I__3895 (
            .O(N__18368),
            .I(N__18365));
    CascadeMux I__3894 (
            .O(N__18365),
            .I(N__18362));
    CascadeBuf I__3893 (
            .O(N__18362),
            .I(N__18359));
    CascadeMux I__3892 (
            .O(N__18359),
            .I(N__18356));
    CascadeBuf I__3891 (
            .O(N__18356),
            .I(N__18353));
    CascadeMux I__3890 (
            .O(N__18353),
            .I(N__18350));
    InMux I__3889 (
            .O(N__18350),
            .I(N__18347));
    LocalMux I__3888 (
            .O(N__18347),
            .I(N__18343));
    InMux I__3887 (
            .O(N__18346),
            .I(N__18339));
    Sp12to4 I__3886 (
            .O(N__18343),
            .I(N__18336));
    InMux I__3885 (
            .O(N__18342),
            .I(N__18333));
    LocalMux I__3884 (
            .O(N__18339),
            .I(N__18328));
    Span12Mux_s11_v I__3883 (
            .O(N__18336),
            .I(N__18328));
    LocalMux I__3882 (
            .O(N__18333),
            .I(M_this_internal_address_qZ0Z_3));
    Odrv12 I__3881 (
            .O(N__18328),
            .I(M_this_internal_address_qZ0Z_3));
    InMux I__3880 (
            .O(N__18323),
            .I(N__18320));
    LocalMux I__3879 (
            .O(N__18320),
            .I(M_this_internal_address_q_RNO_1Z0Z_3));
    InMux I__3878 (
            .O(N__18317),
            .I(un1_M_this_internal_address_q_cry_2));
    InMux I__3877 (
            .O(N__18314),
            .I(un1_M_this_internal_address_q_cry_3));
    InMux I__3876 (
            .O(N__18311),
            .I(un1_M_this_internal_address_q_cry_4));
    InMux I__3875 (
            .O(N__18308),
            .I(un1_M_this_internal_address_q_cry_5));
    InMux I__3874 (
            .O(N__18305),
            .I(N__18302));
    LocalMux I__3873 (
            .O(N__18302),
            .I(N__18299));
    Span4Mux_h I__3872 (
            .O(N__18299),
            .I(N__18296));
    Odrv4 I__3871 (
            .O(N__18296),
            .I(M_this_internal_address_q_RNO_1Z0Z_7));
    InMux I__3870 (
            .O(N__18293),
            .I(un1_M_this_internal_address_q_cry_6));
    CascadeMux I__3869 (
            .O(N__18290),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0_cascade_));
    InMux I__3868 (
            .O(N__18287),
            .I(N__18282));
    InMux I__3867 (
            .O(N__18286),
            .I(N__18277));
    InMux I__3866 (
            .O(N__18285),
            .I(N__18277));
    LocalMux I__3865 (
            .O(N__18282),
            .I(if_generate_plus_mult1_un89_sum_axbxc3));
    LocalMux I__3864 (
            .O(N__18277),
            .I(if_generate_plus_mult1_un89_sum_axbxc3));
    CascadeMux I__3863 (
            .O(N__18272),
            .I(\this_ppu.sprites_N_7_0_cascade_ ));
    InMux I__3862 (
            .O(N__18269),
            .I(N__18265));
    InMux I__3861 (
            .O(N__18268),
            .I(N__18262));
    LocalMux I__3860 (
            .O(N__18265),
            .I(\this_ppu.un5_sprites_addr_1_c2 ));
    LocalMux I__3859 (
            .O(N__18262),
            .I(\this_ppu.un5_sprites_addr_1_c2 ));
    CascadeMux I__3858 (
            .O(N__18257),
            .I(\this_ppu.sprites_m7Z0Z_0_cascade_ ));
    InMux I__3857 (
            .O(N__18254),
            .I(N__18251));
    LocalMux I__3856 (
            .O(N__18251),
            .I(N__18241));
    InMux I__3855 (
            .O(N__18250),
            .I(N__18232));
    InMux I__3854 (
            .O(N__18249),
            .I(N__18232));
    InMux I__3853 (
            .O(N__18248),
            .I(N__18232));
    InMux I__3852 (
            .O(N__18247),
            .I(N__18232));
    InMux I__3851 (
            .O(N__18246),
            .I(N__18229));
    InMux I__3850 (
            .O(N__18245),
            .I(N__18224));
    InMux I__3849 (
            .O(N__18244),
            .I(N__18224));
    Odrv4 I__3848 (
            .O(N__18241),
            .I(if_generate_plus_mult1_un68_sum_axbxc3_ns));
    LocalMux I__3847 (
            .O(N__18232),
            .I(if_generate_plus_mult1_un68_sum_axbxc3_ns));
    LocalMux I__3846 (
            .O(N__18229),
            .I(if_generate_plus_mult1_un68_sum_axbxc3_ns));
    LocalMux I__3845 (
            .O(N__18224),
            .I(if_generate_plus_mult1_un68_sum_axbxc3_ns));
    CascadeMux I__3844 (
            .O(N__18215),
            .I(N__18212));
    CascadeBuf I__3843 (
            .O(N__18212),
            .I(N__18209));
    CascadeMux I__3842 (
            .O(N__18209),
            .I(N__18206));
    CascadeBuf I__3841 (
            .O(N__18206),
            .I(N__18203));
    CascadeMux I__3840 (
            .O(N__18203),
            .I(N__18200));
    CascadeBuf I__3839 (
            .O(N__18200),
            .I(N__18197));
    CascadeMux I__3838 (
            .O(N__18197),
            .I(N__18194));
    CascadeBuf I__3837 (
            .O(N__18194),
            .I(N__18191));
    CascadeMux I__3836 (
            .O(N__18191),
            .I(N__18188));
    CascadeBuf I__3835 (
            .O(N__18188),
            .I(N__18185));
    CascadeMux I__3834 (
            .O(N__18185),
            .I(N__18182));
    CascadeBuf I__3833 (
            .O(N__18182),
            .I(N__18179));
    CascadeMux I__3832 (
            .O(N__18179),
            .I(N__18176));
    CascadeBuf I__3831 (
            .O(N__18176),
            .I(N__18173));
    CascadeMux I__3830 (
            .O(N__18173),
            .I(N__18170));
    CascadeBuf I__3829 (
            .O(N__18170),
            .I(N__18167));
    CascadeMux I__3828 (
            .O(N__18167),
            .I(N__18164));
    CascadeBuf I__3827 (
            .O(N__18164),
            .I(N__18161));
    CascadeMux I__3826 (
            .O(N__18161),
            .I(N__18158));
    CascadeBuf I__3825 (
            .O(N__18158),
            .I(N__18155));
    CascadeMux I__3824 (
            .O(N__18155),
            .I(N__18152));
    CascadeBuf I__3823 (
            .O(N__18152),
            .I(N__18149));
    CascadeMux I__3822 (
            .O(N__18149),
            .I(N__18146));
    CascadeBuf I__3821 (
            .O(N__18146),
            .I(N__18143));
    CascadeMux I__3820 (
            .O(N__18143),
            .I(N__18140));
    CascadeBuf I__3819 (
            .O(N__18140),
            .I(N__18137));
    CascadeMux I__3818 (
            .O(N__18137),
            .I(N__18134));
    CascadeBuf I__3817 (
            .O(N__18134),
            .I(N__18131));
    CascadeMux I__3816 (
            .O(N__18131),
            .I(N__18128));
    CascadeBuf I__3815 (
            .O(N__18128),
            .I(N__18125));
    CascadeMux I__3814 (
            .O(N__18125),
            .I(N__18122));
    InMux I__3813 (
            .O(N__18122),
            .I(N__18119));
    LocalMux I__3812 (
            .O(N__18119),
            .I(N__18116));
    Span12Mux_s10_h I__3811 (
            .O(N__18116),
            .I(N__18113));
    Span12Mux_v I__3810 (
            .O(N__18113),
            .I(N__18110));
    Odrv12 I__3809 (
            .O(N__18110),
            .I(N_140_i));
    CascadeMux I__3808 (
            .O(N__18107),
            .I(N__18102));
    InMux I__3807 (
            .O(N__18106),
            .I(N__18094));
    InMux I__3806 (
            .O(N__18105),
            .I(N__18090));
    InMux I__3805 (
            .O(N__18102),
            .I(N__18087));
    CascadeMux I__3804 (
            .O(N__18101),
            .I(N__18084));
    InMux I__3803 (
            .O(N__18100),
            .I(N__18079));
    InMux I__3802 (
            .O(N__18099),
            .I(N__18076));
    InMux I__3801 (
            .O(N__18098),
            .I(N__18071));
    InMux I__3800 (
            .O(N__18097),
            .I(N__18071));
    LocalMux I__3799 (
            .O(N__18094),
            .I(N__18068));
    CascadeMux I__3798 (
            .O(N__18093),
            .I(N__18063));
    LocalMux I__3797 (
            .O(N__18090),
            .I(N__18057));
    LocalMux I__3796 (
            .O(N__18087),
            .I(N__18057));
    InMux I__3795 (
            .O(N__18084),
            .I(N__18054));
    InMux I__3794 (
            .O(N__18083),
            .I(N__18049));
    InMux I__3793 (
            .O(N__18082),
            .I(N__18049));
    LocalMux I__3792 (
            .O(N__18079),
            .I(N__18046));
    LocalMux I__3791 (
            .O(N__18076),
            .I(N__18041));
    LocalMux I__3790 (
            .O(N__18071),
            .I(N__18041));
    Span12Mux_v I__3789 (
            .O(N__18068),
            .I(N__18038));
    InMux I__3788 (
            .O(N__18067),
            .I(N__18035));
    InMux I__3787 (
            .O(N__18066),
            .I(N__18032));
    InMux I__3786 (
            .O(N__18063),
            .I(N__18027));
    InMux I__3785 (
            .O(N__18062),
            .I(N__18027));
    Span4Mux_v I__3784 (
            .O(N__18057),
            .I(N__18024));
    LocalMux I__3783 (
            .O(N__18054),
            .I(N__18021));
    LocalMux I__3782 (
            .O(N__18049),
            .I(N__18018));
    Span4Mux_v I__3781 (
            .O(N__18046),
            .I(N__18013));
    Span4Mux_h I__3780 (
            .O(N__18041),
            .I(N__18013));
    Odrv12 I__3779 (
            .O(N__18038),
            .I(this_vga_signals_M_hcounter_q_2));
    LocalMux I__3778 (
            .O(N__18035),
            .I(this_vga_signals_M_hcounter_q_2));
    LocalMux I__3777 (
            .O(N__18032),
            .I(this_vga_signals_M_hcounter_q_2));
    LocalMux I__3776 (
            .O(N__18027),
            .I(this_vga_signals_M_hcounter_q_2));
    Odrv4 I__3775 (
            .O(N__18024),
            .I(this_vga_signals_M_hcounter_q_2));
    Odrv4 I__3774 (
            .O(N__18021),
            .I(this_vga_signals_M_hcounter_q_2));
    Odrv12 I__3773 (
            .O(N__18018),
            .I(this_vga_signals_M_hcounter_q_2));
    Odrv4 I__3772 (
            .O(N__18013),
            .I(this_vga_signals_M_hcounter_q_2));
    InMux I__3771 (
            .O(N__17996),
            .I(N__17989));
    InMux I__3770 (
            .O(N__17995),
            .I(N__17989));
    InMux I__3769 (
            .O(N__17994),
            .I(N__17986));
    LocalMux I__3768 (
            .O(N__17989),
            .I(N__17983));
    LocalMux I__3767 (
            .O(N__17986),
            .I(N__17980));
    Span4Mux_v I__3766 (
            .O(N__17983),
            .I(N__17974));
    Span4Mux_h I__3765 (
            .O(N__17980),
            .I(N__17974));
    InMux I__3764 (
            .O(N__17979),
            .I(N__17971));
    Odrv4 I__3763 (
            .O(N__17974),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1));
    LocalMux I__3762 (
            .O(N__17971),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1));
    InMux I__3761 (
            .O(N__17966),
            .I(N__17962));
    InMux I__3760 (
            .O(N__17965),
            .I(N__17959));
    LocalMux I__3759 (
            .O(N__17962),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3));
    LocalMux I__3758 (
            .O(N__17959),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3));
    InMux I__3757 (
            .O(N__17954),
            .I(N__17946));
    InMux I__3756 (
            .O(N__17953),
            .I(N__17946));
    InMux I__3755 (
            .O(N__17952),
            .I(N__17941));
    InMux I__3754 (
            .O(N__17951),
            .I(N__17941));
    LocalMux I__3753 (
            .O(N__17946),
            .I(if_generate_plus_mult1_un75_sum_axbxc3));
    LocalMux I__3752 (
            .O(N__17941),
            .I(if_generate_plus_mult1_un75_sum_axbxc3));
    InMux I__3751 (
            .O(N__17936),
            .I(N__17930));
    InMux I__3750 (
            .O(N__17935),
            .I(N__17920));
    InMux I__3749 (
            .O(N__17934),
            .I(N__17920));
    InMux I__3748 (
            .O(N__17933),
            .I(N__17920));
    LocalMux I__3747 (
            .O(N__17930),
            .I(N__17917));
    InMux I__3746 (
            .O(N__17929),
            .I(N__17910));
    InMux I__3745 (
            .O(N__17928),
            .I(N__17910));
    InMux I__3744 (
            .O(N__17927),
            .I(N__17910));
    LocalMux I__3743 (
            .O(N__17920),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0));
    Odrv4 I__3742 (
            .O(N__17917),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0));
    LocalMux I__3741 (
            .O(N__17910),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0));
    InMux I__3740 (
            .O(N__17903),
            .I(N__17898));
    CascadeMux I__3739 (
            .O(N__17902),
            .I(N__17893));
    InMux I__3738 (
            .O(N__17901),
            .I(N__17890));
    LocalMux I__3737 (
            .O(N__17898),
            .I(N__17885));
    InMux I__3736 (
            .O(N__17897),
            .I(N__17882));
    InMux I__3735 (
            .O(N__17896),
            .I(N__17878));
    InMux I__3734 (
            .O(N__17893),
            .I(N__17875));
    LocalMux I__3733 (
            .O(N__17890),
            .I(N__17872));
    CascadeMux I__3732 (
            .O(N__17889),
            .I(N__17866));
    InMux I__3731 (
            .O(N__17888),
            .I(N__17862));
    Span4Mux_h I__3730 (
            .O(N__17885),
            .I(N__17859));
    LocalMux I__3729 (
            .O(N__17882),
            .I(N__17856));
    InMux I__3728 (
            .O(N__17881),
            .I(N__17853));
    LocalMux I__3727 (
            .O(N__17878),
            .I(N__17848));
    LocalMux I__3726 (
            .O(N__17875),
            .I(N__17848));
    Span4Mux_h I__3725 (
            .O(N__17872),
            .I(N__17845));
    InMux I__3724 (
            .O(N__17871),
            .I(N__17842));
    InMux I__3723 (
            .O(N__17870),
            .I(N__17839));
    InMux I__3722 (
            .O(N__17869),
            .I(N__17832));
    InMux I__3721 (
            .O(N__17866),
            .I(N__17832));
    InMux I__3720 (
            .O(N__17865),
            .I(N__17832));
    LocalMux I__3719 (
            .O(N__17862),
            .I(N__17829));
    Span4Mux_v I__3718 (
            .O(N__17859),
            .I(N__17820));
    Span4Mux_h I__3717 (
            .O(N__17856),
            .I(N__17820));
    LocalMux I__3716 (
            .O(N__17853),
            .I(N__17820));
    Span4Mux_h I__3715 (
            .O(N__17848),
            .I(N__17820));
    Odrv4 I__3714 (
            .O(N__17845),
            .I(this_vga_signals_M_hcounter_q_1));
    LocalMux I__3713 (
            .O(N__17842),
            .I(this_vga_signals_M_hcounter_q_1));
    LocalMux I__3712 (
            .O(N__17839),
            .I(this_vga_signals_M_hcounter_q_1));
    LocalMux I__3711 (
            .O(N__17832),
            .I(this_vga_signals_M_hcounter_q_1));
    Odrv12 I__3710 (
            .O(N__17829),
            .I(this_vga_signals_M_hcounter_q_1));
    Odrv4 I__3709 (
            .O(N__17820),
            .I(this_vga_signals_M_hcounter_q_1));
    CascadeMux I__3708 (
            .O(N__17807),
            .I(N__17804));
    InMux I__3707 (
            .O(N__17804),
            .I(N__17796));
    InMux I__3706 (
            .O(N__17803),
            .I(N__17792));
    CascadeMux I__3705 (
            .O(N__17802),
            .I(N__17789));
    InMux I__3704 (
            .O(N__17801),
            .I(N__17785));
    CascadeMux I__3703 (
            .O(N__17800),
            .I(N__17782));
    InMux I__3702 (
            .O(N__17799),
            .I(N__17779));
    LocalMux I__3701 (
            .O(N__17796),
            .I(N__17776));
    CascadeMux I__3700 (
            .O(N__17795),
            .I(N__17770));
    LocalMux I__3699 (
            .O(N__17792),
            .I(N__17767));
    InMux I__3698 (
            .O(N__17789),
            .I(N__17762));
    InMux I__3697 (
            .O(N__17788),
            .I(N__17762));
    LocalMux I__3696 (
            .O(N__17785),
            .I(N__17759));
    InMux I__3695 (
            .O(N__17782),
            .I(N__17756));
    LocalMux I__3694 (
            .O(N__17779),
            .I(N__17751));
    Span4Mux_v I__3693 (
            .O(N__17776),
            .I(N__17751));
    InMux I__3692 (
            .O(N__17775),
            .I(N__17746));
    InMux I__3691 (
            .O(N__17774),
            .I(N__17746));
    InMux I__3690 (
            .O(N__17773),
            .I(N__17743));
    InMux I__3689 (
            .O(N__17770),
            .I(N__17740));
    Span4Mux_h I__3688 (
            .O(N__17767),
            .I(N__17735));
    LocalMux I__3687 (
            .O(N__17762),
            .I(N__17735));
    Span4Mux_v I__3686 (
            .O(N__17759),
            .I(N__17728));
    LocalMux I__3685 (
            .O(N__17756),
            .I(N__17728));
    Span4Mux_h I__3684 (
            .O(N__17751),
            .I(N__17728));
    LocalMux I__3683 (
            .O(N__17746),
            .I(this_vga_signals_M_hcounter_q_0));
    LocalMux I__3682 (
            .O(N__17743),
            .I(this_vga_signals_M_hcounter_q_0));
    LocalMux I__3681 (
            .O(N__17740),
            .I(this_vga_signals_M_hcounter_q_0));
    Odrv4 I__3680 (
            .O(N__17735),
            .I(this_vga_signals_M_hcounter_q_0));
    Odrv4 I__3679 (
            .O(N__17728),
            .I(this_vga_signals_M_hcounter_q_0));
    CascadeMux I__3678 (
            .O(N__17717),
            .I(\this_ppu.sprites_mZ0Z1_cascade_ ));
    InMux I__3677 (
            .O(N__17714),
            .I(N__17709));
    InMux I__3676 (
            .O(N__17713),
            .I(N__17704));
    InMux I__3675 (
            .O(N__17712),
            .I(N__17704));
    LocalMux I__3674 (
            .O(N__17709),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1));
    LocalMux I__3673 (
            .O(N__17704),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1));
    CascadeMux I__3672 (
            .O(N__17699),
            .I(M_this_internal_address_q_3_ns_1_10_cascade_));
    SRMux I__3671 (
            .O(N__17696),
            .I(N__17692));
    SRMux I__3670 (
            .O(N__17695),
            .I(N__17689));
    LocalMux I__3669 (
            .O(N__17692),
            .I(N__17686));
    LocalMux I__3668 (
            .O(N__17689),
            .I(N__17683));
    Span4Mux_h I__3667 (
            .O(N__17686),
            .I(N__17680));
    Odrv4 I__3666 (
            .O(N__17683),
            .I(M_this_state_q_RNI20CEZ0Z_0));
    Odrv4 I__3665 (
            .O(N__17680),
            .I(M_this_state_q_RNI20CEZ0Z_0));
    SRMux I__3664 (
            .O(N__17675),
            .I(N__17668));
    SRMux I__3663 (
            .O(N__17674),
            .I(N__17665));
    SRMux I__3662 (
            .O(N__17673),
            .I(N__17662));
    SRMux I__3661 (
            .O(N__17672),
            .I(N__17655));
    SRMux I__3660 (
            .O(N__17671),
            .I(N__17652));
    LocalMux I__3659 (
            .O(N__17668),
            .I(N__17649));
    LocalMux I__3658 (
            .O(N__17665),
            .I(N__17644));
    LocalMux I__3657 (
            .O(N__17662),
            .I(N__17644));
    SRMux I__3656 (
            .O(N__17661),
            .I(N__17641));
    SRMux I__3655 (
            .O(N__17660),
            .I(N__17638));
    SRMux I__3654 (
            .O(N__17659),
            .I(N__17632));
    SRMux I__3653 (
            .O(N__17658),
            .I(N__17626));
    LocalMux I__3652 (
            .O(N__17655),
            .I(N__17623));
    LocalMux I__3651 (
            .O(N__17652),
            .I(N__17620));
    Span4Mux_h I__3650 (
            .O(N__17649),
            .I(N__17611));
    Span4Mux_s3_v I__3649 (
            .O(N__17644),
            .I(N__17611));
    LocalMux I__3648 (
            .O(N__17641),
            .I(N__17611));
    LocalMux I__3647 (
            .O(N__17638),
            .I(N__17611));
    SRMux I__3646 (
            .O(N__17637),
            .I(N__17608));
    SRMux I__3645 (
            .O(N__17636),
            .I(N__17605));
    SRMux I__3644 (
            .O(N__17635),
            .I(N__17599));
    LocalMux I__3643 (
            .O(N__17632),
            .I(N__17595));
    SRMux I__3642 (
            .O(N__17631),
            .I(N__17592));
    SRMux I__3641 (
            .O(N__17630),
            .I(N__17586));
    SRMux I__3640 (
            .O(N__17629),
            .I(N__17581));
    LocalMux I__3639 (
            .O(N__17626),
            .I(N__17578));
    Span4Mux_v I__3638 (
            .O(N__17623),
            .I(N__17567));
    Span4Mux_h I__3637 (
            .O(N__17620),
            .I(N__17567));
    Span4Mux_v I__3636 (
            .O(N__17611),
            .I(N__17567));
    LocalMux I__3635 (
            .O(N__17608),
            .I(N__17567));
    LocalMux I__3634 (
            .O(N__17605),
            .I(N__17567));
    SRMux I__3633 (
            .O(N__17604),
            .I(N__17564));
    SRMux I__3632 (
            .O(N__17603),
            .I(N__17561));
    IoInMux I__3631 (
            .O(N__17602),
            .I(N__17556));
    LocalMux I__3630 (
            .O(N__17599),
            .I(N__17553));
    SRMux I__3629 (
            .O(N__17598),
            .I(N__17550));
    Span4Mux_v I__3628 (
            .O(N__17595),
            .I(N__17544));
    LocalMux I__3627 (
            .O(N__17592),
            .I(N__17544));
    SRMux I__3626 (
            .O(N__17591),
            .I(N__17541));
    SRMux I__3625 (
            .O(N__17590),
            .I(N__17537));
    SRMux I__3624 (
            .O(N__17589),
            .I(N__17534));
    LocalMux I__3623 (
            .O(N__17586),
            .I(N__17530));
    SRMux I__3622 (
            .O(N__17585),
            .I(N__17527));
    SRMux I__3621 (
            .O(N__17584),
            .I(N__17524));
    LocalMux I__3620 (
            .O(N__17581),
            .I(N__17519));
    Span4Mux_h I__3619 (
            .O(N__17578),
            .I(N__17510));
    Span4Mux_v I__3618 (
            .O(N__17567),
            .I(N__17510));
    LocalMux I__3617 (
            .O(N__17564),
            .I(N__17510));
    LocalMux I__3616 (
            .O(N__17561),
            .I(N__17510));
    SRMux I__3615 (
            .O(N__17560),
            .I(N__17507));
    SRMux I__3614 (
            .O(N__17559),
            .I(N__17504));
    LocalMux I__3613 (
            .O(N__17556),
            .I(N__17499));
    Span4Mux_v I__3612 (
            .O(N__17553),
            .I(N__17496));
    LocalMux I__3611 (
            .O(N__17550),
            .I(N__17493));
    SRMux I__3610 (
            .O(N__17549),
            .I(N__17489));
    Span4Mux_v I__3609 (
            .O(N__17544),
            .I(N__17484));
    LocalMux I__3608 (
            .O(N__17541),
            .I(N__17484));
    SRMux I__3607 (
            .O(N__17540),
            .I(N__17481));
    LocalMux I__3606 (
            .O(N__17537),
            .I(N__17478));
    LocalMux I__3605 (
            .O(N__17534),
            .I(N__17475));
    SRMux I__3604 (
            .O(N__17533),
            .I(N__17472));
    Span4Mux_h I__3603 (
            .O(N__17530),
            .I(N__17465));
    LocalMux I__3602 (
            .O(N__17527),
            .I(N__17465));
    LocalMux I__3601 (
            .O(N__17524),
            .I(N__17465));
    SRMux I__3600 (
            .O(N__17523),
            .I(N__17462));
    SRMux I__3599 (
            .O(N__17522),
            .I(N__17459));
    Span4Mux_h I__3598 (
            .O(N__17519),
            .I(N__17449));
    Span4Mux_v I__3597 (
            .O(N__17510),
            .I(N__17449));
    LocalMux I__3596 (
            .O(N__17507),
            .I(N__17449));
    LocalMux I__3595 (
            .O(N__17504),
            .I(N__17449));
    SRMux I__3594 (
            .O(N__17503),
            .I(N__17446));
    SRMux I__3593 (
            .O(N__17502),
            .I(N__17443));
    IoSpan4Mux I__3592 (
            .O(N__17499),
            .I(N__17440));
    Span4Mux_v I__3591 (
            .O(N__17496),
            .I(N__17435));
    Span4Mux_v I__3590 (
            .O(N__17493),
            .I(N__17435));
    SRMux I__3589 (
            .O(N__17492),
            .I(N__17431));
    LocalMux I__3588 (
            .O(N__17489),
            .I(N__17428));
    Span4Mux_v I__3587 (
            .O(N__17484),
            .I(N__17423));
    LocalMux I__3586 (
            .O(N__17481),
            .I(N__17423));
    Span4Mux_v I__3585 (
            .O(N__17478),
            .I(N__17416));
    Span4Mux_h I__3584 (
            .O(N__17475),
            .I(N__17416));
    LocalMux I__3583 (
            .O(N__17472),
            .I(N__17416));
    Span4Mux_v I__3582 (
            .O(N__17465),
            .I(N__17409));
    LocalMux I__3581 (
            .O(N__17462),
            .I(N__17409));
    LocalMux I__3580 (
            .O(N__17459),
            .I(N__17409));
    SRMux I__3579 (
            .O(N__17458),
            .I(N__17406));
    Span4Mux_v I__3578 (
            .O(N__17449),
            .I(N__17399));
    LocalMux I__3577 (
            .O(N__17446),
            .I(N__17399));
    LocalMux I__3576 (
            .O(N__17443),
            .I(N__17399));
    Span4Mux_s3_h I__3575 (
            .O(N__17440),
            .I(N__17396));
    Span4Mux_h I__3574 (
            .O(N__17435),
            .I(N__17393));
    InMux I__3573 (
            .O(N__17434),
            .I(N__17390));
    LocalMux I__3572 (
            .O(N__17431),
            .I(N__17387));
    Span4Mux_h I__3571 (
            .O(N__17428),
            .I(N__17384));
    Span4Mux_v I__3570 (
            .O(N__17423),
            .I(N__17379));
    Span4Mux_v I__3569 (
            .O(N__17416),
            .I(N__17379));
    Span4Mux_v I__3568 (
            .O(N__17409),
            .I(N__17372));
    LocalMux I__3567 (
            .O(N__17406),
            .I(N__17372));
    Span4Mux_v I__3566 (
            .O(N__17399),
            .I(N__17372));
    Span4Mux_h I__3565 (
            .O(N__17396),
            .I(N__17369));
    Span4Mux_v I__3564 (
            .O(N__17393),
            .I(N__17364));
    LocalMux I__3563 (
            .O(N__17390),
            .I(N__17364));
    Span12Mux_s11_v I__3562 (
            .O(N__17387),
            .I(N__17361));
    Span4Mux_v I__3561 (
            .O(N__17384),
            .I(N__17354));
    Span4Mux_h I__3560 (
            .O(N__17379),
            .I(N__17354));
    Span4Mux_h I__3559 (
            .O(N__17372),
            .I(N__17354));
    Span4Mux_h I__3558 (
            .O(N__17369),
            .I(N__17349));
    Span4Mux_v I__3557 (
            .O(N__17364),
            .I(N__17349));
    Span12Mux_v I__3556 (
            .O(N__17361),
            .I(N__17343));
    Span4Mux_h I__3555 (
            .O(N__17354),
            .I(N__17340));
    Span4Mux_v I__3554 (
            .O(N__17349),
            .I(N__17337));
    InMux I__3553 (
            .O(N__17348),
            .I(N__17334));
    InMux I__3552 (
            .O(N__17347),
            .I(N__17329));
    InMux I__3551 (
            .O(N__17346),
            .I(N__17329));
    Odrv12 I__3550 (
            .O(N__17343),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3549 (
            .O(N__17340),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3548 (
            .O(N__17337),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3547 (
            .O(N__17334),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3546 (
            .O(N__17329),
            .I(CONSTANT_ONE_NET));
    InMux I__3545 (
            .O(N__17318),
            .I(bfn_15_25_0_));
    InMux I__3544 (
            .O(N__17315),
            .I(N__17312));
    LocalMux I__3543 (
            .O(N__17312),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    CascadeMux I__3542 (
            .O(N__17309),
            .I(N__17306));
    InMux I__3541 (
            .O(N__17306),
            .I(N__17303));
    LocalMux I__3540 (
            .O(N__17303),
            .I(N__17299));
    CascadeMux I__3539 (
            .O(N__17302),
            .I(N__17296));
    Span4Mux_h I__3538 (
            .O(N__17299),
            .I(N__17293));
    InMux I__3537 (
            .O(N__17296),
            .I(N__17290));
    Span4Mux_v I__3536 (
            .O(N__17293),
            .I(N__17287));
    LocalMux I__3535 (
            .O(N__17290),
            .I(N__17284));
    Span4Mux_v I__3534 (
            .O(N__17287),
            .I(N__17281));
    Span4Mux_h I__3533 (
            .O(N__17284),
            .I(N__17278));
    Odrv4 I__3532 (
            .O(N__17281),
            .I(N_13_0));
    Odrv4 I__3531 (
            .O(N__17278),
            .I(N_13_0));
    InMux I__3530 (
            .O(N__17273),
            .I(N__17267));
    InMux I__3529 (
            .O(N__17272),
            .I(N__17267));
    LocalMux I__3528 (
            .O(N__17267),
            .I(M_this_vga_signals_address_5));
    InMux I__3527 (
            .O(N__17264),
            .I(N__17260));
    InMux I__3526 (
            .O(N__17263),
            .I(N__17257));
    LocalMux I__3525 (
            .O(N__17260),
            .I(\this_ppu.un5_sprites_addr_1_c4 ));
    LocalMux I__3524 (
            .O(N__17257),
            .I(\this_ppu.un5_sprites_addr_1_c4 ));
    InMux I__3523 (
            .O(N__17252),
            .I(un1_M_this_data_count_q_cry_3));
    InMux I__3522 (
            .O(N__17249),
            .I(un1_M_this_data_count_q_cry_4));
    InMux I__3521 (
            .O(N__17246),
            .I(un1_M_this_data_count_q_cry_5));
    InMux I__3520 (
            .O(N__17243),
            .I(un1_M_this_data_count_q_cry_6));
    InMux I__3519 (
            .O(N__17240),
            .I(bfn_15_24_0_));
    InMux I__3518 (
            .O(N__17237),
            .I(un1_M_this_data_count_q_cry_8));
    InMux I__3517 (
            .O(N__17234),
            .I(un1_M_this_data_count_q_cry_9));
    InMux I__3516 (
            .O(N__17231),
            .I(un1_M_this_data_count_q_cry_10));
    InMux I__3515 (
            .O(N__17228),
            .I(un1_M_this_data_count_q_cry_11));
    InMux I__3514 (
            .O(N__17225),
            .I(N__17222));
    LocalMux I__3513 (
            .O(N__17222),
            .I(M_this_internal_address_q_3_ns_1_9));
    CascadeMux I__3512 (
            .O(N__17219),
            .I(M_this_internal_address_q_3_ns_1_3_cascade_));
    InMux I__3511 (
            .O(N__17216),
            .I(N__17213));
    LocalMux I__3510 (
            .O(N__17213),
            .I(M_this_internal_address_q_3_ns_1_8));
    InMux I__3509 (
            .O(N__17210),
            .I(un1_M_this_data_count_q_cry_0));
    InMux I__3508 (
            .O(N__17207),
            .I(un1_M_this_data_count_q_cry_1));
    InMux I__3507 (
            .O(N__17204),
            .I(un1_M_this_data_count_q_cry_2));
    InMux I__3506 (
            .O(N__17201),
            .I(N__17195));
    InMux I__3505 (
            .O(N__17200),
            .I(N__17195));
    LocalMux I__3504 (
            .O(N__17195),
            .I(N__17191));
    CascadeMux I__3503 (
            .O(N__17194),
            .I(N__17187));
    Span4Mux_h I__3502 (
            .O(N__17191),
            .I(N__17184));
    InMux I__3501 (
            .O(N__17190),
            .I(N__17179));
    InMux I__3500 (
            .O(N__17187),
            .I(N__17179));
    Odrv4 I__3499 (
            .O(N__17184),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3));
    LocalMux I__3498 (
            .O(N__17179),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3));
    InMux I__3497 (
            .O(N__17174),
            .I(N__17165));
    InMux I__3496 (
            .O(N__17173),
            .I(N__17165));
    InMux I__3495 (
            .O(N__17172),
            .I(N__17160));
    InMux I__3494 (
            .O(N__17171),
            .I(N__17160));
    InMux I__3493 (
            .O(N__17170),
            .I(N__17157));
    LocalMux I__3492 (
            .O(N__17165),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0));
    LocalMux I__3491 (
            .O(N__17160),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0));
    LocalMux I__3490 (
            .O(N__17157),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0));
    InMux I__3489 (
            .O(N__17150),
            .I(N__17133));
    InMux I__3488 (
            .O(N__17149),
            .I(N__17133));
    InMux I__3487 (
            .O(N__17148),
            .I(N__17133));
    InMux I__3486 (
            .O(N__17147),
            .I(N__17128));
    InMux I__3485 (
            .O(N__17146),
            .I(N__17128));
    InMux I__3484 (
            .O(N__17145),
            .I(N__17123));
    InMux I__3483 (
            .O(N__17144),
            .I(N__17123));
    InMux I__3482 (
            .O(N__17143),
            .I(N__17120));
    InMux I__3481 (
            .O(N__17142),
            .I(N__17111));
    InMux I__3480 (
            .O(N__17141),
            .I(N__17111));
    InMux I__3479 (
            .O(N__17140),
            .I(N__17111));
    LocalMux I__3478 (
            .O(N__17133),
            .I(N__17108));
    LocalMux I__3477 (
            .O(N__17128),
            .I(N__17103));
    LocalMux I__3476 (
            .O(N__17123),
            .I(N__17103));
    LocalMux I__3475 (
            .O(N__17120),
            .I(N__17100));
    InMux I__3474 (
            .O(N__17119),
            .I(N__17095));
    InMux I__3473 (
            .O(N__17118),
            .I(N__17095));
    LocalMux I__3472 (
            .O(N__17111),
            .I(N__17092));
    Span4Mux_v I__3471 (
            .O(N__17108),
            .I(N__17087));
    Span4Mux_h I__3470 (
            .O(N__17103),
            .I(N__17087));
    Span12Mux_v I__3469 (
            .O(N__17100),
            .I(N__17083));
    LocalMux I__3468 (
            .O(N__17095),
            .I(N__17080));
    Span4Mux_h I__3467 (
            .O(N__17092),
            .I(N__17077));
    Span4Mux_h I__3466 (
            .O(N__17087),
            .I(N__17074));
    InMux I__3465 (
            .O(N__17086),
            .I(N__17071));
    Span12Mux_h I__3464 (
            .O(N__17083),
            .I(N__17068));
    Odrv12 I__3463 (
            .O(N__17080),
            .I(\this_vga_signals.GZ0Z_210 ));
    Odrv4 I__3462 (
            .O(N__17077),
            .I(\this_vga_signals.GZ0Z_210 ));
    Odrv4 I__3461 (
            .O(N__17074),
            .I(\this_vga_signals.GZ0Z_210 ));
    LocalMux I__3460 (
            .O(N__17071),
            .I(\this_vga_signals.GZ0Z_210 ));
    Odrv12 I__3459 (
            .O(N__17068),
            .I(\this_vga_signals.GZ0Z_210 ));
    SRMux I__3458 (
            .O(N__17057),
            .I(N__17051));
    SRMux I__3457 (
            .O(N__17056),
            .I(N__17048));
    SRMux I__3456 (
            .O(N__17055),
            .I(N__17045));
    SRMux I__3455 (
            .O(N__17054),
            .I(N__17042));
    LocalMux I__3454 (
            .O(N__17051),
            .I(N__17039));
    LocalMux I__3453 (
            .O(N__17048),
            .I(N__17036));
    LocalMux I__3452 (
            .O(N__17045),
            .I(N__17033));
    LocalMux I__3451 (
            .O(N__17042),
            .I(N__17030));
    Span4Mux_v I__3450 (
            .O(N__17039),
            .I(N__17026));
    Span4Mux_h I__3449 (
            .O(N__17036),
            .I(N__17021));
    Span4Mux_v I__3448 (
            .O(N__17033),
            .I(N__17021));
    Span4Mux_v I__3447 (
            .O(N__17030),
            .I(N__17018));
    InMux I__3446 (
            .O(N__17029),
            .I(N__17015));
    Odrv4 I__3445 (
            .O(N__17026),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9 ));
    Odrv4 I__3444 (
            .O(N__17021),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9 ));
    Odrv4 I__3443 (
            .O(N__17018),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9 ));
    LocalMux I__3442 (
            .O(N__17015),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9 ));
    InMux I__3441 (
            .O(N__17006),
            .I(N__17003));
    LocalMux I__3440 (
            .O(N__17003),
            .I(N__16997));
    InMux I__3439 (
            .O(N__17002),
            .I(N__16993));
    InMux I__3438 (
            .O(N__17001),
            .I(N__16989));
    CascadeMux I__3437 (
            .O(N__17000),
            .I(N__16983));
    Span4Mux_v I__3436 (
            .O(N__16997),
            .I(N__16980));
    InMux I__3435 (
            .O(N__16996),
            .I(N__16977));
    LocalMux I__3434 (
            .O(N__16993),
            .I(N__16974));
    InMux I__3433 (
            .O(N__16992),
            .I(N__16971));
    LocalMux I__3432 (
            .O(N__16989),
            .I(N__16968));
    InMux I__3431 (
            .O(N__16988),
            .I(N__16964));
    InMux I__3430 (
            .O(N__16987),
            .I(N__16961));
    InMux I__3429 (
            .O(N__16986),
            .I(N__16956));
    InMux I__3428 (
            .O(N__16983),
            .I(N__16956));
    Span4Mux_h I__3427 (
            .O(N__16980),
            .I(N__16948));
    LocalMux I__3426 (
            .O(N__16977),
            .I(N__16948));
    Span4Mux_v I__3425 (
            .O(N__16974),
            .I(N__16948));
    LocalMux I__3424 (
            .O(N__16971),
            .I(N__16943));
    Span4Mux_v I__3423 (
            .O(N__16968),
            .I(N__16943));
    InMux I__3422 (
            .O(N__16967),
            .I(N__16940));
    LocalMux I__3421 (
            .O(N__16964),
            .I(N__16935));
    LocalMux I__3420 (
            .O(N__16961),
            .I(N__16935));
    LocalMux I__3419 (
            .O(N__16956),
            .I(N__16932));
    InMux I__3418 (
            .O(N__16955),
            .I(N__16929));
    Odrv4 I__3417 (
            .O(N__16948),
            .I(this_vga_signals_M_hcounter_q_3));
    Odrv4 I__3416 (
            .O(N__16943),
            .I(this_vga_signals_M_hcounter_q_3));
    LocalMux I__3415 (
            .O(N__16940),
            .I(this_vga_signals_M_hcounter_q_3));
    Odrv4 I__3414 (
            .O(N__16935),
            .I(this_vga_signals_M_hcounter_q_3));
    Odrv12 I__3413 (
            .O(N__16932),
            .I(this_vga_signals_M_hcounter_q_3));
    LocalMux I__3412 (
            .O(N__16929),
            .I(this_vga_signals_M_hcounter_q_3));
    InMux I__3411 (
            .O(N__16916),
            .I(N__16913));
    LocalMux I__3410 (
            .O(N__16913),
            .I(\this_vga_signals.if_N_9_1 ));
    InMux I__3409 (
            .O(N__16910),
            .I(N__16907));
    LocalMux I__3408 (
            .O(N__16907),
            .I(\this_ppu.sprites_m1_0_xZ0Z1 ));
    CascadeMux I__3407 (
            .O(N__16904),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3_cascade_));
    InMux I__3406 (
            .O(N__16901),
            .I(N__16898));
    LocalMux I__3405 (
            .O(N__16898),
            .I(\this_ppu.sprites_m1_0_xZ0Z0 ));
    InMux I__3404 (
            .O(N__16895),
            .I(N__16892));
    LocalMux I__3403 (
            .O(N__16892),
            .I(M_this_internal_address_q_3_ns_1_2));
    InMux I__3402 (
            .O(N__16889),
            .I(N__16884));
    InMux I__3401 (
            .O(N__16888),
            .I(N__16879));
    InMux I__3400 (
            .O(N__16887),
            .I(N__16879));
    LocalMux I__3399 (
            .O(N__16884),
            .I(\this_pixel_clk.M_counter_qZ0Z_0 ));
    LocalMux I__3398 (
            .O(N__16879),
            .I(\this_pixel_clk.M_counter_qZ0Z_0 ));
    InMux I__3397 (
            .O(N__16874),
            .I(N__16871));
    LocalMux I__3396 (
            .O(N__16871),
            .I(N__16864));
    InMux I__3395 (
            .O(N__16870),
            .I(N__16861));
    CascadeMux I__3394 (
            .O(N__16869),
            .I(N__16857));
    CascadeMux I__3393 (
            .O(N__16868),
            .I(N__16854));
    InMux I__3392 (
            .O(N__16867),
            .I(N__16850));
    Span4Mux_h I__3391 (
            .O(N__16864),
            .I(N__16845));
    LocalMux I__3390 (
            .O(N__16861),
            .I(N__16845));
    InMux I__3389 (
            .O(N__16860),
            .I(N__16842));
    InMux I__3388 (
            .O(N__16857),
            .I(N__16835));
    InMux I__3387 (
            .O(N__16854),
            .I(N__16835));
    InMux I__3386 (
            .O(N__16853),
            .I(N__16835));
    LocalMux I__3385 (
            .O(N__16850),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    Odrv4 I__3384 (
            .O(N__16845),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__3383 (
            .O(N__16842),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    LocalMux I__3382 (
            .O(N__16835),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    CascadeMux I__3381 (
            .O(N__16826),
            .I(if_generate_plus_mult1_un75_sum_axbxc3_cascade_));
    CascadeMux I__3380 (
            .O(N__16823),
            .I(\this_ppu.un5_sprites_addr_1_c2_cascade_ ));
    CascadeMux I__3379 (
            .O(N__16820),
            .I(N__16817));
    InMux I__3378 (
            .O(N__16817),
            .I(N__16812));
    InMux I__3377 (
            .O(N__16816),
            .I(N__16809));
    InMux I__3376 (
            .O(N__16815),
            .I(N__16806));
    LocalMux I__3375 (
            .O(N__16812),
            .I(N__16803));
    LocalMux I__3374 (
            .O(N__16809),
            .I(N__16800));
    LocalMux I__3373 (
            .O(N__16806),
            .I(\this_ppu.N_4_0_1 ));
    Odrv4 I__3372 (
            .O(N__16803),
            .I(\this_ppu.N_4_0_1 ));
    Odrv4 I__3371 (
            .O(N__16800),
            .I(\this_ppu.N_4_0_1 ));
    InMux I__3370 (
            .O(N__16793),
            .I(N__16790));
    LocalMux I__3369 (
            .O(N__16790),
            .I(\this_ppu.sprites_addr_1_i_7_tz_0_9 ));
    InMux I__3368 (
            .O(N__16787),
            .I(N__16784));
    LocalMux I__3367 (
            .O(N__16784),
            .I(N__16781));
    Odrv4 I__3366 (
            .O(N__16781),
            .I(\this_ppu.sprites_addr_1_i_a7Z0Z_9 ));
    InMux I__3365 (
            .O(N__16778),
            .I(N__16775));
    LocalMux I__3364 (
            .O(N__16775),
            .I(N__16770));
    InMux I__3363 (
            .O(N__16774),
            .I(N__16765));
    InMux I__3362 (
            .O(N__16773),
            .I(N__16765));
    Span4Mux_h I__3361 (
            .O(N__16770),
            .I(N__16759));
    LocalMux I__3360 (
            .O(N__16765),
            .I(N__16756));
    InMux I__3359 (
            .O(N__16764),
            .I(N__16753));
    InMux I__3358 (
            .O(N__16763),
            .I(N__16748));
    InMux I__3357 (
            .O(N__16762),
            .I(N__16748));
    Odrv4 I__3356 (
            .O(N__16759),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3));
    Odrv4 I__3355 (
            .O(N__16756),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3));
    LocalMux I__3354 (
            .O(N__16753),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3));
    LocalMux I__3353 (
            .O(N__16748),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3));
    CascadeMux I__3352 (
            .O(N__16739),
            .I(N__16736));
    InMux I__3351 (
            .O(N__16736),
            .I(N__16733));
    LocalMux I__3350 (
            .O(N__16733),
            .I(\this_ppu.un5_sprites_addr1_4 ));
    CascadeMux I__3349 (
            .O(N__16730),
            .I(\this_vga_signals.if_N_8_i_0_cascade_ ));
    InMux I__3348 (
            .O(N__16727),
            .I(N__16722));
    InMux I__3347 (
            .O(N__16726),
            .I(N__16717));
    InMux I__3346 (
            .O(N__16725),
            .I(N__16717));
    LocalMux I__3345 (
            .O(N__16722),
            .I(\this_vga_signals.mult1_un68_sum_axb1_1 ));
    LocalMux I__3344 (
            .O(N__16717),
            .I(\this_vga_signals.mult1_un68_sum_axb1_1 ));
    InMux I__3343 (
            .O(N__16712),
            .I(N__16709));
    LocalMux I__3342 (
            .O(N__16709),
            .I(M_counter_q_RNIFKS8_0));
    CascadeMux I__3341 (
            .O(N__16706),
            .I(M_counter_q_RNIFKS8_0_cascade_));
    InMux I__3340 (
            .O(N__16703),
            .I(N__16691));
    InMux I__3339 (
            .O(N__16702),
            .I(N__16691));
    InMux I__3338 (
            .O(N__16701),
            .I(N__16691));
    InMux I__3337 (
            .O(N__16700),
            .I(N__16691));
    LocalMux I__3336 (
            .O(N__16691),
            .I(this_pixel_clk_M_counter_q_i_1));
    InMux I__3335 (
            .O(N__16688),
            .I(N__16685));
    LocalMux I__3334 (
            .O(N__16685),
            .I(\this_vga_signals.N_455 ));
    CascadeMux I__3333 (
            .O(N__16682),
            .I(N__16679));
    InMux I__3332 (
            .O(N__16679),
            .I(N__16675));
    InMux I__3331 (
            .O(N__16678),
            .I(N__16672));
    LocalMux I__3330 (
            .O(N__16675),
            .I(N__16669));
    LocalMux I__3329 (
            .O(N__16672),
            .I(N__16666));
    Span4Mux_h I__3328 (
            .O(N__16669),
            .I(N__16663));
    Span4Mux_h I__3327 (
            .O(N__16666),
            .I(N__16656));
    Span4Mux_h I__3326 (
            .O(N__16663),
            .I(N__16656));
    InMux I__3325 (
            .O(N__16662),
            .I(N__16651));
    InMux I__3324 (
            .O(N__16661),
            .I(N__16651));
    Odrv4 I__3323 (
            .O(N__16656),
            .I(\this_vga_signals.N_459 ));
    LocalMux I__3322 (
            .O(N__16651),
            .I(\this_vga_signals.N_459 ));
    CascadeMux I__3321 (
            .O(N__16646),
            .I(\this_vga_signals.GZ0Z_210_cascade_ ));
    InMux I__3320 (
            .O(N__16643),
            .I(N__16634));
    InMux I__3319 (
            .O(N__16642),
            .I(N__16631));
    InMux I__3318 (
            .O(N__16641),
            .I(N__16627));
    InMux I__3317 (
            .O(N__16640),
            .I(N__16624));
    InMux I__3316 (
            .O(N__16639),
            .I(N__16621));
    InMux I__3315 (
            .O(N__16638),
            .I(N__16616));
    InMux I__3314 (
            .O(N__16637),
            .I(N__16616));
    LocalMux I__3313 (
            .O(N__16634),
            .I(N__16608));
    LocalMux I__3312 (
            .O(N__16631),
            .I(N__16605));
    InMux I__3311 (
            .O(N__16630),
            .I(N__16602));
    LocalMux I__3310 (
            .O(N__16627),
            .I(N__16599));
    LocalMux I__3309 (
            .O(N__16624),
            .I(N__16592));
    LocalMux I__3308 (
            .O(N__16621),
            .I(N__16592));
    LocalMux I__3307 (
            .O(N__16616),
            .I(N__16592));
    CascadeMux I__3306 (
            .O(N__16615),
            .I(N__16589));
    CascadeMux I__3305 (
            .O(N__16614),
            .I(N__16585));
    InMux I__3304 (
            .O(N__16613),
            .I(N__16582));
    InMux I__3303 (
            .O(N__16612),
            .I(N__16578));
    InMux I__3302 (
            .O(N__16611),
            .I(N__16575));
    Span4Mux_v I__3301 (
            .O(N__16608),
            .I(N__16572));
    Span12Mux_s9_h I__3300 (
            .O(N__16605),
            .I(N__16569));
    LocalMux I__3299 (
            .O(N__16602),
            .I(N__16562));
    Span4Mux_h I__3298 (
            .O(N__16599),
            .I(N__16562));
    Span4Mux_v I__3297 (
            .O(N__16592),
            .I(N__16562));
    InMux I__3296 (
            .O(N__16589),
            .I(N__16555));
    InMux I__3295 (
            .O(N__16588),
            .I(N__16555));
    InMux I__3294 (
            .O(N__16585),
            .I(N__16555));
    LocalMux I__3293 (
            .O(N__16582),
            .I(N__16552));
    InMux I__3292 (
            .O(N__16581),
            .I(N__16549));
    LocalMux I__3291 (
            .O(N__16578),
            .I(N__16544));
    LocalMux I__3290 (
            .O(N__16575),
            .I(N__16544));
    Odrv4 I__3289 (
            .O(N__16572),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv12 I__3288 (
            .O(N__16569),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__3287 (
            .O(N__16562),
            .I(this_vga_signals_M_vcounter_q_9));
    LocalMux I__3286 (
            .O(N__16555),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__3285 (
            .O(N__16552),
            .I(this_vga_signals_M_vcounter_q_9));
    LocalMux I__3284 (
            .O(N__16549),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__3283 (
            .O(N__16544),
            .I(this_vga_signals_M_vcounter_q_9));
    IoInMux I__3282 (
            .O(N__16529),
            .I(N__16526));
    LocalMux I__3281 (
            .O(N__16526),
            .I(N__16523));
    IoSpan4Mux I__3280 (
            .O(N__16523),
            .I(N__16520));
    Span4Mux_s0_h I__3279 (
            .O(N__16520),
            .I(N__16517));
    Sp12to4 I__3278 (
            .O(N__16517),
            .I(N__16514));
    Span12Mux_s8_h I__3277 (
            .O(N__16514),
            .I(N__16511));
    Odrv12 I__3276 (
            .O(N__16511),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIIRV75Z0Z_9 ));
    InMux I__3275 (
            .O(N__16508),
            .I(N__16505));
    LocalMux I__3274 (
            .O(N__16505),
            .I(N__16502));
    Odrv4 I__3273 (
            .O(N__16502),
            .I(\this_ppu.sprites_addr_1_i_2_1Z0Z_9 ));
    CascadeMux I__3272 (
            .O(N__16499),
            .I(\this_ppu.sprites_addr_1_i_0_0Z0Z_9_cascade_ ));
    InMux I__3271 (
            .O(N__16496),
            .I(N__16493));
    LocalMux I__3270 (
            .O(N__16493),
            .I(N__16490));
    Span4Mux_h I__3269 (
            .O(N__16490),
            .I(N__16487));
    Odrv4 I__3268 (
            .O(N__16487),
            .I(\this_ppu.sprites_addr_1_i_a0_2Z0Z_9 ));
    CascadeMux I__3267 (
            .O(N__16484),
            .I(\this_ppu.sprites_addr_1_i_0_2Z0Z_9_cascade_ ));
    CascadeMux I__3266 (
            .O(N__16481),
            .I(N__16478));
    CascadeBuf I__3265 (
            .O(N__16478),
            .I(N__16475));
    CascadeMux I__3264 (
            .O(N__16475),
            .I(N__16472));
    CascadeBuf I__3263 (
            .O(N__16472),
            .I(N__16469));
    CascadeMux I__3262 (
            .O(N__16469),
            .I(N__16466));
    CascadeBuf I__3261 (
            .O(N__16466),
            .I(N__16463));
    CascadeMux I__3260 (
            .O(N__16463),
            .I(N__16460));
    CascadeBuf I__3259 (
            .O(N__16460),
            .I(N__16457));
    CascadeMux I__3258 (
            .O(N__16457),
            .I(N__16454));
    CascadeBuf I__3257 (
            .O(N__16454),
            .I(N__16451));
    CascadeMux I__3256 (
            .O(N__16451),
            .I(N__16448));
    CascadeBuf I__3255 (
            .O(N__16448),
            .I(N__16445));
    CascadeMux I__3254 (
            .O(N__16445),
            .I(N__16442));
    CascadeBuf I__3253 (
            .O(N__16442),
            .I(N__16439));
    CascadeMux I__3252 (
            .O(N__16439),
            .I(N__16436));
    CascadeBuf I__3251 (
            .O(N__16436),
            .I(N__16433));
    CascadeMux I__3250 (
            .O(N__16433),
            .I(N__16430));
    CascadeBuf I__3249 (
            .O(N__16430),
            .I(N__16427));
    CascadeMux I__3248 (
            .O(N__16427),
            .I(N__16424));
    CascadeBuf I__3247 (
            .O(N__16424),
            .I(N__16421));
    CascadeMux I__3246 (
            .O(N__16421),
            .I(N__16418));
    CascadeBuf I__3245 (
            .O(N__16418),
            .I(N__16415));
    CascadeMux I__3244 (
            .O(N__16415),
            .I(N__16412));
    CascadeBuf I__3243 (
            .O(N__16412),
            .I(N__16409));
    CascadeMux I__3242 (
            .O(N__16409),
            .I(N__16406));
    CascadeBuf I__3241 (
            .O(N__16406),
            .I(N__16403));
    CascadeMux I__3240 (
            .O(N__16403),
            .I(N__16400));
    CascadeBuf I__3239 (
            .O(N__16400),
            .I(N__16397));
    CascadeMux I__3238 (
            .O(N__16397),
            .I(N__16394));
    CascadeBuf I__3237 (
            .O(N__16394),
            .I(N__16391));
    CascadeMux I__3236 (
            .O(N__16391),
            .I(N__16388));
    InMux I__3235 (
            .O(N__16388),
            .I(N__16385));
    LocalMux I__3234 (
            .O(N__16385),
            .I(N__16382));
    Span12Mux_h I__3233 (
            .O(N__16382),
            .I(N__16379));
    Span12Mux_v I__3232 (
            .O(N__16379),
            .I(N__16376));
    Odrv12 I__3231 (
            .O(N__16376),
            .I(N_138_0));
    InMux I__3230 (
            .O(N__16373),
            .I(N__16370));
    LocalMux I__3229 (
            .O(N__16370),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_0_1 ));
    InMux I__3228 (
            .O(N__16367),
            .I(N__16364));
    LocalMux I__3227 (
            .O(N__16364),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_x0 ));
    InMux I__3226 (
            .O(N__16361),
            .I(N__16358));
    LocalMux I__3225 (
            .O(N__16358),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_x1 ));
    InMux I__3224 (
            .O(N__16355),
            .I(N__16352));
    LocalMux I__3223 (
            .O(N__16352),
            .I(\this_vga_signals.mult1_un75_sum_ac0_1 ));
    CascadeMux I__3222 (
            .O(N__16349),
            .I(if_generate_plus_mult1_un68_sum_axbxc3_ns_cascade_));
    CascadeMux I__3221 (
            .O(N__16346),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_cascade_));
    InMux I__3220 (
            .O(N__16343),
            .I(N__16339));
    CascadeMux I__3219 (
            .O(N__16342),
            .I(N__16335));
    LocalMux I__3218 (
            .O(N__16339),
            .I(N__16332));
    InMux I__3217 (
            .O(N__16338),
            .I(N__16329));
    InMux I__3216 (
            .O(N__16335),
            .I(N__16326));
    Span4Mux_h I__3215 (
            .O(N__16332),
            .I(N__16323));
    LocalMux I__3214 (
            .O(N__16329),
            .I(N__16320));
    LocalMux I__3213 (
            .O(N__16326),
            .I(N__16311));
    Span4Mux_v I__3212 (
            .O(N__16323),
            .I(N__16304));
    Span4Mux_h I__3211 (
            .O(N__16320),
            .I(N__16304));
    InMux I__3210 (
            .O(N__16319),
            .I(N__16301));
    InMux I__3209 (
            .O(N__16318),
            .I(N__16292));
    InMux I__3208 (
            .O(N__16317),
            .I(N__16292));
    InMux I__3207 (
            .O(N__16316),
            .I(N__16292));
    InMux I__3206 (
            .O(N__16315),
            .I(N__16292));
    CascadeMux I__3205 (
            .O(N__16314),
            .I(N__16287));
    Span4Mux_v I__3204 (
            .O(N__16311),
            .I(N__16281));
    InMux I__3203 (
            .O(N__16310),
            .I(N__16278));
    InMux I__3202 (
            .O(N__16309),
            .I(N__16275));
    Span4Mux_h I__3201 (
            .O(N__16304),
            .I(N__16268));
    LocalMux I__3200 (
            .O(N__16301),
            .I(N__16268));
    LocalMux I__3199 (
            .O(N__16292),
            .I(N__16268));
    InMux I__3198 (
            .O(N__16291),
            .I(N__16257));
    InMux I__3197 (
            .O(N__16290),
            .I(N__16257));
    InMux I__3196 (
            .O(N__16287),
            .I(N__16257));
    InMux I__3195 (
            .O(N__16286),
            .I(N__16257));
    InMux I__3194 (
            .O(N__16285),
            .I(N__16257));
    InMux I__3193 (
            .O(N__16284),
            .I(N__16254));
    Odrv4 I__3192 (
            .O(N__16281),
            .I(this_vga_signals_M_hcounter_q_5));
    LocalMux I__3191 (
            .O(N__16278),
            .I(this_vga_signals_M_hcounter_q_5));
    LocalMux I__3190 (
            .O(N__16275),
            .I(this_vga_signals_M_hcounter_q_5));
    Odrv4 I__3189 (
            .O(N__16268),
            .I(this_vga_signals_M_hcounter_q_5));
    LocalMux I__3188 (
            .O(N__16257),
            .I(this_vga_signals_M_hcounter_q_5));
    LocalMux I__3187 (
            .O(N__16254),
            .I(this_vga_signals_M_hcounter_q_5));
    CascadeMux I__3186 (
            .O(N__16241),
            .I(N__16237));
    CascadeMux I__3185 (
            .O(N__16240),
            .I(N__16234));
    InMux I__3184 (
            .O(N__16237),
            .I(N__16230));
    InMux I__3183 (
            .O(N__16234),
            .I(N__16225));
    InMux I__3182 (
            .O(N__16233),
            .I(N__16225));
    LocalMux I__3181 (
            .O(N__16230),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0 ));
    LocalMux I__3180 (
            .O(N__16225),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0 ));
    InMux I__3179 (
            .O(N__16220),
            .I(N__16217));
    LocalMux I__3178 (
            .O(N__16217),
            .I(N__16211));
    InMux I__3177 (
            .O(N__16216),
            .I(N__16208));
    InMux I__3176 (
            .O(N__16215),
            .I(N__16199));
    InMux I__3175 (
            .O(N__16214),
            .I(N__16194));
    Span4Mux_h I__3174 (
            .O(N__16211),
            .I(N__16191));
    LocalMux I__3173 (
            .O(N__16208),
            .I(N__16188));
    InMux I__3172 (
            .O(N__16207),
            .I(N__16185));
    InMux I__3171 (
            .O(N__16206),
            .I(N__16182));
    InMux I__3170 (
            .O(N__16205),
            .I(N__16179));
    InMux I__3169 (
            .O(N__16204),
            .I(N__16172));
    InMux I__3168 (
            .O(N__16203),
            .I(N__16172));
    InMux I__3167 (
            .O(N__16202),
            .I(N__16172));
    LocalMux I__3166 (
            .O(N__16199),
            .I(N__16164));
    InMux I__3165 (
            .O(N__16198),
            .I(N__16161));
    InMux I__3164 (
            .O(N__16197),
            .I(N__16158));
    LocalMux I__3163 (
            .O(N__16194),
            .I(N__16155));
    Span4Mux_h I__3162 (
            .O(N__16191),
            .I(N__16148));
    Span4Mux_h I__3161 (
            .O(N__16188),
            .I(N__16148));
    LocalMux I__3160 (
            .O(N__16185),
            .I(N__16148));
    LocalMux I__3159 (
            .O(N__16182),
            .I(N__16141));
    LocalMux I__3158 (
            .O(N__16179),
            .I(N__16141));
    LocalMux I__3157 (
            .O(N__16172),
            .I(N__16141));
    InMux I__3156 (
            .O(N__16171),
            .I(N__16130));
    InMux I__3155 (
            .O(N__16170),
            .I(N__16130));
    InMux I__3154 (
            .O(N__16169),
            .I(N__16130));
    InMux I__3153 (
            .O(N__16168),
            .I(N__16130));
    InMux I__3152 (
            .O(N__16167),
            .I(N__16130));
    Odrv4 I__3151 (
            .O(N__16164),
            .I(this_vga_signals_M_hcounter_q_4));
    LocalMux I__3150 (
            .O(N__16161),
            .I(this_vga_signals_M_hcounter_q_4));
    LocalMux I__3149 (
            .O(N__16158),
            .I(this_vga_signals_M_hcounter_q_4));
    Odrv12 I__3148 (
            .O(N__16155),
            .I(this_vga_signals_M_hcounter_q_4));
    Odrv4 I__3147 (
            .O(N__16148),
            .I(this_vga_signals_M_hcounter_q_4));
    Odrv4 I__3146 (
            .O(N__16141),
            .I(this_vga_signals_M_hcounter_q_4));
    LocalMux I__3145 (
            .O(N__16130),
            .I(this_vga_signals_M_hcounter_q_4));
    InMux I__3144 (
            .O(N__16115),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_2 ));
    InMux I__3143 (
            .O(N__16112),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_3 ));
    InMux I__3142 (
            .O(N__16109),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_4 ));
    InMux I__3141 (
            .O(N__16106),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_5 ));
    InMux I__3140 (
            .O(N__16103),
            .I(N__16097));
    CascadeMux I__3139 (
            .O(N__16102),
            .I(N__16094));
    InMux I__3138 (
            .O(N__16101),
            .I(N__16089));
    InMux I__3137 (
            .O(N__16100),
            .I(N__16086));
    LocalMux I__3136 (
            .O(N__16097),
            .I(N__16082));
    InMux I__3135 (
            .O(N__16094),
            .I(N__16077));
    InMux I__3134 (
            .O(N__16093),
            .I(N__16077));
    InMux I__3133 (
            .O(N__16092),
            .I(N__16074));
    LocalMux I__3132 (
            .O(N__16089),
            .I(N__16069));
    LocalMux I__3131 (
            .O(N__16086),
            .I(N__16069));
    InMux I__3130 (
            .O(N__16085),
            .I(N__16066));
    Span4Mux_v I__3129 (
            .O(N__16082),
            .I(N__16057));
    LocalMux I__3128 (
            .O(N__16077),
            .I(N__16057));
    LocalMux I__3127 (
            .O(N__16074),
            .I(N__16053));
    Span4Mux_v I__3126 (
            .O(N__16069),
            .I(N__16048));
    LocalMux I__3125 (
            .O(N__16066),
            .I(N__16048));
    InMux I__3124 (
            .O(N__16065),
            .I(N__16045));
    CascadeMux I__3123 (
            .O(N__16064),
            .I(N__16042));
    CascadeMux I__3122 (
            .O(N__16063),
            .I(N__16039));
    InMux I__3121 (
            .O(N__16062),
            .I(N__16036));
    Span4Mux_h I__3120 (
            .O(N__16057),
            .I(N__16033));
    InMux I__3119 (
            .O(N__16056),
            .I(N__16030));
    Span4Mux_v I__3118 (
            .O(N__16053),
            .I(N__16023));
    Span4Mux_h I__3117 (
            .O(N__16048),
            .I(N__16023));
    LocalMux I__3116 (
            .O(N__16045),
            .I(N__16023));
    InMux I__3115 (
            .O(N__16042),
            .I(N__16018));
    InMux I__3114 (
            .O(N__16039),
            .I(N__16018));
    LocalMux I__3113 (
            .O(N__16036),
            .I(this_vga_signals_M_hcounter_q_7));
    Odrv4 I__3112 (
            .O(N__16033),
            .I(this_vga_signals_M_hcounter_q_7));
    LocalMux I__3111 (
            .O(N__16030),
            .I(this_vga_signals_M_hcounter_q_7));
    Odrv4 I__3110 (
            .O(N__16023),
            .I(this_vga_signals_M_hcounter_q_7));
    LocalMux I__3109 (
            .O(N__16018),
            .I(this_vga_signals_M_hcounter_q_7));
    InMux I__3108 (
            .O(N__16007),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_6 ));
    CascadeMux I__3107 (
            .O(N__16004),
            .I(N__15999));
    CascadeMux I__3106 (
            .O(N__16003),
            .I(N__15996));
    InMux I__3105 (
            .O(N__16002),
            .I(N__15993));
    InMux I__3104 (
            .O(N__15999),
            .I(N__15988));
    InMux I__3103 (
            .O(N__15996),
            .I(N__15985));
    LocalMux I__3102 (
            .O(N__15993),
            .I(N__15980));
    InMux I__3101 (
            .O(N__15992),
            .I(N__15977));
    InMux I__3100 (
            .O(N__15991),
            .I(N__15973));
    LocalMux I__3099 (
            .O(N__15988),
            .I(N__15968));
    LocalMux I__3098 (
            .O(N__15985),
            .I(N__15968));
    InMux I__3097 (
            .O(N__15984),
            .I(N__15965));
    CascadeMux I__3096 (
            .O(N__15983),
            .I(N__15962));
    Span4Mux_v I__3095 (
            .O(N__15980),
            .I(N__15954));
    LocalMux I__3094 (
            .O(N__15977),
            .I(N__15954));
    InMux I__3093 (
            .O(N__15976),
            .I(N__15951));
    LocalMux I__3092 (
            .O(N__15973),
            .I(N__15948));
    Span4Mux_v I__3091 (
            .O(N__15968),
            .I(N__15943));
    LocalMux I__3090 (
            .O(N__15965),
            .I(N__15943));
    InMux I__3089 (
            .O(N__15962),
            .I(N__15940));
    InMux I__3088 (
            .O(N__15961),
            .I(N__15935));
    InMux I__3087 (
            .O(N__15960),
            .I(N__15932));
    InMux I__3086 (
            .O(N__15959),
            .I(N__15929));
    Span4Mux_h I__3085 (
            .O(N__15954),
            .I(N__15924));
    LocalMux I__3084 (
            .O(N__15951),
            .I(N__15924));
    Span4Mux_v I__3083 (
            .O(N__15948),
            .I(N__15917));
    Span4Mux_h I__3082 (
            .O(N__15943),
            .I(N__15917));
    LocalMux I__3081 (
            .O(N__15940),
            .I(N__15917));
    InMux I__3080 (
            .O(N__15939),
            .I(N__15914));
    InMux I__3079 (
            .O(N__15938),
            .I(N__15911));
    LocalMux I__3078 (
            .O(N__15935),
            .I(this_vga_signals_M_hcounter_q_8));
    LocalMux I__3077 (
            .O(N__15932),
            .I(this_vga_signals_M_hcounter_q_8));
    LocalMux I__3076 (
            .O(N__15929),
            .I(this_vga_signals_M_hcounter_q_8));
    Odrv4 I__3075 (
            .O(N__15924),
            .I(this_vga_signals_M_hcounter_q_8));
    Odrv4 I__3074 (
            .O(N__15917),
            .I(this_vga_signals_M_hcounter_q_8));
    LocalMux I__3073 (
            .O(N__15914),
            .I(this_vga_signals_M_hcounter_q_8));
    LocalMux I__3072 (
            .O(N__15911),
            .I(this_vga_signals_M_hcounter_q_8));
    InMux I__3071 (
            .O(N__15896),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_7 ));
    InMux I__3070 (
            .O(N__15893),
            .I(bfn_14_18_0_));
    InMux I__3069 (
            .O(N__15890),
            .I(N__15885));
    InMux I__3068 (
            .O(N__15889),
            .I(N__15882));
    InMux I__3067 (
            .O(N__15888),
            .I(N__15879));
    LocalMux I__3066 (
            .O(N__15885),
            .I(N__15870));
    LocalMux I__3065 (
            .O(N__15882),
            .I(N__15870));
    LocalMux I__3064 (
            .O(N__15879),
            .I(N__15867));
    InMux I__3063 (
            .O(N__15878),
            .I(N__15864));
    InMux I__3062 (
            .O(N__15877),
            .I(N__15860));
    InMux I__3061 (
            .O(N__15876),
            .I(N__15857));
    InMux I__3060 (
            .O(N__15875),
            .I(N__15854));
    Span4Mux_v I__3059 (
            .O(N__15870),
            .I(N__15847));
    Span4Mux_v I__3058 (
            .O(N__15867),
            .I(N__15847));
    LocalMux I__3057 (
            .O(N__15864),
            .I(N__15847));
    InMux I__3056 (
            .O(N__15863),
            .I(N__15841));
    LocalMux I__3055 (
            .O(N__15860),
            .I(N__15838));
    LocalMux I__3054 (
            .O(N__15857),
            .I(N__15833));
    LocalMux I__3053 (
            .O(N__15854),
            .I(N__15833));
    Span4Mux_h I__3052 (
            .O(N__15847),
            .I(N__15830));
    InMux I__3051 (
            .O(N__15846),
            .I(N__15827));
    InMux I__3050 (
            .O(N__15845),
            .I(N__15824));
    InMux I__3049 (
            .O(N__15844),
            .I(N__15821));
    LocalMux I__3048 (
            .O(N__15841),
            .I(this_vga_signals_M_hcounter_q_9));
    Odrv4 I__3047 (
            .O(N__15838),
            .I(this_vga_signals_M_hcounter_q_9));
    Odrv4 I__3046 (
            .O(N__15833),
            .I(this_vga_signals_M_hcounter_q_9));
    Odrv4 I__3045 (
            .O(N__15830),
            .I(this_vga_signals_M_hcounter_q_9));
    LocalMux I__3044 (
            .O(N__15827),
            .I(this_vga_signals_M_hcounter_q_9));
    LocalMux I__3043 (
            .O(N__15824),
            .I(this_vga_signals_M_hcounter_q_9));
    LocalMux I__3042 (
            .O(N__15821),
            .I(this_vga_signals_M_hcounter_q_9));
    InMux I__3041 (
            .O(N__15806),
            .I(N__15802));
    InMux I__3040 (
            .O(N__15805),
            .I(N__15799));
    LocalMux I__3039 (
            .O(N__15802),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0 ));
    LocalMux I__3038 (
            .O(N__15799),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0 ));
    InMux I__3037 (
            .O(N__15794),
            .I(N__15785));
    InMux I__3036 (
            .O(N__15793),
            .I(N__15785));
    InMux I__3035 (
            .O(N__15792),
            .I(N__15782));
    CascadeMux I__3034 (
            .O(N__15791),
            .I(N__15778));
    InMux I__3033 (
            .O(N__15790),
            .I(N__15775));
    LocalMux I__3032 (
            .O(N__15785),
            .I(N__15769));
    LocalMux I__3031 (
            .O(N__15782),
            .I(N__15769));
    InMux I__3030 (
            .O(N__15781),
            .I(N__15760));
    InMux I__3029 (
            .O(N__15778),
            .I(N__15760));
    LocalMux I__3028 (
            .O(N__15775),
            .I(N__15757));
    InMux I__3027 (
            .O(N__15774),
            .I(N__15754));
    Span4Mux_v I__3026 (
            .O(N__15769),
            .I(N__15751));
    InMux I__3025 (
            .O(N__15768),
            .I(N__15748));
    CascadeMux I__3024 (
            .O(N__15767),
            .I(N__15745));
    CascadeMux I__3023 (
            .O(N__15766),
            .I(N__15742));
    InMux I__3022 (
            .O(N__15765),
            .I(N__15739));
    LocalMux I__3021 (
            .O(N__15760),
            .I(N__15736));
    Span4Mux_v I__3020 (
            .O(N__15757),
            .I(N__15731));
    LocalMux I__3019 (
            .O(N__15754),
            .I(N__15731));
    Span4Mux_h I__3018 (
            .O(N__15751),
            .I(N__15726));
    LocalMux I__3017 (
            .O(N__15748),
            .I(N__15726));
    InMux I__3016 (
            .O(N__15745),
            .I(N__15723));
    InMux I__3015 (
            .O(N__15742),
            .I(N__15720));
    LocalMux I__3014 (
            .O(N__15739),
            .I(this_vga_signals_M_hcounter_q_6));
    Odrv4 I__3013 (
            .O(N__15736),
            .I(this_vga_signals_M_hcounter_q_6));
    Odrv4 I__3012 (
            .O(N__15731),
            .I(this_vga_signals_M_hcounter_q_6));
    Odrv4 I__3011 (
            .O(N__15726),
            .I(this_vga_signals_M_hcounter_q_6));
    LocalMux I__3010 (
            .O(N__15723),
            .I(this_vga_signals_M_hcounter_q_6));
    LocalMux I__3009 (
            .O(N__15720),
            .I(this_vga_signals_M_hcounter_q_6));
    CEMux I__3008 (
            .O(N__15707),
            .I(N__15703));
    CEMux I__3007 (
            .O(N__15706),
            .I(N__15700));
    LocalMux I__3006 (
            .O(N__15703),
            .I(N__15697));
    LocalMux I__3005 (
            .O(N__15700),
            .I(N__15694));
    Span4Mux_h I__3004 (
            .O(N__15697),
            .I(N__15691));
    Odrv4 I__3003 (
            .O(N__15694),
            .I(\this_vga_signals.N_517_0 ));
    Odrv4 I__3002 (
            .O(N__15691),
            .I(\this_vga_signals.N_517_0 ));
    InMux I__3001 (
            .O(N__15686),
            .I(N__15682));
    InMux I__3000 (
            .O(N__15685),
            .I(N__15679));
    LocalMux I__2999 (
            .O(N__15682),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1 ));
    LocalMux I__2998 (
            .O(N__15679),
            .I(\this_vga_signals.mult1_un61_sum_axbxc1 ));
    InMux I__2997 (
            .O(N__15674),
            .I(N__15671));
    LocalMux I__2996 (
            .O(N__15671),
            .I(N__15668));
    Odrv12 I__2995 (
            .O(N__15668),
            .I(\this_vga_signals.N_3 ));
    CascadeMux I__2994 (
            .O(N__15665),
            .I(N__15662));
    InMux I__2993 (
            .O(N__15662),
            .I(N__15658));
    CascadeMux I__2992 (
            .O(N__15661),
            .I(N__15654));
    LocalMux I__2991 (
            .O(N__15658),
            .I(N__15651));
    InMux I__2990 (
            .O(N__15657),
            .I(N__15646));
    InMux I__2989 (
            .O(N__15654),
            .I(N__15646));
    Span4Mux_h I__2988 (
            .O(N__15651),
            .I(N__15643));
    LocalMux I__2987 (
            .O(N__15646),
            .I(N__15640));
    Sp12to4 I__2986 (
            .O(N__15643),
            .I(N__15636));
    Span4Mux_h I__2985 (
            .O(N__15640),
            .I(N__15633));
    InMux I__2984 (
            .O(N__15639),
            .I(N__15630));
    Odrv12 I__2983 (
            .O(N__15636),
            .I(\this_vga_signals.mult1_un68_sum_s_3 ));
    Odrv4 I__2982 (
            .O(N__15633),
            .I(\this_vga_signals.mult1_un68_sum_s_3 ));
    LocalMux I__2981 (
            .O(N__15630),
            .I(\this_vga_signals.mult1_un68_sum_s_3 ));
    ClkMux I__2980 (
            .O(N__15623),
            .I(N__15617));
    ClkMux I__2979 (
            .O(N__15622),
            .I(N__15614));
    ClkMux I__2978 (
            .O(N__15621),
            .I(N__15610));
    ClkMux I__2977 (
            .O(N__15620),
            .I(N__15606));
    LocalMux I__2976 (
            .O(N__15617),
            .I(N__15601));
    LocalMux I__2975 (
            .O(N__15614),
            .I(N__15601));
    ClkMux I__2974 (
            .O(N__15613),
            .I(N__15598));
    LocalMux I__2973 (
            .O(N__15610),
            .I(N__15595));
    ClkMux I__2972 (
            .O(N__15609),
            .I(N__15592));
    LocalMux I__2971 (
            .O(N__15606),
            .I(N__15589));
    IoSpan4Mux I__2970 (
            .O(N__15601),
            .I(N__15586));
    LocalMux I__2969 (
            .O(N__15598),
            .I(N__15583));
    Span4Mux_s2_h I__2968 (
            .O(N__15595),
            .I(N__15580));
    LocalMux I__2967 (
            .O(N__15592),
            .I(N__15577));
    Span4Mux_s2_h I__2966 (
            .O(N__15589),
            .I(N__15574));
    IoSpan4Mux I__2965 (
            .O(N__15586),
            .I(N__15569));
    IoSpan4Mux I__2964 (
            .O(N__15583),
            .I(N__15569));
    Span4Mux_v I__2963 (
            .O(N__15580),
            .I(N__15566));
    Span4Mux_s2_h I__2962 (
            .O(N__15577),
            .I(N__15563));
    Sp12to4 I__2961 (
            .O(N__15574),
            .I(N__15560));
    Span4Mux_s1_h I__2960 (
            .O(N__15569),
            .I(N__15557));
    Sp12to4 I__2959 (
            .O(N__15566),
            .I(N__15552));
    Sp12to4 I__2958 (
            .O(N__15563),
            .I(N__15552));
    Span12Mux_v I__2957 (
            .O(N__15560),
            .I(N__15545));
    Sp12to4 I__2956 (
            .O(N__15557),
            .I(N__15545));
    Span12Mux_v I__2955 (
            .O(N__15552),
            .I(N__15545));
    Odrv12 I__2954 (
            .O(N__15545),
            .I(M_this_vga_signals_pixel_clk_0));
    InMux I__2953 (
            .O(N__15542),
            .I(N__15539));
    LocalMux I__2952 (
            .O(N__15539),
            .I(N__15534));
    InMux I__2951 (
            .O(N__15538),
            .I(N__15529));
    InMux I__2950 (
            .O(N__15537),
            .I(N__15529));
    Odrv12 I__2949 (
            .O(N__15534),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    LocalMux I__2948 (
            .O(N__15529),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    CEMux I__2947 (
            .O(N__15524),
            .I(N__15503));
    CEMux I__2946 (
            .O(N__15523),
            .I(N__15503));
    CEMux I__2945 (
            .O(N__15522),
            .I(N__15503));
    CEMux I__2944 (
            .O(N__15521),
            .I(N__15503));
    CEMux I__2943 (
            .O(N__15520),
            .I(N__15503));
    CEMux I__2942 (
            .O(N__15519),
            .I(N__15503));
    CEMux I__2941 (
            .O(N__15518),
            .I(N__15503));
    GlobalMux I__2940 (
            .O(N__15503),
            .I(N__15500));
    gio2CtrlBuf I__2939 (
            .O(N__15500),
            .I(\this_vga_signals.N_517_1_g ));
    InMux I__2938 (
            .O(N__15497),
            .I(N__15494));
    LocalMux I__2937 (
            .O(N__15494),
            .I(N__15483));
    SRMux I__2936 (
            .O(N__15493),
            .I(N__15464));
    SRMux I__2935 (
            .O(N__15492),
            .I(N__15464));
    SRMux I__2934 (
            .O(N__15491),
            .I(N__15464));
    SRMux I__2933 (
            .O(N__15490),
            .I(N__15464));
    SRMux I__2932 (
            .O(N__15489),
            .I(N__15464));
    SRMux I__2931 (
            .O(N__15488),
            .I(N__15464));
    SRMux I__2930 (
            .O(N__15487),
            .I(N__15464));
    SRMux I__2929 (
            .O(N__15486),
            .I(N__15464));
    Glb2LocalMux I__2928 (
            .O(N__15483),
            .I(N__15464));
    GlobalMux I__2927 (
            .O(N__15464),
            .I(N__15461));
    gio2CtrlBuf I__2926 (
            .O(N__15461),
            .I(\this_vga_signals.N_684_g ));
    InMux I__2925 (
            .O(N__15458),
            .I(N__15455));
    LocalMux I__2924 (
            .O(N__15455),
            .I(\this_vga_signals.N_272_0 ));
    CascadeMux I__2923 (
            .O(N__15452),
            .I(N__15443));
    CascadeMux I__2922 (
            .O(N__15451),
            .I(N__15437));
    CascadeMux I__2921 (
            .O(N__15450),
            .I(N__15434));
    CascadeMux I__2920 (
            .O(N__15449),
            .I(N__15419));
    CascadeMux I__2919 (
            .O(N__15448),
            .I(N__15416));
    CascadeMux I__2918 (
            .O(N__15447),
            .I(N__15411));
    InMux I__2917 (
            .O(N__15446),
            .I(N__15408));
    InMux I__2916 (
            .O(N__15443),
            .I(N__15403));
    InMux I__2915 (
            .O(N__15442),
            .I(N__15403));
    CascadeMux I__2914 (
            .O(N__15441),
            .I(N__15399));
    CascadeMux I__2913 (
            .O(N__15440),
            .I(N__15394));
    InMux I__2912 (
            .O(N__15437),
            .I(N__15389));
    InMux I__2911 (
            .O(N__15434),
            .I(N__15389));
    InMux I__2910 (
            .O(N__15433),
            .I(N__15384));
    InMux I__2909 (
            .O(N__15432),
            .I(N__15384));
    InMux I__2908 (
            .O(N__15431),
            .I(N__15381));
    InMux I__2907 (
            .O(N__15430),
            .I(N__15376));
    InMux I__2906 (
            .O(N__15429),
            .I(N__15376));
    InMux I__2905 (
            .O(N__15428),
            .I(N__15373));
    CascadeMux I__2904 (
            .O(N__15427),
            .I(N__15370));
    CascadeMux I__2903 (
            .O(N__15426),
            .I(N__15366));
    CascadeMux I__2902 (
            .O(N__15425),
            .I(N__15363));
    CascadeMux I__2901 (
            .O(N__15424),
            .I(N__15359));
    InMux I__2900 (
            .O(N__15423),
            .I(N__15355));
    InMux I__2899 (
            .O(N__15422),
            .I(N__15352));
    InMux I__2898 (
            .O(N__15419),
            .I(N__15349));
    InMux I__2897 (
            .O(N__15416),
            .I(N__15340));
    InMux I__2896 (
            .O(N__15415),
            .I(N__15340));
    InMux I__2895 (
            .O(N__15414),
            .I(N__15340));
    InMux I__2894 (
            .O(N__15411),
            .I(N__15340));
    LocalMux I__2893 (
            .O(N__15408),
            .I(N__15334));
    LocalMux I__2892 (
            .O(N__15403),
            .I(N__15334));
    InMux I__2891 (
            .O(N__15402),
            .I(N__15329));
    InMux I__2890 (
            .O(N__15399),
            .I(N__15329));
    InMux I__2889 (
            .O(N__15398),
            .I(N__15326));
    InMux I__2888 (
            .O(N__15397),
            .I(N__15323));
    InMux I__2887 (
            .O(N__15394),
            .I(N__15320));
    LocalMux I__2886 (
            .O(N__15389),
            .I(N__15315));
    LocalMux I__2885 (
            .O(N__15384),
            .I(N__15315));
    LocalMux I__2884 (
            .O(N__15381),
            .I(N__15308));
    LocalMux I__2883 (
            .O(N__15376),
            .I(N__15308));
    LocalMux I__2882 (
            .O(N__15373),
            .I(N__15308));
    InMux I__2881 (
            .O(N__15370),
            .I(N__15301));
    InMux I__2880 (
            .O(N__15369),
            .I(N__15301));
    InMux I__2879 (
            .O(N__15366),
            .I(N__15301));
    InMux I__2878 (
            .O(N__15363),
            .I(N__15296));
    InMux I__2877 (
            .O(N__15362),
            .I(N__15296));
    InMux I__2876 (
            .O(N__15359),
            .I(N__15293));
    InMux I__2875 (
            .O(N__15358),
            .I(N__15290));
    LocalMux I__2874 (
            .O(N__15355),
            .I(N__15285));
    LocalMux I__2873 (
            .O(N__15352),
            .I(N__15285));
    LocalMux I__2872 (
            .O(N__15349),
            .I(N__15280));
    LocalMux I__2871 (
            .O(N__15340),
            .I(N__15280));
    InMux I__2870 (
            .O(N__15339),
            .I(N__15277));
    Span4Mux_h I__2869 (
            .O(N__15334),
            .I(N__15272));
    LocalMux I__2868 (
            .O(N__15329),
            .I(N__15272));
    LocalMux I__2867 (
            .O(N__15326),
            .I(N__15265));
    LocalMux I__2866 (
            .O(N__15323),
            .I(N__15265));
    LocalMux I__2865 (
            .O(N__15320),
            .I(N__15265));
    Span4Mux_v I__2864 (
            .O(N__15315),
            .I(N__15261));
    Span4Mux_h I__2863 (
            .O(N__15308),
            .I(N__15256));
    LocalMux I__2862 (
            .O(N__15301),
            .I(N__15256));
    LocalMux I__2861 (
            .O(N__15296),
            .I(N__15251));
    LocalMux I__2860 (
            .O(N__15293),
            .I(N__15251));
    LocalMux I__2859 (
            .O(N__15290),
            .I(N__15244));
    Span4Mux_v I__2858 (
            .O(N__15285),
            .I(N__15244));
    Span4Mux_v I__2857 (
            .O(N__15280),
            .I(N__15244));
    LocalMux I__2856 (
            .O(N__15277),
            .I(N__15237));
    Span4Mux_v I__2855 (
            .O(N__15272),
            .I(N__15237));
    Span4Mux_h I__2854 (
            .O(N__15265),
            .I(N__15237));
    InMux I__2853 (
            .O(N__15264),
            .I(N__15233));
    Span4Mux_h I__2852 (
            .O(N__15261),
            .I(N__15228));
    Span4Mux_v I__2851 (
            .O(N__15256),
            .I(N__15228));
    Span4Mux_h I__2850 (
            .O(N__15251),
            .I(N__15225));
    Span4Mux_h I__2849 (
            .O(N__15244),
            .I(N__15222));
    Span4Mux_v I__2848 (
            .O(N__15237),
            .I(N__15219));
    InMux I__2847 (
            .O(N__15236),
            .I(N__15216));
    LocalMux I__2846 (
            .O(N__15233),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv4 I__2845 (
            .O(N__15228),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv4 I__2844 (
            .O(N__15225),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv4 I__2843 (
            .O(N__15222),
            .I(this_vga_signals_M_vcounter_q_4));
    Odrv4 I__2842 (
            .O(N__15219),
            .I(this_vga_signals_M_vcounter_q_4));
    LocalMux I__2841 (
            .O(N__15216),
            .I(this_vga_signals_M_vcounter_q_4));
    CascadeMux I__2840 (
            .O(N__15203),
            .I(N__15198));
    InMux I__2839 (
            .O(N__15202),
            .I(N__15195));
    InMux I__2838 (
            .O(N__15201),
            .I(N__15192));
    InMux I__2837 (
            .O(N__15198),
            .I(N__15188));
    LocalMux I__2836 (
            .O(N__15195),
            .I(N__15185));
    LocalMux I__2835 (
            .O(N__15192),
            .I(N__15182));
    InMux I__2834 (
            .O(N__15191),
            .I(N__15179));
    LocalMux I__2833 (
            .O(N__15188),
            .I(N__15176));
    Span4Mux_v I__2832 (
            .O(N__15185),
            .I(N__15173));
    Span4Mux_h I__2831 (
            .O(N__15182),
            .I(N__15170));
    LocalMux I__2830 (
            .O(N__15179),
            .I(N__15167));
    Span4Mux_h I__2829 (
            .O(N__15176),
            .I(N__15164));
    Odrv4 I__2828 (
            .O(N__15173),
            .I(N_475));
    Odrv4 I__2827 (
            .O(N__15170),
            .I(N_475));
    Odrv4 I__2826 (
            .O(N__15167),
            .I(N_475));
    Odrv4 I__2825 (
            .O(N__15164),
            .I(N_475));
    CascadeMux I__2824 (
            .O(N__15155),
            .I(N__15147));
    CascadeMux I__2823 (
            .O(N__15154),
            .I(N__15144));
    CascadeMux I__2822 (
            .O(N__15153),
            .I(N__15138));
    InMux I__2821 (
            .O(N__15152),
            .I(N__15132));
    InMux I__2820 (
            .O(N__15151),
            .I(N__15129));
    InMux I__2819 (
            .O(N__15150),
            .I(N__15122));
    InMux I__2818 (
            .O(N__15147),
            .I(N__15119));
    InMux I__2817 (
            .O(N__15144),
            .I(N__15110));
    InMux I__2816 (
            .O(N__15143),
            .I(N__15110));
    InMux I__2815 (
            .O(N__15142),
            .I(N__15110));
    InMux I__2814 (
            .O(N__15141),
            .I(N__15110));
    InMux I__2813 (
            .O(N__15138),
            .I(N__15107));
    InMux I__2812 (
            .O(N__15137),
            .I(N__15101));
    InMux I__2811 (
            .O(N__15136),
            .I(N__15098));
    InMux I__2810 (
            .O(N__15135),
            .I(N__15095));
    LocalMux I__2809 (
            .O(N__15132),
            .I(N__15087));
    LocalMux I__2808 (
            .O(N__15129),
            .I(N__15087));
    InMux I__2807 (
            .O(N__15128),
            .I(N__15084));
    InMux I__2806 (
            .O(N__15127),
            .I(N__15080));
    CascadeMux I__2805 (
            .O(N__15126),
            .I(N__15077));
    CascadeMux I__2804 (
            .O(N__15125),
            .I(N__15074));
    LocalMux I__2803 (
            .O(N__15122),
            .I(N__15071));
    LocalMux I__2802 (
            .O(N__15119),
            .I(N__15068));
    LocalMux I__2801 (
            .O(N__15110),
            .I(N__15065));
    LocalMux I__2800 (
            .O(N__15107),
            .I(N__15060));
    InMux I__2799 (
            .O(N__15106),
            .I(N__15053));
    InMux I__2798 (
            .O(N__15105),
            .I(N__15053));
    InMux I__2797 (
            .O(N__15104),
            .I(N__15053));
    LocalMux I__2796 (
            .O(N__15101),
            .I(N__15050));
    LocalMux I__2795 (
            .O(N__15098),
            .I(N__15045));
    LocalMux I__2794 (
            .O(N__15095),
            .I(N__15045));
    InMux I__2793 (
            .O(N__15094),
            .I(N__15041));
    InMux I__2792 (
            .O(N__15093),
            .I(N__15038));
    InMux I__2791 (
            .O(N__15092),
            .I(N__15035));
    Span4Mux_h I__2790 (
            .O(N__15087),
            .I(N__15030));
    LocalMux I__2789 (
            .O(N__15084),
            .I(N__15030));
    InMux I__2788 (
            .O(N__15083),
            .I(N__15026));
    LocalMux I__2787 (
            .O(N__15080),
            .I(N__15023));
    InMux I__2786 (
            .O(N__15077),
            .I(N__15018));
    InMux I__2785 (
            .O(N__15074),
            .I(N__15018));
    Span4Mux_v I__2784 (
            .O(N__15071),
            .I(N__15011));
    Span4Mux_v I__2783 (
            .O(N__15068),
            .I(N__15011));
    Span4Mux_v I__2782 (
            .O(N__15065),
            .I(N__15011));
    InMux I__2781 (
            .O(N__15064),
            .I(N__15006));
    InMux I__2780 (
            .O(N__15063),
            .I(N__15006));
    Span4Mux_h I__2779 (
            .O(N__15060),
            .I(N__14997));
    LocalMux I__2778 (
            .O(N__15053),
            .I(N__14997));
    Span4Mux_v I__2777 (
            .O(N__15050),
            .I(N__14997));
    Span4Mux_h I__2776 (
            .O(N__15045),
            .I(N__14997));
    InMux I__2775 (
            .O(N__15044),
            .I(N__14994));
    LocalMux I__2774 (
            .O(N__15041),
            .I(N__14989));
    LocalMux I__2773 (
            .O(N__15038),
            .I(N__14989));
    LocalMux I__2772 (
            .O(N__15035),
            .I(N__14986));
    Span4Mux_v I__2771 (
            .O(N__15030),
            .I(N__14983));
    InMux I__2770 (
            .O(N__15029),
            .I(N__14980));
    LocalMux I__2769 (
            .O(N__15026),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv4 I__2768 (
            .O(N__15023),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__2767 (
            .O(N__15018),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv4 I__2766 (
            .O(N__15011),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__2765 (
            .O(N__15006),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv4 I__2764 (
            .O(N__14997),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__2763 (
            .O(N__14994),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv12 I__2762 (
            .O(N__14989),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv12 I__2761 (
            .O(N__14986),
            .I(this_vga_signals_M_vcounter_q_5));
    Odrv4 I__2760 (
            .O(N__14983),
            .I(this_vga_signals_M_vcounter_q_5));
    LocalMux I__2759 (
            .O(N__14980),
            .I(this_vga_signals_M_vcounter_q_5));
    InMux I__2758 (
            .O(N__14957),
            .I(N__14954));
    LocalMux I__2757 (
            .O(N__14954),
            .I(N__14951));
    Span4Mux_v I__2756 (
            .O(N__14951),
            .I(N__14948));
    Odrv4 I__2755 (
            .O(N__14948),
            .I(\this_vga_signals.N_404_0 ));
    InMux I__2754 (
            .O(N__14945),
            .I(N__14941));
    InMux I__2753 (
            .O(N__14944),
            .I(N__14938));
    LocalMux I__2752 (
            .O(N__14941),
            .I(N_204_0));
    LocalMux I__2751 (
            .O(N__14938),
            .I(N_204_0));
    InMux I__2750 (
            .O(N__14933),
            .I(\this_vga_signals.un1_M_hcounter_d_1_cry_1 ));
    CascadeMux I__2749 (
            .O(N__14930),
            .I(\this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ));
    InMux I__2748 (
            .O(N__14927),
            .I(N__14924));
    LocalMux I__2747 (
            .O(N__14924),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ));
    CascadeMux I__2746 (
            .O(N__14921),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ));
    InMux I__2745 (
            .O(N__14918),
            .I(N__14915));
    LocalMux I__2744 (
            .O(N__14915),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1 ));
    CascadeMux I__2743 (
            .O(N__14912),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_cascade_ ));
    InMux I__2742 (
            .O(N__14909),
            .I(N__14904));
    InMux I__2741 (
            .O(N__14908),
            .I(N__14899));
    InMux I__2740 (
            .O(N__14907),
            .I(N__14899));
    LocalMux I__2739 (
            .O(N__14904),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_1 ));
    LocalMux I__2738 (
            .O(N__14899),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_1 ));
    InMux I__2737 (
            .O(N__14894),
            .I(N__14891));
    LocalMux I__2736 (
            .O(N__14891),
            .I(N__14887));
    InMux I__2735 (
            .O(N__14890),
            .I(N__14884));
    Odrv4 I__2734 (
            .O(N__14887),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    LocalMux I__2733 (
            .O(N__14884),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    CascadeMux I__2732 (
            .O(N__14879),
            .I(N__14876));
    InMux I__2731 (
            .O(N__14876),
            .I(N__14873));
    LocalMux I__2730 (
            .O(N__14873),
            .I(N__14870));
    Odrv4 I__2729 (
            .O(N__14870),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ));
    InMux I__2728 (
            .O(N__14867),
            .I(N__14864));
    LocalMux I__2727 (
            .O(N__14864),
            .I(N__14859));
    InMux I__2726 (
            .O(N__14863),
            .I(N__14854));
    InMux I__2725 (
            .O(N__14862),
            .I(N__14854));
    Odrv4 I__2724 (
            .O(N__14859),
            .I(\this_vga_signals.N_336_0 ));
    LocalMux I__2723 (
            .O(N__14854),
            .I(\this_vga_signals.N_336_0 ));
    CascadeMux I__2722 (
            .O(N__14849),
            .I(\this_vga_signals.N_336_0_cascade_ ));
    InMux I__2721 (
            .O(N__14846),
            .I(N__14840));
    InMux I__2720 (
            .O(N__14845),
            .I(N__14833));
    InMux I__2719 (
            .O(N__14844),
            .I(N__14833));
    InMux I__2718 (
            .O(N__14843),
            .I(N__14833));
    LocalMux I__2717 (
            .O(N__14840),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ));
    LocalMux I__2716 (
            .O(N__14833),
            .I(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ));
    InMux I__2715 (
            .O(N__14828),
            .I(N__14825));
    LocalMux I__2714 (
            .O(N__14825),
            .I(\this_vga_signals.N_287 ));
    CascadeMux I__2713 (
            .O(N__14822),
            .I(\this_vga_signals.N_287_cascade_ ));
    InMux I__2712 (
            .O(N__14819),
            .I(N__14816));
    LocalMux I__2711 (
            .O(N__14816),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0 ));
    CascadeMux I__2710 (
            .O(N__14813),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ));
    CascadeMux I__2709 (
            .O(N__14810),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3_cascade_));
    CascadeMux I__2708 (
            .O(N__14807),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_1_cascade_ ));
    InMux I__2707 (
            .O(N__14804),
            .I(N__14794));
    InMux I__2706 (
            .O(N__14803),
            .I(N__14794));
    InMux I__2705 (
            .O(N__14802),
            .I(N__14794));
    InMux I__2704 (
            .O(N__14801),
            .I(N__14791));
    LocalMux I__2703 (
            .O(N__14794),
            .I(\this_vga_signals.SUM_7_i_1_0 ));
    LocalMux I__2702 (
            .O(N__14791),
            .I(\this_vga_signals.SUM_7_i_1_0 ));
    CascadeMux I__2701 (
            .O(N__14786),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ));
    InMux I__2700 (
            .O(N__14783),
            .I(N__14780));
    LocalMux I__2699 (
            .O(N__14780),
            .I(G_504));
    CascadeMux I__2698 (
            .O(N__14777),
            .I(N__14774));
    InMux I__2697 (
            .O(N__14774),
            .I(N__14771));
    LocalMux I__2696 (
            .O(N__14771),
            .I(N__14768));
    Span4Mux_v I__2695 (
            .O(N__14768),
            .I(N__14765));
    Odrv4 I__2694 (
            .O(N__14765),
            .I(\this_vga_signals.mult1_un68_sum_cry_1_s ));
    InMux I__2693 (
            .O(N__14762),
            .I(N__14759));
    LocalMux I__2692 (
            .O(N__14759),
            .I(G_503));
    InMux I__2691 (
            .O(N__14756),
            .I(N__14753));
    LocalMux I__2690 (
            .O(N__14753),
            .I(N__14750));
    Odrv4 I__2689 (
            .O(N__14750),
            .I(\this_vga_signals.mult1_un75_sum_axb_3 ));
    InMux I__2688 (
            .O(N__14747),
            .I(\this_vga_signals.mult1_un75_sum_cry_2 ));
    CascadeMux I__2687 (
            .O(N__14744),
            .I(\this_ppu.M_m12_0_o2_381Z0Z_4_cascade_ ));
    InMux I__2686 (
            .O(N__14741),
            .I(N__14737));
    InMux I__2685 (
            .O(N__14740),
            .I(N__14734));
    LocalMux I__2684 (
            .O(N__14737),
            .I(N__14731));
    LocalMux I__2683 (
            .O(N__14734),
            .I(N_275));
    Odrv4 I__2682 (
            .O(N__14731),
            .I(N_275));
    CascadeMux I__2681 (
            .O(N__14726),
            .I(\this_ppu.M_m12_0_o2_381_5_cascade_ ));
    InMux I__2680 (
            .O(N__14723),
            .I(N__14720));
    LocalMux I__2679 (
            .O(N__14720),
            .I(N__14717));
    Span4Mux_h I__2678 (
            .O(N__14717),
            .I(N__14712));
    InMux I__2677 (
            .O(N__14716),
            .I(N__14709));
    InMux I__2676 (
            .O(N__14715),
            .I(N__14706));
    Odrv4 I__2675 (
            .O(N__14712),
            .I(N_190_0));
    LocalMux I__2674 (
            .O(N__14709),
            .I(N_190_0));
    LocalMux I__2673 (
            .O(N__14706),
            .I(N_190_0));
    InMux I__2672 (
            .O(N__14699),
            .I(N__14696));
    LocalMux I__2671 (
            .O(N__14696),
            .I(N__14693));
    Span4Mux_h I__2670 (
            .O(N__14693),
            .I(N__14690));
    Odrv4 I__2669 (
            .O(N__14690),
            .I(\this_ppu.M_m12_0_o2_381_8 ));
    InMux I__2668 (
            .O(N__14687),
            .I(N__14682));
    InMux I__2667 (
            .O(N__14686),
            .I(N__14677));
    InMux I__2666 (
            .O(N__14685),
            .I(N__14677));
    LocalMux I__2665 (
            .O(N__14682),
            .I(M_this_delay_clk_out_0));
    LocalMux I__2664 (
            .O(N__14677),
            .I(M_this_delay_clk_out_0));
    InMux I__2663 (
            .O(N__14672),
            .I(N__14665));
    InMux I__2662 (
            .O(N__14671),
            .I(N__14665));
    InMux I__2661 (
            .O(N__14670),
            .I(N__14662));
    LocalMux I__2660 (
            .O(N__14665),
            .I(N__14657));
    LocalMux I__2659 (
            .O(N__14662),
            .I(N__14657));
    Span4Mux_v I__2658 (
            .O(N__14657),
            .I(N__14654));
    Span4Mux_h I__2657 (
            .O(N__14654),
            .I(N__14651));
    Span4Mux_h I__2656 (
            .O(N__14651),
            .I(N__14648));
    Odrv4 I__2655 (
            .O(N__14648),
            .I(port_enb_c));
    InMux I__2654 (
            .O(N__14645),
            .I(N__14642));
    LocalMux I__2653 (
            .O(N__14642),
            .I(N__14638));
    InMux I__2652 (
            .O(N__14641),
            .I(N__14635));
    Odrv4 I__2651 (
            .O(N__14638),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__2650 (
            .O(N__14635),
            .I(this_start_data_delay_M_last_q));
    InMux I__2649 (
            .O(N__14630),
            .I(N__14627));
    LocalMux I__2648 (
            .O(N__14627),
            .I(\this_vga_signals.mult1_un61_sum_i_0 ));
    InMux I__2647 (
            .O(N__14624),
            .I(N__14620));
    InMux I__2646 (
            .O(N__14623),
            .I(N__14617));
    LocalMux I__2645 (
            .O(N__14620),
            .I(N__14614));
    LocalMux I__2644 (
            .O(N__14617),
            .I(N__14611));
    Span4Mux_h I__2643 (
            .O(N__14614),
            .I(N__14608));
    Span4Mux_h I__2642 (
            .O(N__14611),
            .I(N__14605));
    Span4Mux_v I__2641 (
            .O(N__14608),
            .I(N__14602));
    Odrv4 I__2640 (
            .O(N__14605),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_0 ));
    Odrv4 I__2639 (
            .O(N__14602),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_0 ));
    CascadeMux I__2638 (
            .O(N__14597),
            .I(N__14594));
    InMux I__2637 (
            .O(N__14594),
            .I(N__14591));
    LocalMux I__2636 (
            .O(N__14591),
            .I(N__14588));
    Span12Mux_h I__2635 (
            .O(N__14588),
            .I(N__14585));
    Odrv12 I__2634 (
            .O(N__14585),
            .I(N_90_0));
    CascadeMux I__2633 (
            .O(N__14582),
            .I(N__14569));
    CascadeMux I__2632 (
            .O(N__14581),
            .I(N__14566));
    CascadeMux I__2631 (
            .O(N__14580),
            .I(N__14558));
    CascadeMux I__2630 (
            .O(N__14579),
            .I(N__14552));
    CascadeMux I__2629 (
            .O(N__14578),
            .I(N__14548));
    CascadeMux I__2628 (
            .O(N__14577),
            .I(N__14545));
    CascadeMux I__2627 (
            .O(N__14576),
            .I(N__14542));
    InMux I__2626 (
            .O(N__14575),
            .I(N__14535));
    InMux I__2625 (
            .O(N__14574),
            .I(N__14535));
    InMux I__2624 (
            .O(N__14573),
            .I(N__14532));
    InMux I__2623 (
            .O(N__14572),
            .I(N__14526));
    InMux I__2622 (
            .O(N__14569),
            .I(N__14526));
    InMux I__2621 (
            .O(N__14566),
            .I(N__14519));
    InMux I__2620 (
            .O(N__14565),
            .I(N__14519));
    InMux I__2619 (
            .O(N__14564),
            .I(N__14519));
    InMux I__2618 (
            .O(N__14563),
            .I(N__14514));
    InMux I__2617 (
            .O(N__14562),
            .I(N__14514));
    CascadeMux I__2616 (
            .O(N__14561),
            .I(N__14509));
    InMux I__2615 (
            .O(N__14558),
            .I(N__14506));
    InMux I__2614 (
            .O(N__14557),
            .I(N__14499));
    InMux I__2613 (
            .O(N__14556),
            .I(N__14499));
    InMux I__2612 (
            .O(N__14555),
            .I(N__14499));
    InMux I__2611 (
            .O(N__14552),
            .I(N__14495));
    InMux I__2610 (
            .O(N__14551),
            .I(N__14488));
    InMux I__2609 (
            .O(N__14548),
            .I(N__14488));
    InMux I__2608 (
            .O(N__14545),
            .I(N__14488));
    InMux I__2607 (
            .O(N__14542),
            .I(N__14483));
    InMux I__2606 (
            .O(N__14541),
            .I(N__14483));
    InMux I__2605 (
            .O(N__14540),
            .I(N__14480));
    LocalMux I__2604 (
            .O(N__14535),
            .I(N__14475));
    LocalMux I__2603 (
            .O(N__14532),
            .I(N__14475));
    InMux I__2602 (
            .O(N__14531),
            .I(N__14472));
    LocalMux I__2601 (
            .O(N__14526),
            .I(N__14465));
    LocalMux I__2600 (
            .O(N__14519),
            .I(N__14465));
    LocalMux I__2599 (
            .O(N__14514),
            .I(N__14462));
    InMux I__2598 (
            .O(N__14513),
            .I(N__14459));
    InMux I__2597 (
            .O(N__14512),
            .I(N__14454));
    InMux I__2596 (
            .O(N__14509),
            .I(N__14454));
    LocalMux I__2595 (
            .O(N__14506),
            .I(N__14449));
    LocalMux I__2594 (
            .O(N__14499),
            .I(N__14449));
    InMux I__2593 (
            .O(N__14498),
            .I(N__14446));
    LocalMux I__2592 (
            .O(N__14495),
            .I(N__14443));
    LocalMux I__2591 (
            .O(N__14488),
            .I(N__14434));
    LocalMux I__2590 (
            .O(N__14483),
            .I(N__14434));
    LocalMux I__2589 (
            .O(N__14480),
            .I(N__14434));
    Span4Mux_h I__2588 (
            .O(N__14475),
            .I(N__14434));
    LocalMux I__2587 (
            .O(N__14472),
            .I(N__14431));
    InMux I__2586 (
            .O(N__14471),
            .I(N__14428));
    InMux I__2585 (
            .O(N__14470),
            .I(N__14425));
    Span4Mux_v I__2584 (
            .O(N__14465),
            .I(N__14420));
    Span4Mux_h I__2583 (
            .O(N__14462),
            .I(N__14420));
    LocalMux I__2582 (
            .O(N__14459),
            .I(N__14415));
    LocalMux I__2581 (
            .O(N__14454),
            .I(N__14415));
    Span4Mux_v I__2580 (
            .O(N__14449),
            .I(N__14410));
    LocalMux I__2579 (
            .O(N__14446),
            .I(N__14410));
    Span4Mux_v I__2578 (
            .O(N__14443),
            .I(N__14403));
    Span4Mux_v I__2577 (
            .O(N__14434),
            .I(N__14403));
    Span4Mux_v I__2576 (
            .O(N__14431),
            .I(N__14403));
    LocalMux I__2575 (
            .O(N__14428),
            .I(N__14400));
    LocalMux I__2574 (
            .O(N__14425),
            .I(this_vga_signals_M_vcounter_q_2));
    Odrv4 I__2573 (
            .O(N__14420),
            .I(this_vga_signals_M_vcounter_q_2));
    Odrv12 I__2572 (
            .O(N__14415),
            .I(this_vga_signals_M_vcounter_q_2));
    Odrv4 I__2571 (
            .O(N__14410),
            .I(this_vga_signals_M_vcounter_q_2));
    Odrv4 I__2570 (
            .O(N__14403),
            .I(this_vga_signals_M_vcounter_q_2));
    Odrv4 I__2569 (
            .O(N__14400),
            .I(this_vga_signals_M_vcounter_q_2));
    CascadeMux I__2568 (
            .O(N__14387),
            .I(N__14380));
    CascadeMux I__2567 (
            .O(N__14386),
            .I(N__14362));
    CascadeMux I__2566 (
            .O(N__14385),
            .I(N__14359));
    InMux I__2565 (
            .O(N__14384),
            .I(N__14356));
    InMux I__2564 (
            .O(N__14383),
            .I(N__14351));
    InMux I__2563 (
            .O(N__14380),
            .I(N__14351));
    InMux I__2562 (
            .O(N__14379),
            .I(N__14348));
    InMux I__2561 (
            .O(N__14378),
            .I(N__14339));
    InMux I__2560 (
            .O(N__14377),
            .I(N__14336));
    InMux I__2559 (
            .O(N__14376),
            .I(N__14330));
    InMux I__2558 (
            .O(N__14375),
            .I(N__14327));
    InMux I__2557 (
            .O(N__14374),
            .I(N__14324));
    InMux I__2556 (
            .O(N__14373),
            .I(N__14321));
    InMux I__2555 (
            .O(N__14372),
            .I(N__14312));
    InMux I__2554 (
            .O(N__14371),
            .I(N__14312));
    InMux I__2553 (
            .O(N__14370),
            .I(N__14312));
    InMux I__2552 (
            .O(N__14369),
            .I(N__14312));
    InMux I__2551 (
            .O(N__14368),
            .I(N__14307));
    InMux I__2550 (
            .O(N__14367),
            .I(N__14307));
    InMux I__2549 (
            .O(N__14366),
            .I(N__14296));
    InMux I__2548 (
            .O(N__14365),
            .I(N__14296));
    InMux I__2547 (
            .O(N__14362),
            .I(N__14291));
    InMux I__2546 (
            .O(N__14359),
            .I(N__14291));
    LocalMux I__2545 (
            .O(N__14356),
            .I(N__14284));
    LocalMux I__2544 (
            .O(N__14351),
            .I(N__14284));
    LocalMux I__2543 (
            .O(N__14348),
            .I(N__14284));
    InMux I__2542 (
            .O(N__14347),
            .I(N__14281));
    InMux I__2541 (
            .O(N__14346),
            .I(N__14276));
    InMux I__2540 (
            .O(N__14345),
            .I(N__14276));
    InMux I__2539 (
            .O(N__14344),
            .I(N__14271));
    InMux I__2538 (
            .O(N__14343),
            .I(N__14271));
    InMux I__2537 (
            .O(N__14342),
            .I(N__14267));
    LocalMux I__2536 (
            .O(N__14339),
            .I(N__14262));
    LocalMux I__2535 (
            .O(N__14336),
            .I(N__14262));
    InMux I__2534 (
            .O(N__14335),
            .I(N__14259));
    InMux I__2533 (
            .O(N__14334),
            .I(N__14256));
    InMux I__2532 (
            .O(N__14333),
            .I(N__14251));
    LocalMux I__2531 (
            .O(N__14330),
            .I(N__14242));
    LocalMux I__2530 (
            .O(N__14327),
            .I(N__14242));
    LocalMux I__2529 (
            .O(N__14324),
            .I(N__14242));
    LocalMux I__2528 (
            .O(N__14321),
            .I(N__14242));
    LocalMux I__2527 (
            .O(N__14312),
            .I(N__14237));
    LocalMux I__2526 (
            .O(N__14307),
            .I(N__14237));
    InMux I__2525 (
            .O(N__14306),
            .I(N__14234));
    InMux I__2524 (
            .O(N__14305),
            .I(N__14227));
    InMux I__2523 (
            .O(N__14304),
            .I(N__14227));
    InMux I__2522 (
            .O(N__14303),
            .I(N__14227));
    InMux I__2521 (
            .O(N__14302),
            .I(N__14224));
    InMux I__2520 (
            .O(N__14301),
            .I(N__14221));
    LocalMux I__2519 (
            .O(N__14296),
            .I(N__14214));
    LocalMux I__2518 (
            .O(N__14291),
            .I(N__14214));
    Span4Mux_h I__2517 (
            .O(N__14284),
            .I(N__14214));
    LocalMux I__2516 (
            .O(N__14281),
            .I(N__14207));
    LocalMux I__2515 (
            .O(N__14276),
            .I(N__14207));
    LocalMux I__2514 (
            .O(N__14271),
            .I(N__14207));
    InMux I__2513 (
            .O(N__14270),
            .I(N__14204));
    LocalMux I__2512 (
            .O(N__14267),
            .I(N__14197));
    Span4Mux_v I__2511 (
            .O(N__14262),
            .I(N__14197));
    LocalMux I__2510 (
            .O(N__14259),
            .I(N__14197));
    LocalMux I__2509 (
            .O(N__14256),
            .I(N__14194));
    InMux I__2508 (
            .O(N__14255),
            .I(N__14191));
    InMux I__2507 (
            .O(N__14254),
            .I(N__14188));
    LocalMux I__2506 (
            .O(N__14251),
            .I(N__14185));
    Span4Mux_v I__2505 (
            .O(N__14242),
            .I(N__14180));
    Span4Mux_h I__2504 (
            .O(N__14237),
            .I(N__14180));
    LocalMux I__2503 (
            .O(N__14234),
            .I(N__14173));
    LocalMux I__2502 (
            .O(N__14227),
            .I(N__14173));
    LocalMux I__2501 (
            .O(N__14224),
            .I(N__14173));
    LocalMux I__2500 (
            .O(N__14221),
            .I(N__14164));
    Span4Mux_v I__2499 (
            .O(N__14214),
            .I(N__14164));
    Span4Mux_v I__2498 (
            .O(N__14207),
            .I(N__14164));
    LocalMux I__2497 (
            .O(N__14204),
            .I(N__14164));
    Span4Mux_v I__2496 (
            .O(N__14197),
            .I(N__14157));
    Span4Mux_v I__2495 (
            .O(N__14194),
            .I(N__14157));
    LocalMux I__2494 (
            .O(N__14191),
            .I(N__14157));
    LocalMux I__2493 (
            .O(N__14188),
            .I(this_vga_signals_M_vcounter_q_3));
    Odrv12 I__2492 (
            .O(N__14185),
            .I(this_vga_signals_M_vcounter_q_3));
    Odrv4 I__2491 (
            .O(N__14180),
            .I(this_vga_signals_M_vcounter_q_3));
    Odrv4 I__2490 (
            .O(N__14173),
            .I(this_vga_signals_M_vcounter_q_3));
    Odrv4 I__2489 (
            .O(N__14164),
            .I(this_vga_signals_M_vcounter_q_3));
    Odrv4 I__2488 (
            .O(N__14157),
            .I(this_vga_signals_M_vcounter_q_3));
    InMux I__2487 (
            .O(N__14144),
            .I(N__14141));
    LocalMux I__2486 (
            .O(N__14141),
            .I(N__14138));
    Span4Mux_h I__2485 (
            .O(N__14138),
            .I(N__14135));
    Odrv4 I__2484 (
            .O(N__14135),
            .I(N_184_0));
    CascadeMux I__2483 (
            .O(N__14132),
            .I(N__14123));
    InMux I__2482 (
            .O(N__14131),
            .I(N__14119));
    InMux I__2481 (
            .O(N__14130),
            .I(N__14115));
    CascadeMux I__2480 (
            .O(N__14129),
            .I(N__14110));
    InMux I__2479 (
            .O(N__14128),
            .I(N__14104));
    InMux I__2478 (
            .O(N__14127),
            .I(N__14101));
    InMux I__2477 (
            .O(N__14126),
            .I(N__14098));
    InMux I__2476 (
            .O(N__14123),
            .I(N__14095));
    InMux I__2475 (
            .O(N__14122),
            .I(N__14092));
    LocalMux I__2474 (
            .O(N__14119),
            .I(N__14088));
    InMux I__2473 (
            .O(N__14118),
            .I(N__14085));
    LocalMux I__2472 (
            .O(N__14115),
            .I(N__14082));
    InMux I__2471 (
            .O(N__14114),
            .I(N__14075));
    InMux I__2470 (
            .O(N__14113),
            .I(N__14075));
    InMux I__2469 (
            .O(N__14110),
            .I(N__14075));
    InMux I__2468 (
            .O(N__14109),
            .I(N__14068));
    InMux I__2467 (
            .O(N__14108),
            .I(N__14068));
    InMux I__2466 (
            .O(N__14107),
            .I(N__14068));
    LocalMux I__2465 (
            .O(N__14104),
            .I(N__14063));
    LocalMux I__2464 (
            .O(N__14101),
            .I(N__14060));
    LocalMux I__2463 (
            .O(N__14098),
            .I(N__14057));
    LocalMux I__2462 (
            .O(N__14095),
            .I(N__14054));
    LocalMux I__2461 (
            .O(N__14092),
            .I(N__14051));
    InMux I__2460 (
            .O(N__14091),
            .I(N__14048));
    Span4Mux_h I__2459 (
            .O(N__14088),
            .I(N__14045));
    LocalMux I__2458 (
            .O(N__14085),
            .I(N__14042));
    Span4Mux_v I__2457 (
            .O(N__14082),
            .I(N__14035));
    LocalMux I__2456 (
            .O(N__14075),
            .I(N__14035));
    LocalMux I__2455 (
            .O(N__14068),
            .I(N__14035));
    InMux I__2454 (
            .O(N__14067),
            .I(N__14032));
    InMux I__2453 (
            .O(N__14066),
            .I(N__14029));
    Span4Mux_v I__2452 (
            .O(N__14063),
            .I(N__14022));
    Span4Mux_v I__2451 (
            .O(N__14060),
            .I(N__14022));
    Span4Mux_v I__2450 (
            .O(N__14057),
            .I(N__14022));
    Span4Mux_v I__2449 (
            .O(N__14054),
            .I(N__14017));
    Span4Mux_v I__2448 (
            .O(N__14051),
            .I(N__14017));
    LocalMux I__2447 (
            .O(N__14048),
            .I(N__14014));
    Span4Mux_v I__2446 (
            .O(N__14045),
            .I(N__14007));
    Span4Mux_v I__2445 (
            .O(N__14042),
            .I(N__14007));
    Span4Mux_v I__2444 (
            .O(N__14035),
            .I(N__14007));
    LocalMux I__2443 (
            .O(N__14032),
            .I(N__14004));
    LocalMux I__2442 (
            .O(N__14029),
            .I(this_vga_signals_M_vcounter_q_1));
    Odrv4 I__2441 (
            .O(N__14022),
            .I(this_vga_signals_M_vcounter_q_1));
    Odrv4 I__2440 (
            .O(N__14017),
            .I(this_vga_signals_M_vcounter_q_1));
    Odrv12 I__2439 (
            .O(N__14014),
            .I(this_vga_signals_M_vcounter_q_1));
    Odrv4 I__2438 (
            .O(N__14007),
            .I(this_vga_signals_M_vcounter_q_1));
    Odrv12 I__2437 (
            .O(N__14004),
            .I(this_vga_signals_M_vcounter_q_1));
    CascadeMux I__2436 (
            .O(N__13991),
            .I(N_184_0_cascade_));
    CascadeMux I__2435 (
            .O(N__13988),
            .I(N__13982));
    InMux I__2434 (
            .O(N__13987),
            .I(N__13978));
    InMux I__2433 (
            .O(N__13986),
            .I(N__13974));
    InMux I__2432 (
            .O(N__13985),
            .I(N__13967));
    InMux I__2431 (
            .O(N__13982),
            .I(N__13967));
    InMux I__2430 (
            .O(N__13981),
            .I(N__13967));
    LocalMux I__2429 (
            .O(N__13978),
            .I(N__13962));
    InMux I__2428 (
            .O(N__13977),
            .I(N__13959));
    LocalMux I__2427 (
            .O(N__13974),
            .I(N__13954));
    LocalMux I__2426 (
            .O(N__13967),
            .I(N__13954));
    InMux I__2425 (
            .O(N__13966),
            .I(N__13951));
    InMux I__2424 (
            .O(N__13965),
            .I(N__13948));
    Sp12to4 I__2423 (
            .O(N__13962),
            .I(N__13943));
    LocalMux I__2422 (
            .O(N__13959),
            .I(N__13943));
    Span4Mux_v I__2421 (
            .O(N__13954),
            .I(N__13938));
    LocalMux I__2420 (
            .O(N__13951),
            .I(N__13938));
    LocalMux I__2419 (
            .O(N__13948),
            .I(this_vga_signals_M_vcounter_q_0));
    Odrv12 I__2418 (
            .O(N__13943),
            .I(this_vga_signals_M_vcounter_q_0));
    Odrv4 I__2417 (
            .O(N__13938),
            .I(this_vga_signals_M_vcounter_q_0));
    InMux I__2416 (
            .O(N__13931),
            .I(N__13920));
    InMux I__2415 (
            .O(N__13930),
            .I(N__13913));
    InMux I__2414 (
            .O(N__13929),
            .I(N__13913));
    InMux I__2413 (
            .O(N__13928),
            .I(N__13913));
    InMux I__2412 (
            .O(N__13927),
            .I(N__13908));
    InMux I__2411 (
            .O(N__13926),
            .I(N__13903));
    InMux I__2410 (
            .O(N__13925),
            .I(N__13903));
    InMux I__2409 (
            .O(N__13924),
            .I(N__13900));
    InMux I__2408 (
            .O(N__13923),
            .I(N__13897));
    LocalMux I__2407 (
            .O(N__13920),
            .I(N__13892));
    LocalMux I__2406 (
            .O(N__13913),
            .I(N__13892));
    InMux I__2405 (
            .O(N__13912),
            .I(N__13887));
    InMux I__2404 (
            .O(N__13911),
            .I(N__13887));
    LocalMux I__2403 (
            .O(N__13908),
            .I(N__13881));
    LocalMux I__2402 (
            .O(N__13903),
            .I(N__13874));
    LocalMux I__2401 (
            .O(N__13900),
            .I(N__13874));
    LocalMux I__2400 (
            .O(N__13897),
            .I(N__13874));
    Span4Mux_v I__2399 (
            .O(N__13892),
            .I(N__13869));
    LocalMux I__2398 (
            .O(N__13887),
            .I(N__13869));
    InMux I__2397 (
            .O(N__13886),
            .I(N__13866));
    InMux I__2396 (
            .O(N__13885),
            .I(N__13863));
    InMux I__2395 (
            .O(N__13884),
            .I(N__13860));
    Odrv4 I__2394 (
            .O(N__13881),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__2393 (
            .O(N__13874),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__2392 (
            .O(N__13869),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2391 (
            .O(N__13866),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2390 (
            .O(N__13863),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__2389 (
            .O(N__13860),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    InMux I__2388 (
            .O(N__13847),
            .I(N__13844));
    LocalMux I__2387 (
            .O(N__13844),
            .I(\this_vga_signals.if_N_8_0 ));
    InMux I__2386 (
            .O(N__13841),
            .I(N__13838));
    LocalMux I__2385 (
            .O(N__13838),
            .I(N__13835));
    Span4Mux_v I__2384 (
            .O(N__13835),
            .I(N__13832));
    Odrv4 I__2383 (
            .O(N__13832),
            .I(\this_vga_signals.mult1_un54_sum_i_0 ));
    IoInMux I__2382 (
            .O(N__13829),
            .I(N__13826));
    LocalMux I__2381 (
            .O(N__13826),
            .I(N__13823));
    IoSpan4Mux I__2380 (
            .O(N__13823),
            .I(N__13820));
    IoSpan4Mux I__2379 (
            .O(N__13820),
            .I(N__13817));
    Span4Mux_s2_v I__2378 (
            .O(N__13817),
            .I(N__13814));
    Sp12to4 I__2377 (
            .O(N__13814),
            .I(N__13811));
    Span12Mux_v I__2376 (
            .O(N__13811),
            .I(N__13808));
    Odrv12 I__2375 (
            .O(N__13808),
            .I(N_31));
    InMux I__2374 (
            .O(N__13805),
            .I(N__13794));
    InMux I__2373 (
            .O(N__13804),
            .I(N__13785));
    InMux I__2372 (
            .O(N__13803),
            .I(N__13782));
    InMux I__2371 (
            .O(N__13802),
            .I(N__13777));
    InMux I__2370 (
            .O(N__13801),
            .I(N__13777));
    InMux I__2369 (
            .O(N__13800),
            .I(N__13774));
    InMux I__2368 (
            .O(N__13799),
            .I(N__13770));
    InMux I__2367 (
            .O(N__13798),
            .I(N__13767));
    InMux I__2366 (
            .O(N__13797),
            .I(N__13764));
    LocalMux I__2365 (
            .O(N__13794),
            .I(N__13761));
    InMux I__2364 (
            .O(N__13793),
            .I(N__13758));
    InMux I__2363 (
            .O(N__13792),
            .I(N__13751));
    InMux I__2362 (
            .O(N__13791),
            .I(N__13751));
    InMux I__2361 (
            .O(N__13790),
            .I(N__13751));
    InMux I__2360 (
            .O(N__13789),
            .I(N__13746));
    InMux I__2359 (
            .O(N__13788),
            .I(N__13746));
    LocalMux I__2358 (
            .O(N__13785),
            .I(N__13743));
    LocalMux I__2357 (
            .O(N__13782),
            .I(N__13736));
    LocalMux I__2356 (
            .O(N__13777),
            .I(N__13736));
    LocalMux I__2355 (
            .O(N__13774),
            .I(N__13736));
    InMux I__2354 (
            .O(N__13773),
            .I(N__13733));
    LocalMux I__2353 (
            .O(N__13770),
            .I(N__13728));
    LocalMux I__2352 (
            .O(N__13767),
            .I(N__13728));
    LocalMux I__2351 (
            .O(N__13764),
            .I(N__13723));
    Span4Mux_v I__2350 (
            .O(N__13761),
            .I(N__13723));
    LocalMux I__2349 (
            .O(N__13758),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2348 (
            .O(N__13751),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2347 (
            .O(N__13746),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2346 (
            .O(N__13743),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2345 (
            .O(N__13736),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2344 (
            .O(N__13733),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2343 (
            .O(N__13728),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2342 (
            .O(N__13723),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__2341 (
            .O(N__13706),
            .I(N__13702));
    CascadeMux I__2340 (
            .O(N__13705),
            .I(N__13694));
    LocalMux I__2339 (
            .O(N__13702),
            .I(N__13691));
    CascadeMux I__2338 (
            .O(N__13701),
            .I(N__13687));
    InMux I__2337 (
            .O(N__13700),
            .I(N__13684));
    InMux I__2336 (
            .O(N__13699),
            .I(N__13678));
    InMux I__2335 (
            .O(N__13698),
            .I(N__13678));
    InMux I__2334 (
            .O(N__13697),
            .I(N__13669));
    InMux I__2333 (
            .O(N__13694),
            .I(N__13669));
    Span4Mux_v I__2332 (
            .O(N__13691),
            .I(N__13666));
    InMux I__2331 (
            .O(N__13690),
            .I(N__13663));
    InMux I__2330 (
            .O(N__13687),
            .I(N__13660));
    LocalMux I__2329 (
            .O(N__13684),
            .I(N__13657));
    InMux I__2328 (
            .O(N__13683),
            .I(N__13652));
    LocalMux I__2327 (
            .O(N__13678),
            .I(N__13648));
    InMux I__2326 (
            .O(N__13677),
            .I(N__13645));
    InMux I__2325 (
            .O(N__13676),
            .I(N__13642));
    InMux I__2324 (
            .O(N__13675),
            .I(N__13637));
    InMux I__2323 (
            .O(N__13674),
            .I(N__13637));
    LocalMux I__2322 (
            .O(N__13669),
            .I(N__13634));
    Span4Mux_v I__2321 (
            .O(N__13666),
            .I(N__13629));
    LocalMux I__2320 (
            .O(N__13663),
            .I(N__13629));
    LocalMux I__2319 (
            .O(N__13660),
            .I(N__13626));
    Span4Mux_h I__2318 (
            .O(N__13657),
            .I(N__13623));
    InMux I__2317 (
            .O(N__13656),
            .I(N__13618));
    InMux I__2316 (
            .O(N__13655),
            .I(N__13618));
    LocalMux I__2315 (
            .O(N__13652),
            .I(N__13615));
    InMux I__2314 (
            .O(N__13651),
            .I(N__13612));
    Span4Mux_h I__2313 (
            .O(N__13648),
            .I(N__13601));
    LocalMux I__2312 (
            .O(N__13645),
            .I(N__13601));
    LocalMux I__2311 (
            .O(N__13642),
            .I(N__13601));
    LocalMux I__2310 (
            .O(N__13637),
            .I(N__13601));
    Span4Mux_h I__2309 (
            .O(N__13634),
            .I(N__13601));
    Odrv4 I__2308 (
            .O(N__13629),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv12 I__2307 (
            .O(N__13626),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv4 I__2306 (
            .O(N__13623),
            .I(this_vga_signals_M_vcounter_q_6));
    LocalMux I__2305 (
            .O(N__13618),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv4 I__2304 (
            .O(N__13615),
            .I(this_vga_signals_M_vcounter_q_6));
    LocalMux I__2303 (
            .O(N__13612),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv4 I__2302 (
            .O(N__13601),
            .I(this_vga_signals_M_vcounter_q_6));
    CascadeMux I__2301 (
            .O(N__13586),
            .I(N__13579));
    InMux I__2300 (
            .O(N__13585),
            .I(N__13575));
    InMux I__2299 (
            .O(N__13584),
            .I(N__13572));
    InMux I__2298 (
            .O(N__13583),
            .I(N__13569));
    InMux I__2297 (
            .O(N__13582),
            .I(N__13564));
    InMux I__2296 (
            .O(N__13579),
            .I(N__13561));
    InMux I__2295 (
            .O(N__13578),
            .I(N__13558));
    LocalMux I__2294 (
            .O(N__13575),
            .I(N__13551));
    LocalMux I__2293 (
            .O(N__13572),
            .I(N__13546));
    LocalMux I__2292 (
            .O(N__13569),
            .I(N__13546));
    InMux I__2291 (
            .O(N__13568),
            .I(N__13539));
    InMux I__2290 (
            .O(N__13567),
            .I(N__13539));
    LocalMux I__2289 (
            .O(N__13564),
            .I(N__13534));
    LocalMux I__2288 (
            .O(N__13561),
            .I(N__13534));
    LocalMux I__2287 (
            .O(N__13558),
            .I(N__13531));
    InMux I__2286 (
            .O(N__13557),
            .I(N__13528));
    InMux I__2285 (
            .O(N__13556),
            .I(N__13523));
    InMux I__2284 (
            .O(N__13555),
            .I(N__13523));
    InMux I__2283 (
            .O(N__13554),
            .I(N__13520));
    Span4Mux_v I__2282 (
            .O(N__13551),
            .I(N__13515));
    Span4Mux_v I__2281 (
            .O(N__13546),
            .I(N__13515));
    InMux I__2280 (
            .O(N__13545),
            .I(N__13510));
    InMux I__2279 (
            .O(N__13544),
            .I(N__13510));
    LocalMux I__2278 (
            .O(N__13539),
            .I(N__13507));
    Odrv4 I__2277 (
            .O(N__13534),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2276 (
            .O(N__13531),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2275 (
            .O(N__13528),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2274 (
            .O(N__13523),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2273 (
            .O(N__13520),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2272 (
            .O(N__13515),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2271 (
            .O(N__13510),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    Odrv4 I__2270 (
            .O(N__13507),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    CascadeMux I__2269 (
            .O(N__13490),
            .I(\this_vga_signals.N_177_0_cascade_ ));
    InMux I__2268 (
            .O(N__13487),
            .I(N__13482));
    InMux I__2267 (
            .O(N__13486),
            .I(N__13478));
    CascadeMux I__2266 (
            .O(N__13485),
            .I(N__13475));
    LocalMux I__2265 (
            .O(N__13482),
            .I(N__13472));
    InMux I__2264 (
            .O(N__13481),
            .I(N__13469));
    LocalMux I__2263 (
            .O(N__13478),
            .I(N__13466));
    InMux I__2262 (
            .O(N__13475),
            .I(N__13463));
    Span4Mux_v I__2261 (
            .O(N__13472),
            .I(N__13458));
    LocalMux I__2260 (
            .O(N__13469),
            .I(N__13458));
    Span4Mux_v I__2259 (
            .O(N__13466),
            .I(N__13453));
    LocalMux I__2258 (
            .O(N__13463),
            .I(N__13453));
    Span4Mux_h I__2257 (
            .O(N__13458),
            .I(N__13450));
    Span4Mux_v I__2256 (
            .O(N__13453),
            .I(N__13447));
    Span4Mux_v I__2255 (
            .O(N__13450),
            .I(N__13444));
    Odrv4 I__2254 (
            .O(N__13447),
            .I(\this_vga_signals.CO0_i_0 ));
    Odrv4 I__2253 (
            .O(N__13444),
            .I(\this_vga_signals.CO0_i_0 ));
    InMux I__2252 (
            .O(N__13439),
            .I(N__13436));
    LocalMux I__2251 (
            .O(N__13436),
            .I(\this_vga_signals.N_269_0 ));
    InMux I__2250 (
            .O(N__13433),
            .I(N__13430));
    LocalMux I__2249 (
            .O(N__13430),
            .I(\this_vga_signals.N_286 ));
    CascadeMux I__2248 (
            .O(N__13427),
            .I(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1_cascade_));
    CascadeMux I__2247 (
            .O(N__13424),
            .I(N__13420));
    CascadeMux I__2246 (
            .O(N__13423),
            .I(N__13417));
    InMux I__2245 (
            .O(N__13420),
            .I(N__13414));
    InMux I__2244 (
            .O(N__13417),
            .I(N__13411));
    LocalMux I__2243 (
            .O(N__13414),
            .I(N__13408));
    LocalMux I__2242 (
            .O(N__13411),
            .I(N__13405));
    Span4Mux_h I__2241 (
            .O(N__13408),
            .I(N__13402));
    Span4Mux_h I__2240 (
            .O(N__13405),
            .I(N__13399));
    Odrv4 I__2239 (
            .O(N__13402),
            .I(\this_vga_signals.N_188_0_0_0 ));
    Odrv4 I__2238 (
            .O(N__13399),
            .I(\this_vga_signals.N_188_0_0_0 ));
    InMux I__2237 (
            .O(N__13394),
            .I(N__13391));
    LocalMux I__2236 (
            .O(N__13391),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_1_0_3 ));
    CascadeMux I__2235 (
            .O(N__13388),
            .I(\this_vga_signals.N_188_0_0_0_cascade_ ));
    CascadeMux I__2234 (
            .O(N__13385),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_1_0_2_cascade_ ));
    CascadeMux I__2233 (
            .O(N__13382),
            .I(N__13379));
    InMux I__2232 (
            .O(N__13379),
            .I(N__13376));
    LocalMux I__2231 (
            .O(N__13376),
            .I(N__13373));
    Odrv12 I__2230 (
            .O(N__13373),
            .I(\this_vga_signals.g1_0_1 ));
    CascadeMux I__2229 (
            .O(N__13370),
            .I(N__13366));
    InMux I__2228 (
            .O(N__13369),
            .I(N__13363));
    InMux I__2227 (
            .O(N__13366),
            .I(N__13360));
    LocalMux I__2226 (
            .O(N__13363),
            .I(N__13355));
    LocalMux I__2225 (
            .O(N__13360),
            .I(N__13351));
    CascadeMux I__2224 (
            .O(N__13359),
            .I(N__13348));
    CascadeMux I__2223 (
            .O(N__13358),
            .I(N__13345));
    Span4Mux_v I__2222 (
            .O(N__13355),
            .I(N__13342));
    InMux I__2221 (
            .O(N__13354),
            .I(N__13339));
    Span4Mux_h I__2220 (
            .O(N__13351),
            .I(N__13336));
    InMux I__2219 (
            .O(N__13348),
            .I(N__13331));
    InMux I__2218 (
            .O(N__13345),
            .I(N__13331));
    Odrv4 I__2217 (
            .O(N__13342),
            .I(N_183_0));
    LocalMux I__2216 (
            .O(N__13339),
            .I(N_183_0));
    Odrv4 I__2215 (
            .O(N__13336),
            .I(N_183_0));
    LocalMux I__2214 (
            .O(N__13331),
            .I(N_183_0));
    CascadeMux I__2213 (
            .O(N__13322),
            .I(N__13318));
    InMux I__2212 (
            .O(N__13321),
            .I(N__13311));
    InMux I__2211 (
            .O(N__13318),
            .I(N__13307));
    InMux I__2210 (
            .O(N__13317),
            .I(N__13304));
    CascadeMux I__2209 (
            .O(N__13316),
            .I(N__13301));
    InMux I__2208 (
            .O(N__13315),
            .I(N__13298));
    CascadeMux I__2207 (
            .O(N__13314),
            .I(N__13294));
    LocalMux I__2206 (
            .O(N__13311),
            .I(N__13289));
    InMux I__2205 (
            .O(N__13310),
            .I(N__13286));
    LocalMux I__2204 (
            .O(N__13307),
            .I(N__13281));
    LocalMux I__2203 (
            .O(N__13304),
            .I(N__13281));
    InMux I__2202 (
            .O(N__13301),
            .I(N__13278));
    LocalMux I__2201 (
            .O(N__13298),
            .I(N__13275));
    CascadeMux I__2200 (
            .O(N__13297),
            .I(N__13272));
    InMux I__2199 (
            .O(N__13294),
            .I(N__13268));
    InMux I__2198 (
            .O(N__13293),
            .I(N__13265));
    InMux I__2197 (
            .O(N__13292),
            .I(N__13262));
    Span4Mux_h I__2196 (
            .O(N__13289),
            .I(N__13259));
    LocalMux I__2195 (
            .O(N__13286),
            .I(N__13250));
    Span4Mux_h I__2194 (
            .O(N__13281),
            .I(N__13250));
    LocalMux I__2193 (
            .O(N__13278),
            .I(N__13250));
    Span4Mux_h I__2192 (
            .O(N__13275),
            .I(N__13250));
    InMux I__2191 (
            .O(N__13272),
            .I(N__13245));
    InMux I__2190 (
            .O(N__13271),
            .I(N__13245));
    LocalMux I__2189 (
            .O(N__13268),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__2188 (
            .O(N__13265),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__2187 (
            .O(N__13262),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__2186 (
            .O(N__13259),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__2185 (
            .O(N__13250),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__2184 (
            .O(N__13245),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    InMux I__2183 (
            .O(N__13232),
            .I(N__13229));
    LocalMux I__2182 (
            .O(N__13229),
            .I(\this_vga_signals.mult1_un40_sum_0_axb1_i ));
    InMux I__2181 (
            .O(N__13226),
            .I(N__13223));
    LocalMux I__2180 (
            .O(N__13223),
            .I(\this_vga_signals.mult1_un40_sum_1_axb1 ));
    CascadeMux I__2179 (
            .O(N__13220),
            .I(\this_vga_signals.mult1_un40_sum_m_x0_1_cascade_ ));
    InMux I__2178 (
            .O(N__13217),
            .I(N__13214));
    LocalMux I__2177 (
            .O(N__13214),
            .I(\this_vga_signals.mult1_un40_sum_m_x1_1 ));
    InMux I__2176 (
            .O(N__13211),
            .I(N__13208));
    LocalMux I__2175 (
            .O(N__13208),
            .I(N__13203));
    InMux I__2174 (
            .O(N__13207),
            .I(N__13200));
    InMux I__2173 (
            .O(N__13206),
            .I(N__13197));
    Odrv4 I__2172 (
            .O(N__13203),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_1 ));
    LocalMux I__2171 (
            .O(N__13200),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_1 ));
    LocalMux I__2170 (
            .O(N__13197),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_1 ));
    CascadeMux I__2169 (
            .O(N__13190),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_1_cascade_ ));
    InMux I__2168 (
            .O(N__13187),
            .I(N__13184));
    LocalMux I__2167 (
            .O(N__13184),
            .I(N__13181));
    Odrv4 I__2166 (
            .O(N__13181),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1 ));
    InMux I__2165 (
            .O(N__13178),
            .I(N__13175));
    LocalMux I__2164 (
            .O(N__13175),
            .I(N__13170));
    InMux I__2163 (
            .O(N__13174),
            .I(N__13165));
    InMux I__2162 (
            .O(N__13173),
            .I(N__13165));
    Odrv4 I__2161 (
            .O(N__13170),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    LocalMux I__2160 (
            .O(N__13165),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    InMux I__2159 (
            .O(N__13160),
            .I(N__13156));
    InMux I__2158 (
            .O(N__13159),
            .I(N__13150));
    LocalMux I__2157 (
            .O(N__13156),
            .I(N__13147));
    CascadeMux I__2156 (
            .O(N__13155),
            .I(N__13142));
    CascadeMux I__2155 (
            .O(N__13154),
            .I(N__13139));
    CascadeMux I__2154 (
            .O(N__13153),
            .I(N__13136));
    LocalMux I__2153 (
            .O(N__13150),
            .I(N__13131));
    Span4Mux_v I__2152 (
            .O(N__13147),
            .I(N__13131));
    InMux I__2151 (
            .O(N__13146),
            .I(N__13128));
    InMux I__2150 (
            .O(N__13145),
            .I(N__13119));
    InMux I__2149 (
            .O(N__13142),
            .I(N__13119));
    InMux I__2148 (
            .O(N__13139),
            .I(N__13119));
    InMux I__2147 (
            .O(N__13136),
            .I(N__13119));
    Odrv4 I__2146 (
            .O(N__13131),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__2145 (
            .O(N__13128),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__2144 (
            .O(N__13119),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    InMux I__2143 (
            .O(N__13112),
            .I(N__13108));
    InMux I__2142 (
            .O(N__13111),
            .I(N__13104));
    LocalMux I__2141 (
            .O(N__13108),
            .I(N__13101));
    InMux I__2140 (
            .O(N__13107),
            .I(N__13098));
    LocalMux I__2139 (
            .O(N__13104),
            .I(N__13095));
    Span4Mux_h I__2138 (
            .O(N__13101),
            .I(N__13092));
    LocalMux I__2137 (
            .O(N__13098),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    Odrv4 I__2136 (
            .O(N__13095),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    Odrv4 I__2135 (
            .O(N__13092),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__2134 (
            .O(N__13085),
            .I(N__13082));
    LocalMux I__2133 (
            .O(N__13082),
            .I(N__13077));
    InMux I__2132 (
            .O(N__13081),
            .I(N__13072));
    InMux I__2131 (
            .O(N__13080),
            .I(N__13072));
    Odrv12 I__2130 (
            .O(N__13077),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__2129 (
            .O(N__13072),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    InMux I__2128 (
            .O(N__13067),
            .I(N__13060));
    InMux I__2127 (
            .O(N__13066),
            .I(N__13060));
    InMux I__2126 (
            .O(N__13065),
            .I(N__13057));
    LocalMux I__2125 (
            .O(N__13060),
            .I(N__13054));
    LocalMux I__2124 (
            .O(N__13057),
            .I(\this_vga_signals.vaddress_7 ));
    Odrv4 I__2123 (
            .O(N__13054),
            .I(\this_vga_signals.vaddress_7 ));
    InMux I__2122 (
            .O(N__13049),
            .I(N__13046));
    LocalMux I__2121 (
            .O(N__13046),
            .I(N__13042));
    InMux I__2120 (
            .O(N__13045),
            .I(N__13039));
    Span4Mux_v I__2119 (
            .O(N__13042),
            .I(N__13035));
    LocalMux I__2118 (
            .O(N__13039),
            .I(N__13032));
    InMux I__2117 (
            .O(N__13038),
            .I(N__13029));
    Odrv4 I__2116 (
            .O(N__13035),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    Odrv12 I__2115 (
            .O(N__13032),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    LocalMux I__2114 (
            .O(N__13029),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__2113 (
            .O(N__13022),
            .I(N__13011));
    InMux I__2112 (
            .O(N__13021),
            .I(N__13011));
    InMux I__2111 (
            .O(N__13020),
            .I(N__13000));
    InMux I__2110 (
            .O(N__13019),
            .I(N__13000));
    InMux I__2109 (
            .O(N__13018),
            .I(N__13000));
    InMux I__2108 (
            .O(N__13017),
            .I(N__13000));
    InMux I__2107 (
            .O(N__13016),
            .I(N__13000));
    LocalMux I__2106 (
            .O(N__13011),
            .I(N__12994));
    LocalMux I__2105 (
            .O(N__13000),
            .I(N__12994));
    InMux I__2104 (
            .O(N__12999),
            .I(N__12988));
    Span4Mux_h I__2103 (
            .O(N__12994),
            .I(N__12985));
    InMux I__2102 (
            .O(N__12993),
            .I(N__12982));
    InMux I__2101 (
            .O(N__12992),
            .I(N__12977));
    InMux I__2100 (
            .O(N__12991),
            .I(N__12977));
    LocalMux I__2099 (
            .O(N__12988),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__2098 (
            .O(N__12985),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__2097 (
            .O(N__12982),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__2096 (
            .O(N__12977),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    InMux I__2095 (
            .O(N__12968),
            .I(N__12962));
    InMux I__2094 (
            .O(N__12967),
            .I(N__12962));
    LocalMux I__2093 (
            .O(N__12962),
            .I(N__12958));
    InMux I__2092 (
            .O(N__12961),
            .I(N__12955));
    Span4Mux_h I__2091 (
            .O(N__12958),
            .I(N__12952));
    LocalMux I__2090 (
            .O(N__12955),
            .I(\this_vga_signals.vaddress_6 ));
    Odrv4 I__2089 (
            .O(N__12952),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__2088 (
            .O(N__12947),
            .I(N__12944));
    LocalMux I__2087 (
            .O(N__12944),
            .I(N__12939));
    InMux I__2086 (
            .O(N__12943),
            .I(N__12936));
    InMux I__2085 (
            .O(N__12942),
            .I(N__12933));
    Span4Mux_h I__2084 (
            .O(N__12939),
            .I(N__12930));
    LocalMux I__2083 (
            .O(N__12936),
            .I(N__12925));
    LocalMux I__2082 (
            .O(N__12933),
            .I(N__12925));
    Span4Mux_v I__2081 (
            .O(N__12930),
            .I(N__12922));
    Span4Mux_v I__2080 (
            .O(N__12925),
            .I(N__12919));
    Odrv4 I__2079 (
            .O(N__12922),
            .I(\this_vga_signals.N_188_0 ));
    Odrv4 I__2078 (
            .O(N__12919),
            .I(\this_vga_signals.N_188_0 ));
    InMux I__2077 (
            .O(N__12914),
            .I(N__12911));
    LocalMux I__2076 (
            .O(N__12911),
            .I(N__12908));
    Odrv4 I__2075 (
            .O(N__12908),
            .I(\this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0 ));
    CascadeMux I__2074 (
            .O(N__12905),
            .I(\this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0_cascade_ ));
    InMux I__2073 (
            .O(N__12902),
            .I(N__12898));
    InMux I__2072 (
            .O(N__12901),
            .I(N__12895));
    LocalMux I__2071 (
            .O(N__12898),
            .I(\this_vga_signals.g1_4 ));
    LocalMux I__2070 (
            .O(N__12895),
            .I(\this_vga_signals.g1_4 ));
    CascadeMux I__2069 (
            .O(N__12890),
            .I(N__12887));
    InMux I__2068 (
            .O(N__12887),
            .I(N__12881));
    InMux I__2067 (
            .O(N__12886),
            .I(N__12881));
    LocalMux I__2066 (
            .O(N__12881),
            .I(N__12878));
    Span4Mux_v I__2065 (
            .O(N__12878),
            .I(N__12874));
    InMux I__2064 (
            .O(N__12877),
            .I(N__12871));
    Odrv4 I__2063 (
            .O(N__12874),
            .I(\this_vga_signals.mult1_un61_sum_s_3 ));
    LocalMux I__2062 (
            .O(N__12871),
            .I(\this_vga_signals.mult1_un61_sum_s_3 ));
    CascadeMux I__2061 (
            .O(N__12866),
            .I(N__12863));
    InMux I__2060 (
            .O(N__12863),
            .I(N__12860));
    LocalMux I__2059 (
            .O(N__12860),
            .I(\this_vga_signals.mult1_un61_sum_i_3 ));
    InMux I__2058 (
            .O(N__12857),
            .I(N__12853));
    InMux I__2057 (
            .O(N__12856),
            .I(N__12848));
    LocalMux I__2056 (
            .O(N__12853),
            .I(N__12845));
    InMux I__2055 (
            .O(N__12852),
            .I(N__12840));
    InMux I__2054 (
            .O(N__12851),
            .I(N__12840));
    LocalMux I__2053 (
            .O(N__12848),
            .I(\this_vga_signals.if_N_3_mux ));
    Odrv4 I__2052 (
            .O(N__12845),
            .I(\this_vga_signals.if_N_3_mux ));
    LocalMux I__2051 (
            .O(N__12840),
            .I(\this_vga_signals.if_N_3_mux ));
    InMux I__2050 (
            .O(N__12833),
            .I(N__12830));
    LocalMux I__2049 (
            .O(N__12830),
            .I(N__12826));
    InMux I__2048 (
            .O(N__12829),
            .I(N__12823));
    Odrv4 I__2047 (
            .O(N__12826),
            .I(\this_vga_signals.g6_0 ));
    LocalMux I__2046 (
            .O(N__12823),
            .I(\this_vga_signals.g6_0 ));
    InMux I__2045 (
            .O(N__12818),
            .I(N__12812));
    InMux I__2044 (
            .O(N__12817),
            .I(N__12809));
    CascadeMux I__2043 (
            .O(N__12816),
            .I(N__12801));
    CascadeMux I__2042 (
            .O(N__12815),
            .I(N__12798));
    LocalMux I__2041 (
            .O(N__12812),
            .I(N__12795));
    LocalMux I__2040 (
            .O(N__12809),
            .I(N__12792));
    InMux I__2039 (
            .O(N__12808),
            .I(N__12789));
    InMux I__2038 (
            .O(N__12807),
            .I(N__12786));
    InMux I__2037 (
            .O(N__12806),
            .I(N__12783));
    InMux I__2036 (
            .O(N__12805),
            .I(N__12774));
    InMux I__2035 (
            .O(N__12804),
            .I(N__12774));
    InMux I__2034 (
            .O(N__12801),
            .I(N__12774));
    InMux I__2033 (
            .O(N__12798),
            .I(N__12774));
    Odrv4 I__2032 (
            .O(N__12795),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__2031 (
            .O(N__12792),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2030 (
            .O(N__12789),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2029 (
            .O(N__12786),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2028 (
            .O(N__12783),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__2027 (
            .O(N__12774),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__2026 (
            .O(N__12761),
            .I(N__12758));
    InMux I__2025 (
            .O(N__12758),
            .I(N__12755));
    LocalMux I__2024 (
            .O(N__12755),
            .I(N__12752));
    Span4Mux_h I__2023 (
            .O(N__12752),
            .I(N__12749));
    Span4Mux_v I__2022 (
            .O(N__12749),
            .I(N__12746));
    Odrv4 I__2021 (
            .O(N__12746),
            .I(M_this_vga_signals_address_13));
    CascadeMux I__2020 (
            .O(N__12743),
            .I(N__12740));
    InMux I__2019 (
            .O(N__12740),
            .I(N__12737));
    LocalMux I__2018 (
            .O(N__12737),
            .I(N__12734));
    Odrv4 I__2017 (
            .O(N__12734),
            .I(\this_vga_signals.g0_0 ));
    InMux I__2016 (
            .O(N__12731),
            .I(N__12728));
    LocalMux I__2015 (
            .O(N__12728),
            .I(\this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0ASZ0 ));
    InMux I__2014 (
            .O(N__12725),
            .I(N__12720));
    InMux I__2013 (
            .O(N__12724),
            .I(N__12717));
    CascadeMux I__2012 (
            .O(N__12723),
            .I(N__12714));
    LocalMux I__2011 (
            .O(N__12720),
            .I(N__12710));
    LocalMux I__2010 (
            .O(N__12717),
            .I(N__12707));
    InMux I__2009 (
            .O(N__12714),
            .I(N__12699));
    InMux I__2008 (
            .O(N__12713),
            .I(N__12699));
    Span4Mux_h I__2007 (
            .O(N__12710),
            .I(N__12694));
    Span4Mux_h I__2006 (
            .O(N__12707),
            .I(N__12694));
    InMux I__2005 (
            .O(N__12706),
            .I(N__12687));
    InMux I__2004 (
            .O(N__12705),
            .I(N__12687));
    InMux I__2003 (
            .O(N__12704),
            .I(N__12687));
    LocalMux I__2002 (
            .O(N__12699),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    Odrv4 I__2001 (
            .O(N__12694),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__2000 (
            .O(N__12687),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    InMux I__1999 (
            .O(N__12680),
            .I(N__12674));
    InMux I__1998 (
            .O(N__12679),
            .I(N__12674));
    LocalMux I__1997 (
            .O(N__12674),
            .I(N__12670));
    InMux I__1996 (
            .O(N__12673),
            .I(N__12667));
    Odrv4 I__1995 (
            .O(N__12670),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__1994 (
            .O(N__12667),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__1993 (
            .O(N__12662),
            .I(N__12657));
    InMux I__1992 (
            .O(N__12661),
            .I(N__12652));
    InMux I__1991 (
            .O(N__12660),
            .I(N__12652));
    LocalMux I__1990 (
            .O(N__12657),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1989 (
            .O(N__12652),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    CascadeMux I__1988 (
            .O(N__12647),
            .I(\this_vga_signals.g0_10_1_cascade_ ));
    InMux I__1987 (
            .O(N__12644),
            .I(N__12641));
    LocalMux I__1986 (
            .O(N__12641),
            .I(N__12636));
    InMux I__1985 (
            .O(N__12640),
            .I(N__12633));
    InMux I__1984 (
            .O(N__12639),
            .I(N__12625));
    Span4Mux_h I__1983 (
            .O(N__12636),
            .I(N__12621));
    LocalMux I__1982 (
            .O(N__12633),
            .I(N__12618));
    InMux I__1981 (
            .O(N__12632),
            .I(N__12615));
    InMux I__1980 (
            .O(N__12631),
            .I(N__12606));
    InMux I__1979 (
            .O(N__12630),
            .I(N__12606));
    InMux I__1978 (
            .O(N__12629),
            .I(N__12606));
    InMux I__1977 (
            .O(N__12628),
            .I(N__12606));
    LocalMux I__1976 (
            .O(N__12625),
            .I(N__12603));
    InMux I__1975 (
            .O(N__12624),
            .I(N__12600));
    Odrv4 I__1974 (
            .O(N__12621),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    Odrv4 I__1973 (
            .O(N__12618),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    LocalMux I__1972 (
            .O(N__12615),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    LocalMux I__1971 (
            .O(N__12606),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    Odrv4 I__1970 (
            .O(N__12603),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    LocalMux I__1969 (
            .O(N__12600),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1 ));
    InMux I__1968 (
            .O(N__12587),
            .I(N__12584));
    LocalMux I__1967 (
            .O(N__12584),
            .I(N__12581));
    Span4Mux_h I__1966 (
            .O(N__12581),
            .I(N__12578));
    Odrv4 I__1965 (
            .O(N__12578),
            .I(\this_vga_signals.if_N_18_1 ));
    InMux I__1964 (
            .O(N__12575),
            .I(N__12572));
    LocalMux I__1963 (
            .O(N__12572),
            .I(\this_vga_signals.m48_i_x4_0 ));
    InMux I__1962 (
            .O(N__12569),
            .I(N__12562));
    InMux I__1961 (
            .O(N__12568),
            .I(N__12562));
    InMux I__1960 (
            .O(N__12567),
            .I(N__12557));
    LocalMux I__1959 (
            .O(N__12562),
            .I(N__12554));
    InMux I__1958 (
            .O(N__12561),
            .I(N__12545));
    InMux I__1957 (
            .O(N__12560),
            .I(N__12542));
    LocalMux I__1956 (
            .O(N__12557),
            .I(N__12539));
    Span4Mux_v I__1955 (
            .O(N__12554),
            .I(N__12529));
    InMux I__1954 (
            .O(N__12553),
            .I(N__12522));
    InMux I__1953 (
            .O(N__12552),
            .I(N__12522));
    InMux I__1952 (
            .O(N__12551),
            .I(N__12522));
    InMux I__1951 (
            .O(N__12550),
            .I(N__12515));
    InMux I__1950 (
            .O(N__12549),
            .I(N__12515));
    InMux I__1949 (
            .O(N__12548),
            .I(N__12515));
    LocalMux I__1948 (
            .O(N__12545),
            .I(N__12510));
    LocalMux I__1947 (
            .O(N__12542),
            .I(N__12510));
    Span4Mux_h I__1946 (
            .O(N__12539),
            .I(N__12507));
    InMux I__1945 (
            .O(N__12538),
            .I(N__12498));
    InMux I__1944 (
            .O(N__12537),
            .I(N__12498));
    InMux I__1943 (
            .O(N__12536),
            .I(N__12498));
    InMux I__1942 (
            .O(N__12535),
            .I(N__12498));
    InMux I__1941 (
            .O(N__12534),
            .I(N__12491));
    InMux I__1940 (
            .O(N__12533),
            .I(N__12491));
    InMux I__1939 (
            .O(N__12532),
            .I(N__12491));
    Odrv4 I__1938 (
            .O(N__12529),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    LocalMux I__1937 (
            .O(N__12522),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    LocalMux I__1936 (
            .O(N__12515),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    Odrv4 I__1935 (
            .O(N__12510),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    Odrv4 I__1934 (
            .O(N__12507),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    LocalMux I__1933 (
            .O(N__12498),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    LocalMux I__1932 (
            .O(N__12491),
            .I(\this_vga_signals.mult1_un47_sum_c3_0 ));
    CascadeMux I__1931 (
            .O(N__12476),
            .I(N__12473));
    InMux I__1930 (
            .O(N__12473),
            .I(N__12470));
    LocalMux I__1929 (
            .O(N__12470),
            .I(\this_vga_signals.g4_1_0 ));
    InMux I__1928 (
            .O(N__12467),
            .I(N__12461));
    InMux I__1927 (
            .O(N__12466),
            .I(N__12461));
    LocalMux I__1926 (
            .O(N__12461),
            .I(N__12458));
    Span4Mux_h I__1925 (
            .O(N__12458),
            .I(N__12453));
    InMux I__1924 (
            .O(N__12457),
            .I(N__12448));
    InMux I__1923 (
            .O(N__12456),
            .I(N__12448));
    Odrv4 I__1922 (
            .O(N__12453),
            .I(\this_vga_signals.g0_1 ));
    LocalMux I__1921 (
            .O(N__12448),
            .I(\this_vga_signals.g0_1 ));
    InMux I__1920 (
            .O(N__12443),
            .I(\this_vga_signals.mult1_un68_sum_cry_0 ));
    InMux I__1919 (
            .O(N__12440),
            .I(N__12437));
    LocalMux I__1918 (
            .O(N__12437),
            .I(N__12434));
    Span12Mux_h I__1917 (
            .O(N__12434),
            .I(N__12431));
    Odrv12 I__1916 (
            .O(N__12431),
            .I(\this_vga_signals.mult1_un61_sum_cry_1_s ));
    InMux I__1915 (
            .O(N__12428),
            .I(\this_vga_signals.mult1_un68_sum_cry_1 ));
    InMux I__1914 (
            .O(N__12425),
            .I(N__12422));
    LocalMux I__1913 (
            .O(N__12422),
            .I(N__12419));
    Span4Mux_v I__1912 (
            .O(N__12419),
            .I(N__12416));
    Odrv4 I__1911 (
            .O(N__12416),
            .I(\this_vga_signals.mult1_un68_sum_axb_3 ));
    InMux I__1910 (
            .O(N__12413),
            .I(\this_vga_signals.mult1_un68_sum_cry_2 ));
    InMux I__1909 (
            .O(N__12410),
            .I(N__12407));
    LocalMux I__1908 (
            .O(N__12407),
            .I(N__12401));
    InMux I__1907 (
            .O(N__12406),
            .I(N__12398));
    InMux I__1906 (
            .O(N__12405),
            .I(N__12395));
    InMux I__1905 (
            .O(N__12404),
            .I(N__12392));
    Odrv4 I__1904 (
            .O(N__12401),
            .I(\this_vga_signals.vaddress_8 ));
    LocalMux I__1903 (
            .O(N__12398),
            .I(\this_vga_signals.vaddress_8 ));
    LocalMux I__1902 (
            .O(N__12395),
            .I(\this_vga_signals.vaddress_8 ));
    LocalMux I__1901 (
            .O(N__12392),
            .I(\this_vga_signals.vaddress_8 ));
    InMux I__1900 (
            .O(N__12383),
            .I(N__12380));
    LocalMux I__1899 (
            .O(N__12380),
            .I(\this_vga_signals.N_3_2 ));
    InMux I__1898 (
            .O(N__12377),
            .I(N__12369));
    CascadeMux I__1897 (
            .O(N__12376),
            .I(N__12358));
    InMux I__1896 (
            .O(N__12375),
            .I(N__12348));
    InMux I__1895 (
            .O(N__12374),
            .I(N__12348));
    InMux I__1894 (
            .O(N__12373),
            .I(N__12348));
    InMux I__1893 (
            .O(N__12372),
            .I(N__12348));
    LocalMux I__1892 (
            .O(N__12369),
            .I(N__12345));
    InMux I__1891 (
            .O(N__12368),
            .I(N__12340));
    InMux I__1890 (
            .O(N__12367),
            .I(N__12340));
    InMux I__1889 (
            .O(N__12366),
            .I(N__12337));
    InMux I__1888 (
            .O(N__12365),
            .I(N__12330));
    InMux I__1887 (
            .O(N__12364),
            .I(N__12330));
    InMux I__1886 (
            .O(N__12363),
            .I(N__12330));
    InMux I__1885 (
            .O(N__12362),
            .I(N__12323));
    InMux I__1884 (
            .O(N__12361),
            .I(N__12323));
    InMux I__1883 (
            .O(N__12358),
            .I(N__12323));
    InMux I__1882 (
            .O(N__12357),
            .I(N__12320));
    LocalMux I__1881 (
            .O(N__12348),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    Odrv4 I__1880 (
            .O(N__12345),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__1879 (
            .O(N__12340),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__1878 (
            .O(N__12337),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__1877 (
            .O(N__12330),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__1876 (
            .O(N__12323),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    LocalMux I__1875 (
            .O(N__12320),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ));
    InMux I__1874 (
            .O(N__12305),
            .I(N__12302));
    LocalMux I__1873 (
            .O(N__12302),
            .I(\this_vga_signals.g0_16_x1 ));
    InMux I__1872 (
            .O(N__12299),
            .I(N__12295));
    InMux I__1871 (
            .O(N__12298),
            .I(N__12292));
    LocalMux I__1870 (
            .O(N__12295),
            .I(\this_vga_signals.N_81_1 ));
    LocalMux I__1869 (
            .O(N__12292),
            .I(\this_vga_signals.N_81_1 ));
    InMux I__1868 (
            .O(N__12287),
            .I(N__12284));
    LocalMux I__1867 (
            .O(N__12284),
            .I(\this_vga_signals.g1_2 ));
    InMux I__1866 (
            .O(N__12281),
            .I(N__12277));
    InMux I__1865 (
            .O(N__12280),
            .I(N__12274));
    LocalMux I__1864 (
            .O(N__12277),
            .I(\this_vga_signals.if_N_7_i ));
    LocalMux I__1863 (
            .O(N__12274),
            .I(\this_vga_signals.if_N_7_i ));
    InMux I__1862 (
            .O(N__12269),
            .I(N__12265));
    InMux I__1861 (
            .O(N__12268),
            .I(N__12262));
    LocalMux I__1860 (
            .O(N__12265),
            .I(\this_vga_signals.if_N_11 ));
    LocalMux I__1859 (
            .O(N__12262),
            .I(\this_vga_signals.if_N_11 ));
    CascadeMux I__1858 (
            .O(N__12257),
            .I(\this_vga_signals.if_i3_mux_0_1_cascade_ ));
    InMux I__1857 (
            .O(N__12254),
            .I(N__12251));
    LocalMux I__1856 (
            .O(N__12251),
            .I(\this_vga_signals.m48_i_x4_3 ));
    CascadeMux I__1855 (
            .O(N__12248),
            .I(N__12245));
    InMux I__1854 (
            .O(N__12245),
            .I(N__12242));
    LocalMux I__1853 (
            .O(N__12242),
            .I(N__12239));
    Odrv4 I__1852 (
            .O(N__12239),
            .I(\this_vga_signals.if_i3_mux_0_1 ));
    InMux I__1851 (
            .O(N__12236),
            .I(N__12230));
    InMux I__1850 (
            .O(N__12235),
            .I(N__12230));
    LocalMux I__1849 (
            .O(N__12230),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0_0 ));
    InMux I__1848 (
            .O(N__12227),
            .I(N__12224));
    LocalMux I__1847 (
            .O(N__12224),
            .I(\this_vga_signals.N_57_0 ));
    InMux I__1846 (
            .O(N__12221),
            .I(N__12218));
    LocalMux I__1845 (
            .O(N__12218),
            .I(\this_vga_signals.N_57_i_i_0 ));
    CascadeMux I__1844 (
            .O(N__12215),
            .I(\this_vga_signals.g1_0_cascade_ ));
    InMux I__1843 (
            .O(N__12212),
            .I(N__12209));
    LocalMux I__1842 (
            .O(N__12209),
            .I(\this_vga_signals.if_N_6_mux_0_0_0 ));
    InMux I__1841 (
            .O(N__12206),
            .I(N__12203));
    LocalMux I__1840 (
            .O(N__12203),
            .I(\this_vga_signals.g2_1_0_0 ));
    InMux I__1839 (
            .O(N__12200),
            .I(N__12195));
    InMux I__1838 (
            .O(N__12199),
            .I(N__12184));
    InMux I__1837 (
            .O(N__12198),
            .I(N__12184));
    LocalMux I__1836 (
            .O(N__12195),
            .I(N__12181));
    InMux I__1835 (
            .O(N__12194),
            .I(N__12176));
    InMux I__1834 (
            .O(N__12193),
            .I(N__12176));
    CascadeMux I__1833 (
            .O(N__12192),
            .I(N__12161));
    InMux I__1832 (
            .O(N__12191),
            .I(N__12156));
    InMux I__1831 (
            .O(N__12190),
            .I(N__12156));
    InMux I__1830 (
            .O(N__12189),
            .I(N__12153));
    LocalMux I__1829 (
            .O(N__12184),
            .I(N__12150));
    Span4Mux_v I__1828 (
            .O(N__12181),
            .I(N__12145));
    LocalMux I__1827 (
            .O(N__12176),
            .I(N__12145));
    InMux I__1826 (
            .O(N__12175),
            .I(N__12140));
    InMux I__1825 (
            .O(N__12174),
            .I(N__12140));
    InMux I__1824 (
            .O(N__12173),
            .I(N__12137));
    InMux I__1823 (
            .O(N__12172),
            .I(N__12126));
    InMux I__1822 (
            .O(N__12171),
            .I(N__12126));
    InMux I__1821 (
            .O(N__12170),
            .I(N__12126));
    InMux I__1820 (
            .O(N__12169),
            .I(N__12126));
    InMux I__1819 (
            .O(N__12168),
            .I(N__12126));
    InMux I__1818 (
            .O(N__12167),
            .I(N__12117));
    InMux I__1817 (
            .O(N__12166),
            .I(N__12117));
    InMux I__1816 (
            .O(N__12165),
            .I(N__12117));
    InMux I__1815 (
            .O(N__12164),
            .I(N__12117));
    InMux I__1814 (
            .O(N__12161),
            .I(N__12114));
    LocalMux I__1813 (
            .O(N__12156),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1812 (
            .O(N__12153),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__1811 (
            .O(N__12150),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__1810 (
            .O(N__12145),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1809 (
            .O(N__12140),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1808 (
            .O(N__12137),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1807 (
            .O(N__12126),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1806 (
            .O(N__12117),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1805 (
            .O(N__12114),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    InMux I__1804 (
            .O(N__12095),
            .I(N__12092));
    LocalMux I__1803 (
            .O(N__12092),
            .I(N__12085));
    InMux I__1802 (
            .O(N__12091),
            .I(N__12079));
    InMux I__1801 (
            .O(N__12090),
            .I(N__12074));
    InMux I__1800 (
            .O(N__12089),
            .I(N__12074));
    CascadeMux I__1799 (
            .O(N__12088),
            .I(N__12062));
    Span4Mux_v I__1798 (
            .O(N__12085),
            .I(N__12058));
    InMux I__1797 (
            .O(N__12084),
            .I(N__12053));
    InMux I__1796 (
            .O(N__12083),
            .I(N__12053));
    InMux I__1795 (
            .O(N__12082),
            .I(N__12050));
    LocalMux I__1794 (
            .O(N__12079),
            .I(N__12047));
    LocalMux I__1793 (
            .O(N__12074),
            .I(N__12044));
    InMux I__1792 (
            .O(N__12073),
            .I(N__12041));
    InMux I__1791 (
            .O(N__12072),
            .I(N__12036));
    InMux I__1790 (
            .O(N__12071),
            .I(N__12036));
    InMux I__1789 (
            .O(N__12070),
            .I(N__12029));
    InMux I__1788 (
            .O(N__12069),
            .I(N__12029));
    InMux I__1787 (
            .O(N__12068),
            .I(N__12029));
    InMux I__1786 (
            .O(N__12067),
            .I(N__12020));
    InMux I__1785 (
            .O(N__12066),
            .I(N__12020));
    InMux I__1784 (
            .O(N__12065),
            .I(N__12020));
    InMux I__1783 (
            .O(N__12062),
            .I(N__12020));
    InMux I__1782 (
            .O(N__12061),
            .I(N__12017));
    Odrv4 I__1781 (
            .O(N__12058),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1780 (
            .O(N__12053),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1779 (
            .O(N__12050),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    Odrv4 I__1778 (
            .O(N__12047),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    Odrv4 I__1777 (
            .O(N__12044),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1776 (
            .O(N__12041),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1775 (
            .O(N__12036),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1774 (
            .O(N__12029),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1773 (
            .O(N__12020),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1772 (
            .O(N__12017),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    InMux I__1771 (
            .O(N__11996),
            .I(N__11992));
    CascadeMux I__1770 (
            .O(N__11995),
            .I(N__11989));
    LocalMux I__1769 (
            .O(N__11992),
            .I(N__11986));
    InMux I__1768 (
            .O(N__11989),
            .I(N__11983));
    Odrv4 I__1767 (
            .O(N__11986),
            .I(\this_vga_signals.N_5_i_1_0 ));
    LocalMux I__1766 (
            .O(N__11983),
            .I(\this_vga_signals.N_5_i_1_0 ));
    CascadeMux I__1765 (
            .O(N__11978),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_1_0_x1_cascade_ ));
    InMux I__1764 (
            .O(N__11975),
            .I(N__11972));
    LocalMux I__1763 (
            .O(N__11972),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_1_0 ));
    InMux I__1762 (
            .O(N__11969),
            .I(N__11966));
    LocalMux I__1761 (
            .O(N__11966),
            .I(\this_vga_signals.mult1_un61_sum_ac0_2_2_1 ));
    CascadeMux I__1760 (
            .O(N__11963),
            .I(\this_vga_signals.mult1_un61_sum_ac0_2_2_1_cascade_ ));
    InMux I__1759 (
            .O(N__11960),
            .I(N__11957));
    LocalMux I__1758 (
            .O(N__11957),
            .I(N__11950));
    InMux I__1757 (
            .O(N__11956),
            .I(N__11943));
    InMux I__1756 (
            .O(N__11955),
            .I(N__11943));
    InMux I__1755 (
            .O(N__11954),
            .I(N__11943));
    InMux I__1754 (
            .O(N__11953),
            .I(N__11940));
    Odrv4 I__1753 (
            .O(N__11950),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0));
    LocalMux I__1752 (
            .O(N__11943),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0));
    LocalMux I__1751 (
            .O(N__11940),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0));
    InMux I__1750 (
            .O(N__11933),
            .I(N__11930));
    LocalMux I__1749 (
            .O(N__11930),
            .I(N__11926));
    InMux I__1748 (
            .O(N__11929),
            .I(N__11923));
    Odrv4 I__1747 (
            .O(N__11926),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    LocalMux I__1746 (
            .O(N__11923),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    InMux I__1745 (
            .O(N__11918),
            .I(N__11909));
    InMux I__1744 (
            .O(N__11917),
            .I(N__11909));
    InMux I__1743 (
            .O(N__11916),
            .I(N__11909));
    LocalMux I__1742 (
            .O(N__11909),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_2 ));
    InMux I__1741 (
            .O(N__11906),
            .I(N__11903));
    LocalMux I__1740 (
            .O(N__11903),
            .I(\this_vga_signals.mult1_un61_sum_ac0_sx ));
    InMux I__1739 (
            .O(N__11900),
            .I(N__11896));
    InMux I__1738 (
            .O(N__11899),
            .I(N__11893));
    LocalMux I__1737 (
            .O(N__11896),
            .I(\this_vga_signals.mult1_un61_sum_ac0_2_4_tz ));
    LocalMux I__1736 (
            .O(N__11893),
            .I(\this_vga_signals.mult1_un61_sum_ac0_2_4_tz ));
    InMux I__1735 (
            .O(N__11888),
            .I(N__11884));
    InMux I__1734 (
            .O(N__11887),
            .I(N__11881));
    LocalMux I__1733 (
            .O(N__11884),
            .I(N__11874));
    LocalMux I__1732 (
            .O(N__11881),
            .I(N__11874));
    InMux I__1731 (
            .O(N__11880),
            .I(N__11871));
    InMux I__1730 (
            .O(N__11879),
            .I(N__11868));
    Odrv4 I__1729 (
            .O(N__11874),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    LocalMux I__1728 (
            .O(N__11871),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    LocalMux I__1727 (
            .O(N__11868),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_3 ));
    CascadeMux I__1726 (
            .O(N__11861),
            .I(\this_vga_signals.mult1_un61_sum_ac0_2_cascade_ ));
    InMux I__1725 (
            .O(N__11858),
            .I(N__11854));
    CascadeMux I__1724 (
            .O(N__11857),
            .I(N__11850));
    LocalMux I__1723 (
            .O(N__11854),
            .I(N__11845));
    InMux I__1722 (
            .O(N__11853),
            .I(N__11841));
    InMux I__1721 (
            .O(N__11850),
            .I(N__11836));
    InMux I__1720 (
            .O(N__11849),
            .I(N__11836));
    InMux I__1719 (
            .O(N__11848),
            .I(N__11832));
    Span4Mux_v I__1718 (
            .O(N__11845),
            .I(N__11826));
    InMux I__1717 (
            .O(N__11844),
            .I(N__11823));
    LocalMux I__1716 (
            .O(N__11841),
            .I(N__11820));
    LocalMux I__1715 (
            .O(N__11836),
            .I(N__11817));
    InMux I__1714 (
            .O(N__11835),
            .I(N__11814));
    LocalMux I__1713 (
            .O(N__11832),
            .I(N__11811));
    InMux I__1712 (
            .O(N__11831),
            .I(N__11806));
    InMux I__1711 (
            .O(N__11830),
            .I(N__11806));
    InMux I__1710 (
            .O(N__11829),
            .I(N__11803));
    Odrv4 I__1709 (
            .O(N__11826),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    LocalMux I__1708 (
            .O(N__11823),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    Odrv4 I__1707 (
            .O(N__11820),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    Odrv4 I__1706 (
            .O(N__11817),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    LocalMux I__1705 (
            .O(N__11814),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    Odrv4 I__1704 (
            .O(N__11811),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    LocalMux I__1703 (
            .O(N__11806),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    LocalMux I__1702 (
            .O(N__11803),
            .I(this_vga_signals_un4_lcounter_if_i3_mux));
    InMux I__1701 (
            .O(N__11786),
            .I(N__11783));
    LocalMux I__1700 (
            .O(N__11783),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    InMux I__1699 (
            .O(N__11780),
            .I(N__11777));
    LocalMux I__1698 (
            .O(N__11777),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    InMux I__1697 (
            .O(N__11774),
            .I(N__11771));
    LocalMux I__1696 (
            .O(N__11771),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    InMux I__1695 (
            .O(N__11768),
            .I(N__11764));
    InMux I__1694 (
            .O(N__11767),
            .I(N__11761));
    LocalMux I__1693 (
            .O(N__11764),
            .I(\this_vga_signals.N_81_0 ));
    LocalMux I__1692 (
            .O(N__11761),
            .I(\this_vga_signals.N_81_0 ));
    InMux I__1691 (
            .O(N__11756),
            .I(N__11749));
    InMux I__1690 (
            .O(N__11755),
            .I(N__11749));
    InMux I__1689 (
            .O(N__11754),
            .I(N__11746));
    LocalMux I__1688 (
            .O(N__11749),
            .I(N__11743));
    LocalMux I__1687 (
            .O(N__11746),
            .I(\this_vga_signals.N_370_0 ));
    Odrv4 I__1686 (
            .O(N__11743),
            .I(\this_vga_signals.N_370_0 ));
    InMux I__1685 (
            .O(N__11738),
            .I(N__11735));
    LocalMux I__1684 (
            .O(N__11735),
            .I(\this_vga_signals.mult1_un40_sum1_2 ));
    CascadeMux I__1683 (
            .O(N__11732),
            .I(N__11729));
    InMux I__1682 (
            .O(N__11729),
            .I(N__11716));
    InMux I__1681 (
            .O(N__11728),
            .I(N__11716));
    InMux I__1680 (
            .O(N__11727),
            .I(N__11716));
    InMux I__1679 (
            .O(N__11726),
            .I(N__11716));
    InMux I__1678 (
            .O(N__11725),
            .I(N__11712));
    LocalMux I__1677 (
            .O(N__11716),
            .I(N__11709));
    InMux I__1676 (
            .O(N__11715),
            .I(N__11706));
    LocalMux I__1675 (
            .O(N__11712),
            .I(this_vga_signals_M_vcounter_q_7_rep1));
    Odrv4 I__1674 (
            .O(N__11709),
            .I(this_vga_signals_M_vcounter_q_7_rep1));
    LocalMux I__1673 (
            .O(N__11706),
            .I(this_vga_signals_M_vcounter_q_7_rep1));
    InMux I__1672 (
            .O(N__11699),
            .I(N__11685));
    InMux I__1671 (
            .O(N__11698),
            .I(N__11685));
    InMux I__1670 (
            .O(N__11697),
            .I(N__11685));
    InMux I__1669 (
            .O(N__11696),
            .I(N__11685));
    InMux I__1668 (
            .O(N__11695),
            .I(N__11680));
    InMux I__1667 (
            .O(N__11694),
            .I(N__11680));
    LocalMux I__1666 (
            .O(N__11685),
            .I(this_vga_signals_M_vcounter_q_8_rep1));
    LocalMux I__1665 (
            .O(N__11680),
            .I(this_vga_signals_M_vcounter_q_8_rep1));
    InMux I__1664 (
            .O(N__11675),
            .I(N__11671));
    InMux I__1663 (
            .O(N__11674),
            .I(N__11668));
    LocalMux I__1662 (
            .O(N__11671),
            .I(\this_vga_signals.N_330_0 ));
    LocalMux I__1661 (
            .O(N__11668),
            .I(\this_vga_signals.N_330_0 ));
    CascadeMux I__1660 (
            .O(N__11663),
            .I(N__11660));
    InMux I__1659 (
            .O(N__11660),
            .I(N__11657));
    LocalMux I__1658 (
            .O(N__11657),
            .I(N__11654));
    Span4Mux_v I__1657 (
            .O(N__11654),
            .I(N__11651));
    Odrv4 I__1656 (
            .O(N__11651),
            .I(\this_vga_signals.vsync_1_0_a2_6_a2_0 ));
    CascadeMux I__1655 (
            .O(N__11648),
            .I(\this_vga_signals.if_m11_1_cascade_ ));
    InMux I__1654 (
            .O(N__11645),
            .I(N__11642));
    LocalMux I__1653 (
            .O(N__11642),
            .I(N__11639));
    Span4Mux_h I__1652 (
            .O(N__11639),
            .I(N__11636));
    Odrv4 I__1651 (
            .O(N__11636),
            .I(\this_vga_signals.mult1_un47_sum_i_0 ));
    CascadeMux I__1650 (
            .O(N__11633),
            .I(\this_vga_signals.mult1_un61_sum_ac0_2_2_cascade_ ));
    InMux I__1649 (
            .O(N__11630),
            .I(N__11627));
    LocalMux I__1648 (
            .O(N__11627),
            .I(N__11624));
    Odrv4 I__1647 (
            .O(N__11624),
            .I(\this_vga_signals.mult1_un61_sum_axb2_i ));
    CascadeMux I__1646 (
            .O(N__11621),
            .I(N__11617));
    InMux I__1645 (
            .O(N__11620),
            .I(N__11613));
    InMux I__1644 (
            .O(N__11617),
            .I(N__11610));
    InMux I__1643 (
            .O(N__11616),
            .I(N__11606));
    LocalMux I__1642 (
            .O(N__11613),
            .I(N__11603));
    LocalMux I__1641 (
            .O(N__11610),
            .I(N__11600));
    InMux I__1640 (
            .O(N__11609),
            .I(N__11597));
    LocalMux I__1639 (
            .O(N__11606),
            .I(N__11592));
    Span4Mux_v I__1638 (
            .O(N__11603),
            .I(N__11585));
    Span4Mux_h I__1637 (
            .O(N__11600),
            .I(N__11585));
    LocalMux I__1636 (
            .O(N__11597),
            .I(N__11585));
    InMux I__1635 (
            .O(N__11596),
            .I(N__11580));
    InMux I__1634 (
            .O(N__11595),
            .I(N__11580));
    Odrv4 I__1633 (
            .O(N__11592),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    Odrv4 I__1632 (
            .O(N__11585),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__1631 (
            .O(N__11580),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    CascadeMux I__1630 (
            .O(N__11573),
            .I(N__11570));
    InMux I__1629 (
            .O(N__11570),
            .I(N__11564));
    InMux I__1628 (
            .O(N__11569),
            .I(N__11564));
    LocalMux I__1627 (
            .O(N__11564),
            .I(\this_vga_signals.if_m5_0_1 ));
    CascadeMux I__1626 (
            .O(N__11561),
            .I(N__11558));
    InMux I__1625 (
            .O(N__11558),
            .I(N__11554));
    InMux I__1624 (
            .O(N__11557),
            .I(N__11551));
    LocalMux I__1623 (
            .O(N__11554),
            .I(N__11548));
    LocalMux I__1622 (
            .O(N__11551),
            .I(\this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1 ));
    Odrv4 I__1621 (
            .O(N__11548),
            .I(\this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1 ));
    CascadeMux I__1620 (
            .O(N__11543),
            .I(\this_vga_signals.mult1_un40_sum_0_axb1_i_cascade_ ));
    InMux I__1619 (
            .O(N__11540),
            .I(N__11535));
    InMux I__1618 (
            .O(N__11539),
            .I(N__11530));
    InMux I__1617 (
            .O(N__11538),
            .I(N__11530));
    LocalMux I__1616 (
            .O(N__11535),
            .I(\this_vga_signals.mult1_un47_sum_ac0_1 ));
    LocalMux I__1615 (
            .O(N__11530),
            .I(\this_vga_signals.mult1_un47_sum_ac0_1 ));
    CascadeMux I__1614 (
            .O(N__11525),
            .I(N__11521));
    CascadeMux I__1613 (
            .O(N__11524),
            .I(N__11517));
    InMux I__1612 (
            .O(N__11521),
            .I(N__11512));
    InMux I__1611 (
            .O(N__11520),
            .I(N__11512));
    InMux I__1610 (
            .O(N__11517),
            .I(N__11509));
    LocalMux I__1609 (
            .O(N__11512),
            .I(N__11506));
    LocalMux I__1608 (
            .O(N__11509),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c ));
    Odrv4 I__1607 (
            .O(N__11506),
            .I(\this_vga_signals.mult1_un47_sum_ac0_3_c ));
    CascadeMux I__1606 (
            .O(N__11501),
            .I(N_475_cascade_));
    CascadeMux I__1605 (
            .O(N__11498),
            .I(\this_vga_signals.if_N_3_mux_cascade_ ));
    InMux I__1604 (
            .O(N__11495),
            .I(N__11491));
    InMux I__1603 (
            .O(N__11494),
            .I(N__11488));
    LocalMux I__1602 (
            .O(N__11491),
            .I(N__11483));
    LocalMux I__1601 (
            .O(N__11488),
            .I(N__11483));
    Odrv4 I__1600 (
            .O(N__11483),
            .I(\this_vga_signals.mult1_un47_sum_axb2_0 ));
    InMux I__1599 (
            .O(N__11480),
            .I(N__11477));
    LocalMux I__1598 (
            .O(N__11477),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_x1 ));
    CascadeMux I__1597 (
            .O(N__11474),
            .I(\this_vga_signals.mult1_un47_sum_axb2_0_cascade_ ));
    InMux I__1596 (
            .O(N__11471),
            .I(N__11468));
    LocalMux I__1595 (
            .O(N__11468),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_x0 ));
    InMux I__1594 (
            .O(N__11465),
            .I(N__11459));
    InMux I__1593 (
            .O(N__11464),
            .I(N__11459));
    LocalMux I__1592 (
            .O(N__11459),
            .I(N__11456));
    Odrv4 I__1591 (
            .O(N__11456),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    InMux I__1590 (
            .O(N__11453),
            .I(N__11450));
    LocalMux I__1589 (
            .O(N__11450),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_1_0_x1 ));
    CascadeMux I__1588 (
            .O(N__11447),
            .I(N__11444));
    InMux I__1587 (
            .O(N__11444),
            .I(N__11440));
    CascadeMux I__1586 (
            .O(N__11443),
            .I(N__11436));
    LocalMux I__1585 (
            .O(N__11440),
            .I(N__11432));
    InMux I__1584 (
            .O(N__11439),
            .I(N__11425));
    InMux I__1583 (
            .O(N__11436),
            .I(N__11425));
    InMux I__1582 (
            .O(N__11435),
            .I(N__11425));
    Odrv4 I__1581 (
            .O(N__11432),
            .I(this_vga_signals_M_vcounter_q_fast_6));
    LocalMux I__1580 (
            .O(N__11425),
            .I(this_vga_signals_M_vcounter_q_fast_6));
    InMux I__1579 (
            .O(N__11420),
            .I(N__11417));
    LocalMux I__1578 (
            .O(N__11417),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_1_0_x0 ));
    InMux I__1577 (
            .O(N__11414),
            .I(N__11411));
    LocalMux I__1576 (
            .O(N__11411),
            .I(\this_vga_signals.if_m10_0_a4_1_0_x1 ));
    CascadeMux I__1575 (
            .O(N__11408),
            .I(\this_vga_signals.if_m10_0_a4_1_0_x0_cascade_ ));
    InMux I__1574 (
            .O(N__11405),
            .I(N__11402));
    LocalMux I__1573 (
            .O(N__11402),
            .I(\this_vga_signals.if_m10_0_a4_1 ));
    InMux I__1572 (
            .O(N__11399),
            .I(N__11394));
    InMux I__1571 (
            .O(N__11398),
            .I(N__11391));
    InMux I__1570 (
            .O(N__11397),
            .I(N__11388));
    LocalMux I__1569 (
            .O(N__11394),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__1568 (
            .O(N__11391),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__1567 (
            .O(N__11388),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    InMux I__1566 (
            .O(N__11381),
            .I(N__11375));
    InMux I__1565 (
            .O(N__11380),
            .I(N__11375));
    LocalMux I__1564 (
            .O(N__11375),
            .I(\this_vga_signals.g0_0_a3_0 ));
    CascadeMux I__1563 (
            .O(N__11372),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNISGOSZ0Z_4_cascade_ ));
    CascadeMux I__1562 (
            .O(N__11369),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1_x0_cascade_ ));
    InMux I__1561 (
            .O(N__11366),
            .I(N__11363));
    LocalMux I__1560 (
            .O(N__11363),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1_x1 ));
    CascadeMux I__1559 (
            .O(N__11360),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_1_cascade_ ));
    CascadeMux I__1558 (
            .O(N__11357),
            .I(\this_vga_signals.if_m10_0_x2_0_0_cascade_ ));
    CascadeMux I__1557 (
            .O(N__11354),
            .I(N__11351));
    InMux I__1556 (
            .O(N__11351),
            .I(N__11348));
    LocalMux I__1555 (
            .O(N__11348),
            .I(\this_vga_signals.mult1_un47_sum_c2_0 ));
    CascadeMux I__1554 (
            .O(N__11345),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ));
    CascadeMux I__1553 (
            .O(N__11342),
            .I(\this_vga_signals.mult1_un47_sum_c3_0_cascade_ ));
    InMux I__1552 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1551 (
            .O(N__11336),
            .I(N__11333));
    Odrv4 I__1550 (
            .O(N__11333),
            .I(\this_vga_signals.if_m2_1 ));
    InMux I__1549 (
            .O(N__11330),
            .I(N__11326));
    CascadeMux I__1548 (
            .O(N__11329),
            .I(N__11321));
    LocalMux I__1547 (
            .O(N__11326),
            .I(N__11318));
    CascadeMux I__1546 (
            .O(N__11325),
            .I(N__11315));
    InMux I__1545 (
            .O(N__11324),
            .I(N__11311));
    InMux I__1544 (
            .O(N__11321),
            .I(N__11308));
    Span4Mux_v I__1543 (
            .O(N__11318),
            .I(N__11305));
    InMux I__1542 (
            .O(N__11315),
            .I(N__11300));
    InMux I__1541 (
            .O(N__11314),
            .I(N__11300));
    LocalMux I__1540 (
            .O(N__11311),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__1539 (
            .O(N__11308),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    Odrv4 I__1538 (
            .O(N__11305),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__1537 (
            .O(N__11300),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    CascadeMux I__1536 (
            .O(N__11291),
            .I(\this_vga_signals.g1_2_cascade_ ));
    CascadeMux I__1535 (
            .O(N__11288),
            .I(N__11280));
    InMux I__1534 (
            .O(N__11287),
            .I(N__11266));
    InMux I__1533 (
            .O(N__11286),
            .I(N__11266));
    InMux I__1532 (
            .O(N__11285),
            .I(N__11263));
    InMux I__1531 (
            .O(N__11284),
            .I(N__11258));
    InMux I__1530 (
            .O(N__11283),
            .I(N__11258));
    InMux I__1529 (
            .O(N__11280),
            .I(N__11249));
    InMux I__1528 (
            .O(N__11279),
            .I(N__11249));
    InMux I__1527 (
            .O(N__11278),
            .I(N__11249));
    InMux I__1526 (
            .O(N__11277),
            .I(N__11249));
    InMux I__1525 (
            .O(N__11276),
            .I(N__11244));
    InMux I__1524 (
            .O(N__11275),
            .I(N__11244));
    InMux I__1523 (
            .O(N__11274),
            .I(N__11235));
    InMux I__1522 (
            .O(N__11273),
            .I(N__11235));
    InMux I__1521 (
            .O(N__11272),
            .I(N__11235));
    InMux I__1520 (
            .O(N__11271),
            .I(N__11235));
    LocalMux I__1519 (
            .O(N__11266),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1518 (
            .O(N__11263),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1517 (
            .O(N__11258),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1516 (
            .O(N__11249),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1515 (
            .O(N__11244),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    LocalMux I__1514 (
            .O(N__11235),
            .I(\this_vga_signals.mult1_un61_sum_c3 ));
    CascadeMux I__1513 (
            .O(N__11222),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ));
    InMux I__1512 (
            .O(N__11219),
            .I(N__11216));
    LocalMux I__1511 (
            .O(N__11216),
            .I(\this_vga_signals.g1_1 ));
    InMux I__1510 (
            .O(N__11213),
            .I(N__11210));
    LocalMux I__1509 (
            .O(N__11210),
            .I(N__11207));
    Odrv4 I__1508 (
            .O(N__11207),
            .I(\this_vga_signals.N_4_i_0_x ));
    CascadeMux I__1507 (
            .O(N__11204),
            .I(N__11201));
    InMux I__1506 (
            .O(N__11201),
            .I(N__11195));
    InMux I__1505 (
            .O(N__11200),
            .I(N__11195));
    LocalMux I__1504 (
            .O(N__11195),
            .I(N__11190));
    InMux I__1503 (
            .O(N__11194),
            .I(N__11185));
    InMux I__1502 (
            .O(N__11193),
            .I(N__11185));
    Odrv4 I__1501 (
            .O(N__11190),
            .I(\this_vga_signals.N_4_i_0_1 ));
    LocalMux I__1500 (
            .O(N__11185),
            .I(\this_vga_signals.N_4_i_0_1 ));
    CascadeMux I__1499 (
            .O(N__11180),
            .I(\this_vga_signals.mult1_un54_sum_ac0_3_0_1_cascade_ ));
    CascadeMux I__1498 (
            .O(N__11177),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    InMux I__1497 (
            .O(N__11174),
            .I(N__11171));
    LocalMux I__1496 (
            .O(N__11171),
            .I(\this_vga_signals.N_57_i_i_0_0 ));
    CascadeMux I__1495 (
            .O(N__11168),
            .I(\this_vga_signals.g0_1_0_cascade_ ));
    InMux I__1494 (
            .O(N__11165),
            .I(N__11162));
    LocalMux I__1493 (
            .O(N__11162),
            .I(\this_vga_signals.N_5_0_0_1 ));
    CascadeMux I__1492 (
            .O(N__11159),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_3_0_0_0_cascade_ ));
    CascadeMux I__1491 (
            .O(N__11156),
            .I(N__11153));
    InMux I__1490 (
            .O(N__11153),
            .I(N__11150));
    LocalMux I__1489 (
            .O(N__11150),
            .I(N__11147));
    Odrv4 I__1488 (
            .O(N__11147),
            .I(this_vga_signals_address_0_i_7));
    InMux I__1487 (
            .O(N__11144),
            .I(N__11141));
    LocalMux I__1486 (
            .O(N__11141),
            .I(\this_vga_signals.N_6_0_0 ));
    InMux I__1485 (
            .O(N__11138),
            .I(N__11135));
    LocalMux I__1484 (
            .O(N__11135),
            .I(\this_vga_signals.mult1_un75_sum_c2_0_0_0_1 ));
    CascadeMux I__1483 (
            .O(N__11132),
            .I(N__11129));
    InMux I__1482 (
            .O(N__11129),
            .I(N__11126));
    LocalMux I__1481 (
            .O(N__11126),
            .I(\this_vga_signals.g3_3_0 ));
    CascadeMux I__1480 (
            .O(N__11123),
            .I(N__11120));
    InMux I__1479 (
            .O(N__11120),
            .I(N__11117));
    LocalMux I__1478 (
            .O(N__11117),
            .I(\this_vga_signals.g3_1_0 ));
    CascadeMux I__1477 (
            .O(N__11114),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_i_cascade_ ));
    CascadeMux I__1476 (
            .O(N__11111),
            .I(N__11108));
    CascadeBuf I__1475 (
            .O(N__11108),
            .I(N__11105));
    CascadeMux I__1474 (
            .O(N__11105),
            .I(N__11102));
    CascadeBuf I__1473 (
            .O(N__11102),
            .I(N__11099));
    CascadeMux I__1472 (
            .O(N__11099),
            .I(N__11096));
    CascadeBuf I__1471 (
            .O(N__11096),
            .I(N__11093));
    CascadeMux I__1470 (
            .O(N__11093),
            .I(N__11090));
    CascadeBuf I__1469 (
            .O(N__11090),
            .I(N__11087));
    CascadeMux I__1468 (
            .O(N__11087),
            .I(N__11084));
    CascadeBuf I__1467 (
            .O(N__11084),
            .I(N__11081));
    CascadeMux I__1466 (
            .O(N__11081),
            .I(N__11078));
    CascadeBuf I__1465 (
            .O(N__11078),
            .I(N__11075));
    CascadeMux I__1464 (
            .O(N__11075),
            .I(N__11072));
    CascadeBuf I__1463 (
            .O(N__11072),
            .I(N__11069));
    CascadeMux I__1462 (
            .O(N__11069),
            .I(N__11066));
    CascadeBuf I__1461 (
            .O(N__11066),
            .I(N__11063));
    CascadeMux I__1460 (
            .O(N__11063),
            .I(N__11060));
    CascadeBuf I__1459 (
            .O(N__11060),
            .I(N__11057));
    CascadeMux I__1458 (
            .O(N__11057),
            .I(N__11054));
    CascadeBuf I__1457 (
            .O(N__11054),
            .I(N__11051));
    CascadeMux I__1456 (
            .O(N__11051),
            .I(N__11048));
    CascadeBuf I__1455 (
            .O(N__11048),
            .I(N__11045));
    CascadeMux I__1454 (
            .O(N__11045),
            .I(N__11042));
    CascadeBuf I__1453 (
            .O(N__11042),
            .I(N__11039));
    CascadeMux I__1452 (
            .O(N__11039),
            .I(N__11036));
    CascadeBuf I__1451 (
            .O(N__11036),
            .I(N__11033));
    CascadeMux I__1450 (
            .O(N__11033),
            .I(N__11030));
    CascadeBuf I__1449 (
            .O(N__11030),
            .I(N__11027));
    CascadeMux I__1448 (
            .O(N__11027),
            .I(N__11024));
    CascadeBuf I__1447 (
            .O(N__11024),
            .I(N__11021));
    CascadeMux I__1446 (
            .O(N__11021),
            .I(N__11018));
    InMux I__1445 (
            .O(N__11018),
            .I(N__11014));
    CascadeMux I__1444 (
            .O(N__11017),
            .I(N__11011));
    LocalMux I__1443 (
            .O(N__11014),
            .I(N__11008));
    InMux I__1442 (
            .O(N__11011),
            .I(N__11005));
    Span4Mux_v I__1441 (
            .O(N__11008),
            .I(N__11002));
    LocalMux I__1440 (
            .O(N__11005),
            .I(N__10999));
    Span4Mux_h I__1439 (
            .O(N__11002),
            .I(N__10996));
    Sp12to4 I__1438 (
            .O(N__10999),
            .I(N__10991));
    Sp12to4 I__1437 (
            .O(N__10996),
            .I(N__10988));
    InMux I__1436 (
            .O(N__10995),
            .I(N__10985));
    InMux I__1435 (
            .O(N__10994),
            .I(N__10982));
    Span12Mux_v I__1434 (
            .O(N__10991),
            .I(N__10977));
    Span12Mux_h I__1433 (
            .O(N__10988),
            .I(N__10977));
    LocalMux I__1432 (
            .O(N__10985),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__1431 (
            .O(N__10982),
            .I(M_this_ppu_vram_addr_0));
    Odrv12 I__1430 (
            .O(N__10977),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__1429 (
            .O(N__10970),
            .I(N__10967));
    CascadeBuf I__1428 (
            .O(N__10967),
            .I(N__10964));
    CascadeMux I__1427 (
            .O(N__10964),
            .I(N__10961));
    CascadeBuf I__1426 (
            .O(N__10961),
            .I(N__10958));
    CascadeMux I__1425 (
            .O(N__10958),
            .I(N__10955));
    CascadeBuf I__1424 (
            .O(N__10955),
            .I(N__10952));
    CascadeMux I__1423 (
            .O(N__10952),
            .I(N__10949));
    CascadeBuf I__1422 (
            .O(N__10949),
            .I(N__10946));
    CascadeMux I__1421 (
            .O(N__10946),
            .I(N__10943));
    CascadeBuf I__1420 (
            .O(N__10943),
            .I(N__10940));
    CascadeMux I__1419 (
            .O(N__10940),
            .I(N__10937));
    CascadeBuf I__1418 (
            .O(N__10937),
            .I(N__10934));
    CascadeMux I__1417 (
            .O(N__10934),
            .I(N__10931));
    CascadeBuf I__1416 (
            .O(N__10931),
            .I(N__10928));
    CascadeMux I__1415 (
            .O(N__10928),
            .I(N__10925));
    CascadeBuf I__1414 (
            .O(N__10925),
            .I(N__10922));
    CascadeMux I__1413 (
            .O(N__10922),
            .I(N__10919));
    CascadeBuf I__1412 (
            .O(N__10919),
            .I(N__10916));
    CascadeMux I__1411 (
            .O(N__10916),
            .I(N__10913));
    CascadeBuf I__1410 (
            .O(N__10913),
            .I(N__10910));
    CascadeMux I__1409 (
            .O(N__10910),
            .I(N__10907));
    CascadeBuf I__1408 (
            .O(N__10907),
            .I(N__10904));
    CascadeMux I__1407 (
            .O(N__10904),
            .I(N__10901));
    CascadeBuf I__1406 (
            .O(N__10901),
            .I(N__10898));
    CascadeMux I__1405 (
            .O(N__10898),
            .I(N__10895));
    CascadeBuf I__1404 (
            .O(N__10895),
            .I(N__10892));
    CascadeMux I__1403 (
            .O(N__10892),
            .I(N__10889));
    CascadeBuf I__1402 (
            .O(N__10889),
            .I(N__10886));
    CascadeMux I__1401 (
            .O(N__10886),
            .I(N__10883));
    CascadeBuf I__1400 (
            .O(N__10883),
            .I(N__10879));
    CascadeMux I__1399 (
            .O(N__10882),
            .I(N__10876));
    CascadeMux I__1398 (
            .O(N__10879),
            .I(N__10873));
    InMux I__1397 (
            .O(N__10876),
            .I(N__10870));
    InMux I__1396 (
            .O(N__10873),
            .I(N__10867));
    LocalMux I__1395 (
            .O(N__10870),
            .I(N__10864));
    LocalMux I__1394 (
            .O(N__10867),
            .I(N__10861));
    Sp12to4 I__1393 (
            .O(N__10864),
            .I(N__10856));
    Span12Mux_s11_h I__1392 (
            .O(N__10861),
            .I(N__10853));
    InMux I__1391 (
            .O(N__10860),
            .I(N__10850));
    InMux I__1390 (
            .O(N__10859),
            .I(N__10847));
    Span12Mux_v I__1389 (
            .O(N__10856),
            .I(N__10842));
    Span12Mux_h I__1388 (
            .O(N__10853),
            .I(N__10842));
    LocalMux I__1387 (
            .O(N__10850),
            .I(M_this_ppu_vram_addr_3));
    LocalMux I__1386 (
            .O(N__10847),
            .I(M_this_ppu_vram_addr_3));
    Odrv12 I__1385 (
            .O(N__10842),
            .I(M_this_ppu_vram_addr_3));
    CascadeMux I__1384 (
            .O(N__10835),
            .I(N__10832));
    CascadeBuf I__1383 (
            .O(N__10832),
            .I(N__10829));
    CascadeMux I__1382 (
            .O(N__10829),
            .I(N__10826));
    CascadeBuf I__1381 (
            .O(N__10826),
            .I(N__10823));
    CascadeMux I__1380 (
            .O(N__10823),
            .I(N__10820));
    CascadeBuf I__1379 (
            .O(N__10820),
            .I(N__10817));
    CascadeMux I__1378 (
            .O(N__10817),
            .I(N__10814));
    CascadeBuf I__1377 (
            .O(N__10814),
            .I(N__10811));
    CascadeMux I__1376 (
            .O(N__10811),
            .I(N__10808));
    CascadeBuf I__1375 (
            .O(N__10808),
            .I(N__10805));
    CascadeMux I__1374 (
            .O(N__10805),
            .I(N__10802));
    CascadeBuf I__1373 (
            .O(N__10802),
            .I(N__10799));
    CascadeMux I__1372 (
            .O(N__10799),
            .I(N__10796));
    CascadeBuf I__1371 (
            .O(N__10796),
            .I(N__10793));
    CascadeMux I__1370 (
            .O(N__10793),
            .I(N__10790));
    CascadeBuf I__1369 (
            .O(N__10790),
            .I(N__10787));
    CascadeMux I__1368 (
            .O(N__10787),
            .I(N__10784));
    CascadeBuf I__1367 (
            .O(N__10784),
            .I(N__10781));
    CascadeMux I__1366 (
            .O(N__10781),
            .I(N__10778));
    CascadeBuf I__1365 (
            .O(N__10778),
            .I(N__10775));
    CascadeMux I__1364 (
            .O(N__10775),
            .I(N__10772));
    CascadeBuf I__1363 (
            .O(N__10772),
            .I(N__10769));
    CascadeMux I__1362 (
            .O(N__10769),
            .I(N__10766));
    CascadeBuf I__1361 (
            .O(N__10766),
            .I(N__10763));
    CascadeMux I__1360 (
            .O(N__10763),
            .I(N__10760));
    CascadeBuf I__1359 (
            .O(N__10760),
            .I(N__10757));
    CascadeMux I__1358 (
            .O(N__10757),
            .I(N__10754));
    CascadeBuf I__1357 (
            .O(N__10754),
            .I(N__10751));
    CascadeMux I__1356 (
            .O(N__10751),
            .I(N__10748));
    CascadeBuf I__1355 (
            .O(N__10748),
            .I(N__10745));
    CascadeMux I__1354 (
            .O(N__10745),
            .I(N__10742));
    InMux I__1353 (
            .O(N__10742),
            .I(N__10739));
    LocalMux I__1352 (
            .O(N__10739),
            .I(N__10735));
    CascadeMux I__1351 (
            .O(N__10738),
            .I(N__10732));
    Span4Mux_s3_v I__1350 (
            .O(N__10735),
            .I(N__10729));
    InMux I__1349 (
            .O(N__10732),
            .I(N__10725));
    Span4Mux_h I__1348 (
            .O(N__10729),
            .I(N__10722));
    CascadeMux I__1347 (
            .O(N__10728),
            .I(N__10718));
    LocalMux I__1346 (
            .O(N__10725),
            .I(N__10715));
    Sp12to4 I__1345 (
            .O(N__10722),
            .I(N__10712));
    InMux I__1344 (
            .O(N__10721),
            .I(N__10709));
    InMux I__1343 (
            .O(N__10718),
            .I(N__10706));
    Sp12to4 I__1342 (
            .O(N__10715),
            .I(N__10703));
    Span12Mux_h I__1341 (
            .O(N__10712),
            .I(N__10700));
    LocalMux I__1340 (
            .O(N__10709),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__1339 (
            .O(N__10706),
            .I(M_this_ppu_vram_addr_1));
    Odrv12 I__1338 (
            .O(N__10703),
            .I(M_this_ppu_vram_addr_1));
    Odrv12 I__1337 (
            .O(N__10700),
            .I(M_this_ppu_vram_addr_1));
    InMux I__1336 (
            .O(N__10691),
            .I(N__10688));
    LocalMux I__1335 (
            .O(N__10688),
            .I(\this_ppu.un1_M_state_d8_5_0 ));
    CascadeMux I__1334 (
            .O(N__10685),
            .I(M_this_sprites_ram_read_data_0_cascade_));
    InMux I__1333 (
            .O(N__10682),
            .I(N__10679));
    LocalMux I__1332 (
            .O(N__10679),
            .I(N__10676));
    Span12Mux_v I__1331 (
            .O(N__10676),
            .I(N__10673));
    Odrv12 I__1330 (
            .O(N__10673),
            .I(M_this_vram_write_data_0));
    InMux I__1329 (
            .O(N__10670),
            .I(N__10667));
    LocalMux I__1328 (
            .O(N__10667),
            .I(N__10664));
    Span12Mux_h I__1327 (
            .O(N__10664),
            .I(N__10661));
    Odrv12 I__1326 (
            .O(N__10661),
            .I(port_clk_c));
    InMux I__1325 (
            .O(N__10658),
            .I(N__10655));
    LocalMux I__1324 (
            .O(N__10655),
            .I(N__10652));
    Span4Mux_v I__1323 (
            .O(N__10652),
            .I(N__10649));
    Odrv4 I__1322 (
            .O(N__10649),
            .I(\this_vga_signals.vsync_1_0_a2_6_a2_1_0 ));
    IoInMux I__1321 (
            .O(N__10646),
            .I(N__10643));
    LocalMux I__1320 (
            .O(N__10643),
            .I(N__10640));
    Span4Mux_s0_v I__1319 (
            .O(N__10640),
            .I(N__10637));
    Sp12to4 I__1318 (
            .O(N__10637),
            .I(N__10634));
    Span12Mux_s7_h I__1317 (
            .O(N__10634),
            .I(N__10631));
    Span12Mux_v I__1316 (
            .O(N__10631),
            .I(N__10628));
    Odrv12 I__1315 (
            .O(N__10628),
            .I(this_vga_signals_vsync_1_i));
    InMux I__1314 (
            .O(N__10625),
            .I(N__10622));
    LocalMux I__1313 (
            .O(N__10622),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    InMux I__1312 (
            .O(N__10619),
            .I(N__10616));
    LocalMux I__1311 (
            .O(N__10616),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    CascadeMux I__1310 (
            .O(N__10613),
            .I(\this_vga_signals.g0_16_x0_cascade_ ));
    InMux I__1309 (
            .O(N__10610),
            .I(N__10607));
    LocalMux I__1308 (
            .O(N__10607),
            .I(\this_vga_signals.g3_0 ));
    CascadeMux I__1307 (
            .O(N__10604),
            .I(this_vga_signals_un4_lcounter_if_i1_mux_cascade_));
    InMux I__1306 (
            .O(N__10601),
            .I(N__10595));
    InMux I__1305 (
            .O(N__10600),
            .I(N__10592));
    InMux I__1304 (
            .O(N__10599),
            .I(N__10587));
    InMux I__1303 (
            .O(N__10598),
            .I(N__10587));
    LocalMux I__1302 (
            .O(N__10595),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0));
    LocalMux I__1301 (
            .O(N__10592),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0));
    LocalMux I__1300 (
            .O(N__10587),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0));
    CascadeMux I__1299 (
            .O(N__10580),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_cascade_));
    InMux I__1298 (
            .O(N__10577),
            .I(N__10573));
    InMux I__1297 (
            .O(N__10576),
            .I(N__10570));
    LocalMux I__1296 (
            .O(N__10573),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1));
    LocalMux I__1295 (
            .O(N__10570),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1));
    InMux I__1294 (
            .O(N__10565),
            .I(N__10562));
    LocalMux I__1293 (
            .O(N__10562),
            .I(\this_ppu.M_m7Z0Z_1 ));
    InMux I__1292 (
            .O(N__10559),
            .I(N__10556));
    LocalMux I__1291 (
            .O(N__10556),
            .I(N__10553));
    Odrv4 I__1290 (
            .O(N__10553),
            .I(\this_ppu.M_m12_0_o2_381_10Z0Z_1 ));
    CascadeMux I__1289 (
            .O(N__10550),
            .I(\this_ppu.M_N_11_mux_cascade_ ));
    InMux I__1288 (
            .O(N__10547),
            .I(N__10543));
    InMux I__1287 (
            .O(N__10546),
            .I(N__10540));
    LocalMux I__1286 (
            .O(N__10543),
            .I(\this_ppu.M_m12_0_o2_381_10 ));
    LocalMux I__1285 (
            .O(N__10540),
            .I(\this_ppu.M_m12_0_o2_381_10 ));
    InMux I__1284 (
            .O(N__10535),
            .I(N__10531));
    InMux I__1283 (
            .O(N__10534),
            .I(N__10528));
    LocalMux I__1282 (
            .O(N__10531),
            .I(this_vga_signals_un4_lcounter_if_i1_mux));
    LocalMux I__1281 (
            .O(N__10528),
            .I(this_vga_signals_un4_lcounter_if_i1_mux));
    CascadeMux I__1280 (
            .O(N__10523),
            .I(N__10520));
    InMux I__1279 (
            .O(N__10520),
            .I(N__10515));
    InMux I__1278 (
            .O(N__10519),
            .I(N__10512));
    InMux I__1277 (
            .O(N__10518),
            .I(N__10509));
    LocalMux I__1276 (
            .O(N__10515),
            .I(N__10504));
    LocalMux I__1275 (
            .O(N__10512),
            .I(N__10504));
    LocalMux I__1274 (
            .O(N__10509),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1));
    Odrv4 I__1273 (
            .O(N__10504),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1));
    InMux I__1272 (
            .O(N__10499),
            .I(N__10496));
    LocalMux I__1271 (
            .O(N__10496),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_1));
    InMux I__1270 (
            .O(N__10493),
            .I(N__10486));
    InMux I__1269 (
            .O(N__10492),
            .I(N__10486));
    InMux I__1268 (
            .O(N__10491),
            .I(N__10483));
    LocalMux I__1267 (
            .O(N__10486),
            .I(this_vga_signals_un4_lcounter_if_N_7_i_i));
    LocalMux I__1266 (
            .O(N__10483),
            .I(this_vga_signals_un4_lcounter_if_N_7_i_i));
    CascadeMux I__1265 (
            .O(N__10478),
            .I(N__10475));
    CascadeBuf I__1264 (
            .O(N__10475),
            .I(N__10472));
    CascadeMux I__1263 (
            .O(N__10472),
            .I(N__10469));
    CascadeBuf I__1262 (
            .O(N__10469),
            .I(N__10466));
    CascadeMux I__1261 (
            .O(N__10466),
            .I(N__10463));
    CascadeBuf I__1260 (
            .O(N__10463),
            .I(N__10460));
    CascadeMux I__1259 (
            .O(N__10460),
            .I(N__10457));
    CascadeBuf I__1258 (
            .O(N__10457),
            .I(N__10454));
    CascadeMux I__1257 (
            .O(N__10454),
            .I(N__10451));
    CascadeBuf I__1256 (
            .O(N__10451),
            .I(N__10448));
    CascadeMux I__1255 (
            .O(N__10448),
            .I(N__10445));
    CascadeBuf I__1254 (
            .O(N__10445),
            .I(N__10442));
    CascadeMux I__1253 (
            .O(N__10442),
            .I(N__10439));
    CascadeBuf I__1252 (
            .O(N__10439),
            .I(N__10436));
    CascadeMux I__1251 (
            .O(N__10436),
            .I(N__10433));
    CascadeBuf I__1250 (
            .O(N__10433),
            .I(N__10430));
    CascadeMux I__1249 (
            .O(N__10430),
            .I(N__10427));
    CascadeBuf I__1248 (
            .O(N__10427),
            .I(N__10424));
    CascadeMux I__1247 (
            .O(N__10424),
            .I(N__10421));
    CascadeBuf I__1246 (
            .O(N__10421),
            .I(N__10418));
    CascadeMux I__1245 (
            .O(N__10418),
            .I(N__10415));
    CascadeBuf I__1244 (
            .O(N__10415),
            .I(N__10412));
    CascadeMux I__1243 (
            .O(N__10412),
            .I(N__10409));
    CascadeBuf I__1242 (
            .O(N__10409),
            .I(N__10406));
    CascadeMux I__1241 (
            .O(N__10406),
            .I(N__10403));
    CascadeBuf I__1240 (
            .O(N__10403),
            .I(N__10400));
    CascadeMux I__1239 (
            .O(N__10400),
            .I(N__10397));
    CascadeBuf I__1238 (
            .O(N__10397),
            .I(N__10394));
    CascadeMux I__1237 (
            .O(N__10394),
            .I(N__10391));
    CascadeBuf I__1236 (
            .O(N__10391),
            .I(N__10388));
    CascadeMux I__1235 (
            .O(N__10388),
            .I(N__10385));
    InMux I__1234 (
            .O(N__10385),
            .I(N__10382));
    LocalMux I__1233 (
            .O(N__10382),
            .I(N__10378));
    CascadeMux I__1232 (
            .O(N__10381),
            .I(N__10375));
    Span4Mux_h I__1231 (
            .O(N__10378),
            .I(N__10372));
    InMux I__1230 (
            .O(N__10375),
            .I(N__10369));
    Span4Mux_h I__1229 (
            .O(N__10372),
            .I(N__10366));
    LocalMux I__1228 (
            .O(N__10369),
            .I(N__10361));
    Sp12to4 I__1227 (
            .O(N__10366),
            .I(N__10358));
    InMux I__1226 (
            .O(N__10365),
            .I(N__10355));
    InMux I__1225 (
            .O(N__10364),
            .I(N__10352));
    Span12Mux_v I__1224 (
            .O(N__10361),
            .I(N__10347));
    Span12Mux_v I__1223 (
            .O(N__10358),
            .I(N__10347));
    LocalMux I__1222 (
            .O(N__10355),
            .I(M_this_ppu_vram_addr_5));
    LocalMux I__1221 (
            .O(N__10352),
            .I(M_this_ppu_vram_addr_5));
    Odrv12 I__1220 (
            .O(N__10347),
            .I(M_this_ppu_vram_addr_5));
    CascadeMux I__1219 (
            .O(N__10340),
            .I(N__10337));
    CascadeBuf I__1218 (
            .O(N__10337),
            .I(N__10334));
    CascadeMux I__1217 (
            .O(N__10334),
            .I(N__10331));
    CascadeBuf I__1216 (
            .O(N__10331),
            .I(N__10328));
    CascadeMux I__1215 (
            .O(N__10328),
            .I(N__10325));
    CascadeBuf I__1214 (
            .O(N__10325),
            .I(N__10322));
    CascadeMux I__1213 (
            .O(N__10322),
            .I(N__10319));
    CascadeBuf I__1212 (
            .O(N__10319),
            .I(N__10316));
    CascadeMux I__1211 (
            .O(N__10316),
            .I(N__10313));
    CascadeBuf I__1210 (
            .O(N__10313),
            .I(N__10310));
    CascadeMux I__1209 (
            .O(N__10310),
            .I(N__10307));
    CascadeBuf I__1208 (
            .O(N__10307),
            .I(N__10304));
    CascadeMux I__1207 (
            .O(N__10304),
            .I(N__10301));
    CascadeBuf I__1206 (
            .O(N__10301),
            .I(N__10298));
    CascadeMux I__1205 (
            .O(N__10298),
            .I(N__10295));
    CascadeBuf I__1204 (
            .O(N__10295),
            .I(N__10292));
    CascadeMux I__1203 (
            .O(N__10292),
            .I(N__10289));
    CascadeBuf I__1202 (
            .O(N__10289),
            .I(N__10286));
    CascadeMux I__1201 (
            .O(N__10286),
            .I(N__10283));
    CascadeBuf I__1200 (
            .O(N__10283),
            .I(N__10280));
    CascadeMux I__1199 (
            .O(N__10280),
            .I(N__10277));
    CascadeBuf I__1198 (
            .O(N__10277),
            .I(N__10274));
    CascadeMux I__1197 (
            .O(N__10274),
            .I(N__10271));
    CascadeBuf I__1196 (
            .O(N__10271),
            .I(N__10268));
    CascadeMux I__1195 (
            .O(N__10268),
            .I(N__10265));
    CascadeBuf I__1194 (
            .O(N__10265),
            .I(N__10262));
    CascadeMux I__1193 (
            .O(N__10262),
            .I(N__10259));
    CascadeBuf I__1192 (
            .O(N__10259),
            .I(N__10256));
    CascadeMux I__1191 (
            .O(N__10256),
            .I(N__10253));
    CascadeBuf I__1190 (
            .O(N__10253),
            .I(N__10250));
    CascadeMux I__1189 (
            .O(N__10250),
            .I(N__10247));
    InMux I__1188 (
            .O(N__10247),
            .I(N__10243));
    CascadeMux I__1187 (
            .O(N__10246),
            .I(N__10240));
    LocalMux I__1186 (
            .O(N__10243),
            .I(N__10237));
    InMux I__1185 (
            .O(N__10240),
            .I(N__10234));
    Span4Mux_s2_v I__1184 (
            .O(N__10237),
            .I(N__10231));
    LocalMux I__1183 (
            .O(N__10234),
            .I(N__10228));
    Span4Mux_h I__1182 (
            .O(N__10231),
            .I(N__10225));
    Span4Mux_v I__1181 (
            .O(N__10228),
            .I(N__10220));
    Sp12to4 I__1180 (
            .O(N__10225),
            .I(N__10217));
    InMux I__1179 (
            .O(N__10224),
            .I(N__10214));
    InMux I__1178 (
            .O(N__10223),
            .I(N__10211));
    Span4Mux_v I__1177 (
            .O(N__10220),
            .I(N__10208));
    Span12Mux_v I__1176 (
            .O(N__10217),
            .I(N__10205));
    LocalMux I__1175 (
            .O(N__10214),
            .I(M_this_ppu_vram_addr_4));
    LocalMux I__1174 (
            .O(N__10211),
            .I(M_this_ppu_vram_addr_4));
    Odrv4 I__1173 (
            .O(N__10208),
            .I(M_this_ppu_vram_addr_4));
    Odrv12 I__1172 (
            .O(N__10205),
            .I(M_this_ppu_vram_addr_4));
    CascadeMux I__1171 (
            .O(N__10196),
            .I(N__10193));
    CascadeBuf I__1170 (
            .O(N__10193),
            .I(N__10190));
    CascadeMux I__1169 (
            .O(N__10190),
            .I(N__10187));
    CascadeBuf I__1168 (
            .O(N__10187),
            .I(N__10184));
    CascadeMux I__1167 (
            .O(N__10184),
            .I(N__10181));
    CascadeBuf I__1166 (
            .O(N__10181),
            .I(N__10178));
    CascadeMux I__1165 (
            .O(N__10178),
            .I(N__10175));
    CascadeBuf I__1164 (
            .O(N__10175),
            .I(N__10172));
    CascadeMux I__1163 (
            .O(N__10172),
            .I(N__10169));
    CascadeBuf I__1162 (
            .O(N__10169),
            .I(N__10166));
    CascadeMux I__1161 (
            .O(N__10166),
            .I(N__10163));
    CascadeBuf I__1160 (
            .O(N__10163),
            .I(N__10160));
    CascadeMux I__1159 (
            .O(N__10160),
            .I(N__10157));
    CascadeBuf I__1158 (
            .O(N__10157),
            .I(N__10154));
    CascadeMux I__1157 (
            .O(N__10154),
            .I(N__10151));
    CascadeBuf I__1156 (
            .O(N__10151),
            .I(N__10148));
    CascadeMux I__1155 (
            .O(N__10148),
            .I(N__10145));
    CascadeBuf I__1154 (
            .O(N__10145),
            .I(N__10142));
    CascadeMux I__1153 (
            .O(N__10142),
            .I(N__10139));
    CascadeBuf I__1152 (
            .O(N__10139),
            .I(N__10136));
    CascadeMux I__1151 (
            .O(N__10136),
            .I(N__10133));
    CascadeBuf I__1150 (
            .O(N__10133),
            .I(N__10130));
    CascadeMux I__1149 (
            .O(N__10130),
            .I(N__10127));
    CascadeBuf I__1148 (
            .O(N__10127),
            .I(N__10124));
    CascadeMux I__1147 (
            .O(N__10124),
            .I(N__10121));
    CascadeBuf I__1146 (
            .O(N__10121),
            .I(N__10118));
    CascadeMux I__1145 (
            .O(N__10118),
            .I(N__10115));
    CascadeBuf I__1144 (
            .O(N__10115),
            .I(N__10112));
    CascadeMux I__1143 (
            .O(N__10112),
            .I(N__10109));
    CascadeBuf I__1142 (
            .O(N__10109),
            .I(N__10106));
    CascadeMux I__1141 (
            .O(N__10106),
            .I(N__10103));
    InMux I__1140 (
            .O(N__10103),
            .I(N__10100));
    LocalMux I__1139 (
            .O(N__10100),
            .I(N__10096));
    CascadeMux I__1138 (
            .O(N__10099),
            .I(N__10093));
    Span4Mux_s2_v I__1137 (
            .O(N__10096),
            .I(N__10090));
    InMux I__1136 (
            .O(N__10093),
            .I(N__10087));
    Span4Mux_h I__1135 (
            .O(N__10090),
            .I(N__10084));
    LocalMux I__1134 (
            .O(N__10087),
            .I(N__10080));
    Span4Mux_v I__1133 (
            .O(N__10084),
            .I(N__10077));
    CascadeMux I__1132 (
            .O(N__10083),
            .I(N__10074));
    Span4Mux_v I__1131 (
            .O(N__10080),
            .I(N__10070));
    Sp12to4 I__1130 (
            .O(N__10077),
            .I(N__10067));
    InMux I__1129 (
            .O(N__10074),
            .I(N__10064));
    InMux I__1128 (
            .O(N__10073),
            .I(N__10061));
    Sp12to4 I__1127 (
            .O(N__10070),
            .I(N__10056));
    Span12Mux_h I__1126 (
            .O(N__10067),
            .I(N__10056));
    LocalMux I__1125 (
            .O(N__10064),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__1124 (
            .O(N__10061),
            .I(M_this_ppu_vram_addr_6));
    Odrv12 I__1123 (
            .O(N__10056),
            .I(M_this_ppu_vram_addr_6));
    CascadeMux I__1122 (
            .O(N__10049),
            .I(N__10046));
    CascadeBuf I__1121 (
            .O(N__10046),
            .I(N__10043));
    CascadeMux I__1120 (
            .O(N__10043),
            .I(N__10040));
    CascadeBuf I__1119 (
            .O(N__10040),
            .I(N__10037));
    CascadeMux I__1118 (
            .O(N__10037),
            .I(N__10034));
    CascadeBuf I__1117 (
            .O(N__10034),
            .I(N__10031));
    CascadeMux I__1116 (
            .O(N__10031),
            .I(N__10028));
    CascadeBuf I__1115 (
            .O(N__10028),
            .I(N__10025));
    CascadeMux I__1114 (
            .O(N__10025),
            .I(N__10022));
    CascadeBuf I__1113 (
            .O(N__10022),
            .I(N__10019));
    CascadeMux I__1112 (
            .O(N__10019),
            .I(N__10016));
    CascadeBuf I__1111 (
            .O(N__10016),
            .I(N__10013));
    CascadeMux I__1110 (
            .O(N__10013),
            .I(N__10010));
    CascadeBuf I__1109 (
            .O(N__10010),
            .I(N__10007));
    CascadeMux I__1108 (
            .O(N__10007),
            .I(N__10004));
    CascadeBuf I__1107 (
            .O(N__10004),
            .I(N__10001));
    CascadeMux I__1106 (
            .O(N__10001),
            .I(N__9998));
    CascadeBuf I__1105 (
            .O(N__9998),
            .I(N__9995));
    CascadeMux I__1104 (
            .O(N__9995),
            .I(N__9992));
    CascadeBuf I__1103 (
            .O(N__9992),
            .I(N__9989));
    CascadeMux I__1102 (
            .O(N__9989),
            .I(N__9986));
    CascadeBuf I__1101 (
            .O(N__9986),
            .I(N__9983));
    CascadeMux I__1100 (
            .O(N__9983),
            .I(N__9980));
    CascadeBuf I__1099 (
            .O(N__9980),
            .I(N__9977));
    CascadeMux I__1098 (
            .O(N__9977),
            .I(N__9974));
    CascadeBuf I__1097 (
            .O(N__9974),
            .I(N__9971));
    CascadeMux I__1096 (
            .O(N__9971),
            .I(N__9968));
    CascadeBuf I__1095 (
            .O(N__9968),
            .I(N__9965));
    CascadeMux I__1094 (
            .O(N__9965),
            .I(N__9962));
    CascadeBuf I__1093 (
            .O(N__9962),
            .I(N__9959));
    CascadeMux I__1092 (
            .O(N__9959),
            .I(N__9956));
    InMux I__1091 (
            .O(N__9956),
            .I(N__9953));
    LocalMux I__1090 (
            .O(N__9953),
            .I(N__9949));
    CascadeMux I__1089 (
            .O(N__9952),
            .I(N__9946));
    Span4Mux_s2_v I__1088 (
            .O(N__9949),
            .I(N__9943));
    InMux I__1087 (
            .O(N__9946),
            .I(N__9940));
    Span4Mux_h I__1086 (
            .O(N__9943),
            .I(N__9937));
    LocalMux I__1085 (
            .O(N__9940),
            .I(N__9932));
    Sp12to4 I__1084 (
            .O(N__9937),
            .I(N__9929));
    InMux I__1083 (
            .O(N__9936),
            .I(N__9926));
    InMux I__1082 (
            .O(N__9935),
            .I(N__9923));
    Span12Mux_s8_h I__1081 (
            .O(N__9932),
            .I(N__9920));
    Span12Mux_h I__1080 (
            .O(N__9929),
            .I(N__9917));
    LocalMux I__1079 (
            .O(N__9926),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__1078 (
            .O(N__9923),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__1077 (
            .O(N__9920),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__1076 (
            .O(N__9917),
            .I(M_this_ppu_vram_addr_2));
    CascadeMux I__1075 (
            .O(N__9908),
            .I(\this_ppu.un1_M_state_d8_4_0_cascade_ ));
    InMux I__1074 (
            .O(N__9905),
            .I(N__9902));
    LocalMux I__1073 (
            .O(N__9902),
            .I(\this_ppu.M_N_3_mux_0_0 ));
    InMux I__1072 (
            .O(N__9899),
            .I(N__9896));
    LocalMux I__1071 (
            .O(N__9896),
            .I(N__9891));
    InMux I__1070 (
            .O(N__9895),
            .I(N__9888));
    InMux I__1069 (
            .O(N__9894),
            .I(N__9885));
    Odrv4 I__1068 (
            .O(N__9891),
            .I(\this_vga_signals.CO1_5_0 ));
    LocalMux I__1067 (
            .O(N__9888),
            .I(\this_vga_signals.CO1_5_0 ));
    LocalMux I__1066 (
            .O(N__9885),
            .I(\this_vga_signals.CO1_5_0 ));
    CascadeMux I__1065 (
            .O(N__9878),
            .I(\this_vga_signals.mult1_un40_sum0_2_cascade_ ));
    CascadeMux I__1064 (
            .O(N__9875),
            .I(\this_vga_signals.mult1_un40_sum_m_ns_2_cascade_ ));
    InMux I__1063 (
            .O(N__9872),
            .I(N__9869));
    LocalMux I__1062 (
            .O(N__9869),
            .I(N__9865));
    InMux I__1061 (
            .O(N__9868),
            .I(N__9862));
    Span4Mux_h I__1060 (
            .O(N__9865),
            .I(N__9859));
    LocalMux I__1059 (
            .O(N__9862),
            .I(N__9856));
    Odrv4 I__1058 (
            .O(N__9859),
            .I(\this_vga_signals.N_196_0 ));
    Odrv4 I__1057 (
            .O(N__9856),
            .I(\this_vga_signals.N_196_0 ));
    CascadeMux I__1056 (
            .O(N__9851),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0_cascade_));
    InMux I__1055 (
            .O(N__9848),
            .I(N__9842));
    InMux I__1054 (
            .O(N__9847),
            .I(N__9842));
    LocalMux I__1053 (
            .O(N__9842),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1));
    CascadeMux I__1052 (
            .O(N__9839),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_cascade_));
    InMux I__1051 (
            .O(N__9836),
            .I(N__9832));
    InMux I__1050 (
            .O(N__9835),
            .I(N__9829));
    LocalMux I__1049 (
            .O(N__9832),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0));
    LocalMux I__1048 (
            .O(N__9829),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0));
    CascadeMux I__1047 (
            .O(N__9824),
            .I(\this_vga_signals.mult1_un40_sum_0_c3_0_cascade_ ));
    CascadeMux I__1046 (
            .O(N__9821),
            .I(N__9818));
    InMux I__1045 (
            .O(N__9818),
            .I(N__9814));
    InMux I__1044 (
            .O(N__9817),
            .I(N__9811));
    LocalMux I__1043 (
            .O(N__9814),
            .I(N__9808));
    LocalMux I__1042 (
            .O(N__9811),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    Odrv4 I__1041 (
            .O(N__9808),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    InMux I__1040 (
            .O(N__9803),
            .I(N__9799));
    InMux I__1039 (
            .O(N__9802),
            .I(N__9796));
    LocalMux I__1038 (
            .O(N__9799),
            .I(N__9793));
    LocalMux I__1037 (
            .O(N__9796),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    Odrv4 I__1036 (
            .O(N__9793),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__1035 (
            .O(N__9788),
            .I(N__9785));
    LocalMux I__1034 (
            .O(N__9785),
            .I(N__9781));
    InMux I__1033 (
            .O(N__9784),
            .I(N__9778));
    Odrv4 I__1032 (
            .O(N__9781),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__1031 (
            .O(N__9778),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    InMux I__1030 (
            .O(N__9773),
            .I(N__9770));
    LocalMux I__1029 (
            .O(N__9770),
            .I(\this_vga_signals.mult1_un40_sum_0_c3_0 ));
    InMux I__1028 (
            .O(N__9767),
            .I(N__9764));
    LocalMux I__1027 (
            .O(N__9764),
            .I(\this_vga_signals.mult1_un40_sum_1_c2_0 ));
    CascadeMux I__1026 (
            .O(N__9761),
            .I(\this_vga_signals.mult1_un40_sum_m_x1_3_cascade_ ));
    InMux I__1025 (
            .O(N__9758),
            .I(N__9755));
    LocalMux I__1024 (
            .O(N__9755),
            .I(\this_vga_signals.mult1_un40_sum_m_x0_3 ));
    InMux I__1023 (
            .O(N__9752),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__1022 (
            .O(N__9749),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__1021 (
            .O(N__9746),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__1020 (
            .O(N__9743),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__1019 (
            .O(N__9740),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__1018 (
            .O(N__9737),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__1017 (
            .O(N__9734),
            .I(bfn_10_15_0_));
    InMux I__1016 (
            .O(N__9731),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    CascadeMux I__1015 (
            .O(N__9728),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_1_0_cascade_ ));
    CascadeMux I__1014 (
            .O(N__9725),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    InMux I__1013 (
            .O(N__9722),
            .I(N__9719));
    LocalMux I__1012 (
            .O(N__9719),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_1_0_0 ));
    InMux I__1011 (
            .O(N__9716),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    CascadeMux I__1010 (
            .O(N__9713),
            .I(\this_vga_signals.g0_3_0_a3_2_cascade_ ));
    InMux I__1009 (
            .O(N__9710),
            .I(N__9707));
    LocalMux I__1008 (
            .O(N__9707),
            .I(\this_vga_signals.g2_1 ));
    InMux I__1007 (
            .O(N__9704),
            .I(N__9701));
    LocalMux I__1006 (
            .O(N__9701),
            .I(N__9698));
    Odrv4 I__1005 (
            .O(N__9698),
            .I(\this_vga_signals.g1_0_0_0 ));
    CascadeMux I__1004 (
            .O(N__9695),
            .I(\this_vga_signals.N_188_0_cascade_ ));
    CascadeMux I__1003 (
            .O(N__9692),
            .I(N__9689));
    InMux I__1002 (
            .O(N__9689),
            .I(N__9686));
    LocalMux I__1001 (
            .O(N__9686),
            .I(\this_vga_signals.if_m10_0_a4_0_0 ));
    CascadeMux I__1000 (
            .O(N__9683),
            .I(\this_vga_signals.g1_3_0_cascade_ ));
    InMux I__999 (
            .O(N__9680),
            .I(N__9677));
    LocalMux I__998 (
            .O(N__9677),
            .I(\this_vga_signals.if_m10_0_a4_1_1 ));
    InMux I__997 (
            .O(N__9674),
            .I(N__9671));
    LocalMux I__996 (
            .O(N__9671),
            .I(\this_vga_signals.if_N_18_0 ));
    CascadeMux I__995 (
            .O(N__9668),
            .I(N__9664));
    InMux I__994 (
            .O(N__9667),
            .I(N__9661));
    InMux I__993 (
            .O(N__9664),
            .I(N__9658));
    LocalMux I__992 (
            .O(N__9661),
            .I(\this_vga_signals.N_3_1 ));
    LocalMux I__991 (
            .O(N__9658),
            .I(\this_vga_signals.N_3_1 ));
    CascadeMux I__990 (
            .O(N__9653),
            .I(N__9650));
    InMux I__989 (
            .O(N__9650),
            .I(N__9644));
    InMux I__988 (
            .O(N__9649),
            .I(N__9644));
    LocalMux I__987 (
            .O(N__9644),
            .I(\this_vga_signals.m6_2 ));
    CascadeMux I__986 (
            .O(N__9641),
            .I(N__9638));
    InMux I__985 (
            .O(N__9638),
            .I(N__9635));
    LocalMux I__984 (
            .O(N__9635),
            .I(N__9632));
    Odrv4 I__983 (
            .O(N__9632),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_0_0 ));
    InMux I__982 (
            .O(N__9629),
            .I(N__9626));
    LocalMux I__981 (
            .O(N__9626),
            .I(N__9621));
    InMux I__980 (
            .O(N__9625),
            .I(N__9618));
    InMux I__979 (
            .O(N__9624),
            .I(N__9615));
    Odrv4 I__978 (
            .O(N__9621),
            .I(\this_vga_signals.if_i3_mux_0_0 ));
    LocalMux I__977 (
            .O(N__9618),
            .I(\this_vga_signals.if_i3_mux_0_0 ));
    LocalMux I__976 (
            .O(N__9615),
            .I(\this_vga_signals.if_i3_mux_0_0 ));
    InMux I__975 (
            .O(N__9608),
            .I(N__9605));
    LocalMux I__974 (
            .O(N__9605),
            .I(\this_vga_signals.M_vcounter_q_RNI820378Z0Z_2 ));
    CascadeMux I__973 (
            .O(N__9602),
            .I(\this_vga_signals.N_3_0_cascade_ ));
    CascadeMux I__972 (
            .O(N__9599),
            .I(\this_vga_signals.g1_cascade_ ));
    InMux I__971 (
            .O(N__9596),
            .I(N__9593));
    LocalMux I__970 (
            .O(N__9593),
            .I(\this_vga_signals.mult1_un68_sum_c3_0 ));
    InMux I__969 (
            .O(N__9590),
            .I(N__9587));
    LocalMux I__968 (
            .O(N__9587),
            .I(\this_vga_signals.M_vcounter_q_RNI820378_0Z0Z_2 ));
    InMux I__967 (
            .O(N__9584),
            .I(N__9580));
    InMux I__966 (
            .O(N__9583),
            .I(N__9577));
    LocalMux I__965 (
            .O(N__9580),
            .I(\this_vga_signals.N_9_0_0 ));
    LocalMux I__964 (
            .O(N__9577),
            .I(\this_vga_signals.N_9_0_0 ));
    CascadeMux I__963 (
            .O(N__9572),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIDB4TM3Z0Z_5_cascade_ ));
    InMux I__962 (
            .O(N__9569),
            .I(N__9566));
    LocalMux I__961 (
            .O(N__9566),
            .I(\this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0Z0Z_5 ));
    InMux I__960 (
            .O(N__9563),
            .I(N__9560));
    LocalMux I__959 (
            .O(N__9560),
            .I(N__9557));
    Odrv4 I__958 (
            .O(N__9557),
            .I(\this_vga_signals.N_5 ));
    CascadeMux I__957 (
            .O(N__9554),
            .I(\this_vga_signals.g0_0_x2_0_0_a3_3_cascade_ ));
    CascadeMux I__956 (
            .O(N__9551),
            .I(\this_vga_signals.N_9_i_0_0_cascade_ ));
    InMux I__955 (
            .O(N__9548),
            .I(N__9545));
    LocalMux I__954 (
            .O(N__9545),
            .I(\this_vga_signals.N_9_i_0_0 ));
    CascadeMux I__953 (
            .O(N__9542),
            .I(\this_vga_signals.g0_2_x0_cascade_ ));
    InMux I__952 (
            .O(N__9539),
            .I(N__9536));
    LocalMux I__951 (
            .O(N__9536),
            .I(\this_vga_signals.g0_2_x1 ));
    InMux I__950 (
            .O(N__9533),
            .I(\this_ppu.un1_M_current_q_cry_0 ));
    InMux I__949 (
            .O(N__9530),
            .I(\this_ppu.un1_M_current_q_cry_1 ));
    InMux I__948 (
            .O(N__9527),
            .I(\this_ppu.un1_M_current_q_cry_2 ));
    InMux I__947 (
            .O(N__9524),
            .I(\this_ppu.un1_M_current_q_cry_3 ));
    InMux I__946 (
            .O(N__9521),
            .I(\this_ppu.un1_M_current_q_cry_4 ));
    InMux I__945 (
            .O(N__9518),
            .I(\this_ppu.un1_M_current_q_cry_5 ));
    SRMux I__944 (
            .O(N__9515),
            .I(N__9512));
    LocalMux I__943 (
            .O(N__9512),
            .I(N__9509));
    Odrv12 I__942 (
            .O(N__9509),
            .I(\this_ppu.N_256_1_i ));
    InMux I__941 (
            .O(N__9506),
            .I(N__9501));
    InMux I__940 (
            .O(N__9505),
            .I(N__9496));
    InMux I__939 (
            .O(N__9504),
            .I(N__9496));
    LocalMux I__938 (
            .O(N__9501),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0 ));
    LocalMux I__937 (
            .O(N__9496),
            .I(\this_vga_signals.mult1_un68_sum_axb1_0 ));
    CascadeMux I__936 (
            .O(N__9491),
            .I(N__9488));
    InMux I__935 (
            .O(N__9488),
            .I(N__9485));
    LocalMux I__934 (
            .O(N__9485),
            .I(N__9482));
    Odrv4 I__933 (
            .O(N__9482),
            .I(M_this_vga_signals_address_10));
    CascadeMux I__932 (
            .O(N__9479),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0_cascade_));
    InMux I__931 (
            .O(N__9476),
            .I(N__9470));
    InMux I__930 (
            .O(N__9475),
            .I(N__9470));
    LocalMux I__929 (
            .O(N__9470),
            .I(\this_ppu.N_277 ));
    CascadeMux I__928 (
            .O(N__9467),
            .I(\this_ppu.M_mZ0Z1_cascade_ ));
    IoInMux I__927 (
            .O(N__9464),
            .I(N__9461));
    LocalMux I__926 (
            .O(N__9461),
            .I(N__9458));
    IoSpan4Mux I__925 (
            .O(N__9458),
            .I(N__9455));
    IoSpan4Mux I__924 (
            .O(N__9455),
            .I(N__9452));
    Span4Mux_s3_v I__923 (
            .O(N__9452),
            .I(N__9449));
    Sp12to4 I__922 (
            .O(N__9449),
            .I(N__9446));
    Odrv12 I__921 (
            .O(N__9446),
            .I(N_92));
    CascadeMux I__920 (
            .O(N__9443),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_cascade_));
    InMux I__919 (
            .O(N__9440),
            .I(N__9437));
    LocalMux I__918 (
            .O(N__9437),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0));
    InMux I__917 (
            .O(N__9434),
            .I(N__9431));
    LocalMux I__916 (
            .O(N__9431),
            .I(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1));
    CascadeMux I__915 (
            .O(N__9428),
            .I(\this_ppu.M_N_16_1_cascade_ ));
    InMux I__914 (
            .O(N__9425),
            .I(N__9422));
    LocalMux I__913 (
            .O(N__9422),
            .I(N__9418));
    InMux I__912 (
            .O(N__9421),
            .I(N__9415));
    Odrv4 I__911 (
            .O(N__9418),
            .I(\this_ppu.M_m9_i_x3Z0Z_0 ));
    LocalMux I__910 (
            .O(N__9415),
            .I(\this_ppu.M_m9_i_x3Z0Z_0 ));
    InMux I__909 (
            .O(N__9410),
            .I(N__9407));
    LocalMux I__908 (
            .O(N__9407),
            .I(\this_ppu.M_mZ0Z1 ));
    CascadeMux I__907 (
            .O(N__9404),
            .I(\this_ppu.M_m1_e_0_1_0_cascade_ ));
    InMux I__906 (
            .O(N__9401),
            .I(N__9398));
    LocalMux I__905 (
            .O(N__9398),
            .I(\this_ppu.M_m1_e_0_1_1 ));
    InMux I__904 (
            .O(N__9395),
            .I(N__9389));
    InMux I__903 (
            .O(N__9394),
            .I(N__9389));
    LocalMux I__902 (
            .O(N__9389),
            .I(\this_ppu.M_m12_0_x3_out_0 ));
    InMux I__901 (
            .O(N__9386),
            .I(N__9383));
    LocalMux I__900 (
            .O(N__9383),
            .I(\this_ppu.M_N_16_1 ));
    InMux I__899 (
            .O(N__9380),
            .I(N__9377));
    LocalMux I__898 (
            .O(N__9377),
            .I(\this_ppu.M_m1_e_0_0 ));
    CascadeMux I__897 (
            .O(N__9374),
            .I(\this_ppu.M_N_6_0_cascade_ ));
    InMux I__896 (
            .O(N__9371),
            .I(N__9368));
    LocalMux I__895 (
            .O(N__9368),
            .I(\this_ppu.M_N_13_mux ));
    InMux I__894 (
            .O(N__9365),
            .I(N__9362));
    LocalMux I__893 (
            .O(N__9362),
            .I(\this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_0 ));
    CascadeMux I__892 (
            .O(N__9359),
            .I(\this_ppu.M_N_15_mux_cascade_ ));
    CascadeMux I__891 (
            .O(N__9356),
            .I(\this_ppu.M_m12_0_x3_s_0_1Z0Z_0_cascade_ ));
    CascadeMux I__890 (
            .O(N__9353),
            .I(\this_ppu.M_m12_0_x3_out_0_cascade_ ));
    CascadeMux I__889 (
            .O(N__9350),
            .I(\this_vga_signals.if_m12_cascade_ ));
    CascadeMux I__888 (
            .O(N__9347),
            .I(N__9344));
    InMux I__887 (
            .O(N__9344),
            .I(N__9341));
    LocalMux I__886 (
            .O(N__9341),
            .I(\this_vga_signals.mult1_un54_sum_cry_1_s ));
    InMux I__885 (
            .O(N__9338),
            .I(\this_vga_signals.mult1_un54_sum_cry_0 ));
    InMux I__884 (
            .O(N__9335),
            .I(N__9332));
    LocalMux I__883 (
            .O(N__9332),
            .I(N__9329));
    Odrv12 I__882 (
            .O(N__9329),
            .I(\this_vga_signals.mult1_un47_sum_cry_1_s ));
    InMux I__881 (
            .O(N__9326),
            .I(N__9323));
    LocalMux I__880 (
            .O(N__9323),
            .I(\this_vga_signals.mult1_un61_sum_axb_3 ));
    InMux I__879 (
            .O(N__9320),
            .I(\this_vga_signals.mult1_un54_sum_cry_1 ));
    InMux I__878 (
            .O(N__9317),
            .I(N__9314));
    LocalMux I__877 (
            .O(N__9314),
            .I(N__9311));
    Odrv4 I__876 (
            .O(N__9311),
            .I(\this_vga_signals.mult1_un54_sum_axb_3 ));
    InMux I__875 (
            .O(N__9308),
            .I(\this_vga_signals.mult1_un54_sum_cry_2 ));
    CascadeMux I__874 (
            .O(N__9305),
            .I(N__9302));
    InMux I__873 (
            .O(N__9302),
            .I(N__9295));
    InMux I__872 (
            .O(N__9301),
            .I(N__9295));
    InMux I__871 (
            .O(N__9300),
            .I(N__9292));
    LocalMux I__870 (
            .O(N__9295),
            .I(\this_vga_signals.mult1_un54_sum_s_3 ));
    LocalMux I__869 (
            .O(N__9292),
            .I(\this_vga_signals.mult1_un54_sum_s_3 ));
    InMux I__868 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__867 (
            .O(N__9284),
            .I(N__9281));
    Span4Mux_v I__866 (
            .O(N__9281),
            .I(N__9278));
    Odrv4 I__865 (
            .O(N__9278),
            .I(\this_vga_signals.M_hcounter_q_i_0_5 ));
    CascadeMux I__864 (
            .O(N__9275),
            .I(N__9272));
    InMux I__863 (
            .O(N__9272),
            .I(N__9266));
    InMux I__862 (
            .O(N__9271),
            .I(N__9266));
    LocalMux I__861 (
            .O(N__9266),
            .I(N__9262));
    InMux I__860 (
            .O(N__9265),
            .I(N__9259));
    Odrv12 I__859 (
            .O(N__9262),
            .I(\this_vga_signals.mult1_un47_sum_s_3 ));
    LocalMux I__858 (
            .O(N__9259),
            .I(\this_vga_signals.mult1_un47_sum_s_3 ));
    CascadeMux I__857 (
            .O(N__9254),
            .I(N__9251));
    InMux I__856 (
            .O(N__9251),
            .I(N__9248));
    LocalMux I__855 (
            .O(N__9248),
            .I(\this_vga_signals.mult1_un47_sum_i_3 ));
    InMux I__854 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__853 (
            .O(N__9242),
            .I(\this_vga_signals.mult1_un40_sum_axb_2 ));
    CascadeMux I__852 (
            .O(N__9239),
            .I(N__9236));
    InMux I__851 (
            .O(N__9236),
            .I(N__9233));
    LocalMux I__850 (
            .O(N__9233),
            .I(N__9230));
    Odrv4 I__849 (
            .O(N__9230),
            .I(\this_vga_signals.mult1_un40_sum_axb_1_l_fx ));
    CascadeMux I__848 (
            .O(N__9227),
            .I(N__9224));
    InMux I__847 (
            .O(N__9224),
            .I(N__9217));
    InMux I__846 (
            .O(N__9223),
            .I(N__9217));
    CascadeMux I__845 (
            .O(N__9222),
            .I(N__9214));
    LocalMux I__844 (
            .O(N__9217),
            .I(N__9211));
    InMux I__843 (
            .O(N__9214),
            .I(N__9208));
    Odrv4 I__842 (
            .O(N__9211),
            .I(\this_vga_signals.mult1_un40_sum_cry_2_THRU_CO ));
    LocalMux I__841 (
            .O(N__9208),
            .I(\this_vga_signals.mult1_un40_sum_cry_2_THRU_CO ));
    CascadeMux I__840 (
            .O(N__9203),
            .I(N__9200));
    InMux I__839 (
            .O(N__9200),
            .I(N__9197));
    LocalMux I__838 (
            .O(N__9197),
            .I(\this_vga_signals.mult1_un40_sum_s_3 ));
    InMux I__837 (
            .O(N__9194),
            .I(\this_vga_signals.mult1_un61_sum_cry_0 ));
    InMux I__836 (
            .O(N__9191),
            .I(\this_vga_signals.mult1_un61_sum_cry_1 ));
    InMux I__835 (
            .O(N__9188),
            .I(\this_vga_signals.mult1_un61_sum_cry_2 ));
    InMux I__834 (
            .O(N__9185),
            .I(N__9181));
    InMux I__833 (
            .O(N__9184),
            .I(N__9178));
    LocalMux I__832 (
            .O(N__9181),
            .I(N__9172));
    LocalMux I__831 (
            .O(N__9178),
            .I(N__9172));
    InMux I__830 (
            .O(N__9177),
            .I(N__9169));
    Odrv4 I__829 (
            .O(N__9172),
            .I(\this_vga_signals.N_70_0 ));
    LocalMux I__828 (
            .O(N__9169),
            .I(\this_vga_signals.N_70_0 ));
    InMux I__827 (
            .O(N__9164),
            .I(N__9161));
    LocalMux I__826 (
            .O(N__9161),
            .I(\this_vga_signals.mult1_un54_sum_i_3 ));
    CascadeMux I__825 (
            .O(N__9158),
            .I(N_70_cascade_));
    InMux I__824 (
            .O(N__9155),
            .I(N__9152));
    LocalMux I__823 (
            .O(N__9152),
            .I(\this_vga_signals.mult1_un40_sum_cry_1_THRU_CO ));
    CascadeMux I__822 (
            .O(N__9149),
            .I(N__9146));
    InMux I__821 (
            .O(N__9146),
            .I(N__9141));
    InMux I__820 (
            .O(N__9145),
            .I(N__9136));
    InMux I__819 (
            .O(N__9144),
            .I(N__9136));
    LocalMux I__818 (
            .O(N__9141),
            .I(G_501));
    LocalMux I__817 (
            .O(N__9136),
            .I(G_501));
    InMux I__816 (
            .O(N__9131),
            .I(N__9126));
    InMux I__815 (
            .O(N__9130),
            .I(N__9121));
    InMux I__814 (
            .O(N__9129),
            .I(N__9121));
    LocalMux I__813 (
            .O(N__9126),
            .I(N_70));
    LocalMux I__812 (
            .O(N__9121),
            .I(N_70));
    CEMux I__811 (
            .O(N__9116),
            .I(N__9113));
    LocalMux I__810 (
            .O(N__9113),
            .I(N__9110));
    Span4Mux_v I__809 (
            .O(N__9110),
            .I(N__9107));
    Odrv4 I__808 (
            .O(N__9107),
            .I(N_26));
    InMux I__807 (
            .O(N__9104),
            .I(\this_vga_signals.mult1_un47_sum_cry_0 ));
    InMux I__806 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__805 (
            .O(N__9098),
            .I(N__9095));
    Odrv4 I__804 (
            .O(N__9095),
            .I(\this_vga_signals.mult1_un40_sum_cry_1_s ));
    InMux I__803 (
            .O(N__9092),
            .I(\this_vga_signals.mult1_un47_sum_cry_1 ));
    InMux I__802 (
            .O(N__9089),
            .I(N__9086));
    LocalMux I__801 (
            .O(N__9086),
            .I(\this_vga_signals.mult1_un47_sum_axb_3 ));
    InMux I__800 (
            .O(N__9083),
            .I(\this_vga_signals.mult1_un47_sum_cry_2 ));
    InMux I__799 (
            .O(N__9080),
            .I(N__9074));
    InMux I__798 (
            .O(N__9079),
            .I(N__9074));
    LocalMux I__797 (
            .O(N__9074),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1 ));
    InMux I__796 (
            .O(N__9071),
            .I(N__9068));
    LocalMux I__795 (
            .O(N__9068),
            .I(\this_vga_signals.g2_0_x1 ));
    CascadeMux I__794 (
            .O(N__9065),
            .I(\this_vga_signals.g2_0_x0_cascade_ ));
    InMux I__793 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__792 (
            .O(N__9059),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0 ));
    InMux I__791 (
            .O(N__9056),
            .I(N__9053));
    LocalMux I__790 (
            .O(N__9053),
            .I(\this_vga_signals.g2_0 ));
    CascadeMux I__789 (
            .O(N__9050),
            .I(N__9047));
    InMux I__788 (
            .O(N__9047),
            .I(N__9044));
    LocalMux I__787 (
            .O(N__9044),
            .I(N__9041));
    Odrv4 I__786 (
            .O(N__9041),
            .I(M_this_vga_signals_address_12));
    InMux I__785 (
            .O(N__9038),
            .I(N__9035));
    LocalMux I__784 (
            .O(N__9035),
            .I(\this_vga_signals.g0_2 ));
    CascadeMux I__783 (
            .O(N__9032),
            .I(N__9029));
    InMux I__782 (
            .O(N__9029),
            .I(N__9026));
    LocalMux I__781 (
            .O(N__9026),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_1 ));
    InMux I__780 (
            .O(N__9023),
            .I(\this_vga_signals.mult1_un40_sum_cry_0 ));
    InMux I__779 (
            .O(N__9020),
            .I(\this_vga_signals.mult1_un40_sum_cry_1 ));
    InMux I__778 (
            .O(N__9017),
            .I(\this_vga_signals.mult1_un40_sum_cry_2 ));
    CascadeMux I__777 (
            .O(N__9014),
            .I(\this_vga_signals.if_N_6_mux_0_0_cascade_ ));
    CascadeMux I__776 (
            .O(N__9011),
            .I(N__9008));
    InMux I__775 (
            .O(N__9008),
            .I(N__9005));
    LocalMux I__774 (
            .O(N__9005),
            .I(M_this_vga_signals_address_8));
    CascadeMux I__773 (
            .O(N__9002),
            .I(N__8999));
    InMux I__772 (
            .O(N__8999),
            .I(N__8996));
    LocalMux I__771 (
            .O(N__8996),
            .I(M_this_vga_signals_address_11));
    InMux I__770 (
            .O(N__8993),
            .I(N__8990));
    LocalMux I__769 (
            .O(N__8990),
            .I(\this_vga_signals.g0_0_a2_1 ));
    CascadeMux I__768 (
            .O(N__8987),
            .I(N__8984));
    InMux I__767 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__766 (
            .O(N__8981),
            .I(M_this_vga_signals_address_9));
    CascadeMux I__765 (
            .O(N__8978),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_cascade_ ));
    InMux I__764 (
            .O(N__8975),
            .I(N__8972));
    LocalMux I__763 (
            .O(N__8972),
            .I(\this_vga_ramdac.m16 ));
    IoInMux I__762 (
            .O(N__8969),
            .I(N__8966));
    LocalMux I__761 (
            .O(N__8966),
            .I(N__8963));
    IoSpan4Mux I__760 (
            .O(N__8963),
            .I(N__8960));
    IoSpan4Mux I__759 (
            .O(N__8960),
            .I(N__8957));
    Span4Mux_s2_h I__758 (
            .O(N__8957),
            .I(N__8954));
    Odrv4 I__757 (
            .O(N__8954),
            .I(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_2 ));
    InMux I__756 (
            .O(N__8951),
            .I(N__8948));
    LocalMux I__755 (
            .O(N__8948),
            .I(\this_vga_ramdac.m19 ));
    IoInMux I__754 (
            .O(N__8945),
            .I(N__8942));
    LocalMux I__753 (
            .O(N__8942),
            .I(N__8939));
    Span4Mux_s2_h I__752 (
            .O(N__8939),
            .I(N__8936));
    Sp12to4 I__751 (
            .O(N__8936),
            .I(N__8933));
    Span12Mux_v I__750 (
            .O(N__8933),
            .I(N__8930));
    Odrv12 I__749 (
            .O(N__8930),
            .I(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_3 ));
    IoInMux I__748 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__747 (
            .O(N__8924),
            .I(N__8921));
    Span4Mux_s2_h I__746 (
            .O(N__8921),
            .I(N__8918));
    Odrv4 I__745 (
            .O(N__8918),
            .I(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_1 ));
    InMux I__744 (
            .O(N__8915),
            .I(N__8912));
    LocalMux I__743 (
            .O(N__8912),
            .I(\this_vga_ramdac.i2_mux ));
    InMux I__742 (
            .O(N__8909),
            .I(N__8906));
    LocalMux I__741 (
            .O(N__8906),
            .I(N__8900));
    InMux I__740 (
            .O(N__8905),
            .I(N__8897));
    InMux I__739 (
            .O(N__8904),
            .I(N__8892));
    InMux I__738 (
            .O(N__8903),
            .I(N__8892));
    Span4Mux_s3_h I__737 (
            .O(N__8900),
            .I(N__8885));
    LocalMux I__736 (
            .O(N__8897),
            .I(N__8885));
    LocalMux I__735 (
            .O(N__8892),
            .I(N__8882));
    InMux I__734 (
            .O(N__8891),
            .I(N__8877));
    InMux I__733 (
            .O(N__8890),
            .I(N__8877));
    Span4Mux_v I__732 (
            .O(N__8885),
            .I(N__8870));
    Span4Mux_s3_h I__731 (
            .O(N__8882),
            .I(N__8870));
    LocalMux I__730 (
            .O(N__8877),
            .I(N__8870));
    Span4Mux_h I__729 (
            .O(N__8870),
            .I(N__8867));
    Odrv4 I__728 (
            .O(N__8867),
            .I(M_this_vram_read_data_0));
    InMux I__727 (
            .O(N__8864),
            .I(N__8856));
    InMux I__726 (
            .O(N__8863),
            .I(N__8856));
    InMux I__725 (
            .O(N__8862),
            .I(N__8851));
    InMux I__724 (
            .O(N__8861),
            .I(N__8851));
    LocalMux I__723 (
            .O(N__8856),
            .I(N__8846));
    LocalMux I__722 (
            .O(N__8851),
            .I(N__8843));
    InMux I__721 (
            .O(N__8850),
            .I(N__8838));
    InMux I__720 (
            .O(N__8849),
            .I(N__8838));
    Span4Mux_v I__719 (
            .O(N__8846),
            .I(N__8835));
    Span4Mux_s3_h I__718 (
            .O(N__8843),
            .I(N__8830));
    LocalMux I__717 (
            .O(N__8838),
            .I(N__8830));
    Span4Mux_h I__716 (
            .O(N__8835),
            .I(N__8825));
    Span4Mux_h I__715 (
            .O(N__8830),
            .I(N__8825));
    Odrv4 I__714 (
            .O(N__8825),
            .I(M_this_vram_read_data_2));
    InMux I__713 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__712 (
            .O(N__8819),
            .I(N__8812));
    InMux I__711 (
            .O(N__8818),
            .I(N__8809));
    CascadeMux I__710 (
            .O(N__8817),
            .I(N__8805));
    InMux I__709 (
            .O(N__8816),
            .I(N__8800));
    InMux I__708 (
            .O(N__8815),
            .I(N__8800));
    Span4Mux_s3_h I__707 (
            .O(N__8812),
            .I(N__8795));
    LocalMux I__706 (
            .O(N__8809),
            .I(N__8795));
    InMux I__705 (
            .O(N__8808),
            .I(N__8790));
    InMux I__704 (
            .O(N__8805),
            .I(N__8790));
    LocalMux I__703 (
            .O(N__8800),
            .I(N__8787));
    Span4Mux_v I__702 (
            .O(N__8795),
            .I(N__8784));
    LocalMux I__701 (
            .O(N__8790),
            .I(N__8779));
    Span4Mux_s3_h I__700 (
            .O(N__8787),
            .I(N__8779));
    Span4Mux_h I__699 (
            .O(N__8784),
            .I(N__8774));
    Span4Mux_h I__698 (
            .O(N__8779),
            .I(N__8774));
    Odrv4 I__697 (
            .O(N__8774),
            .I(M_this_vram_read_data_1));
    CascadeMux I__696 (
            .O(N__8771),
            .I(N__8768));
    InMux I__695 (
            .O(N__8768),
            .I(N__8763));
    CascadeMux I__694 (
            .O(N__8767),
            .I(N__8759));
    CascadeMux I__693 (
            .O(N__8766),
            .I(N__8756));
    LocalMux I__692 (
            .O(N__8763),
            .I(N__8752));
    InMux I__691 (
            .O(N__8762),
            .I(N__8749));
    InMux I__690 (
            .O(N__8759),
            .I(N__8744));
    InMux I__689 (
            .O(N__8756),
            .I(N__8744));
    CascadeMux I__688 (
            .O(N__8755),
            .I(N__8740));
    Span4Mux_s3_h I__687 (
            .O(N__8752),
            .I(N__8735));
    LocalMux I__686 (
            .O(N__8749),
            .I(N__8735));
    LocalMux I__685 (
            .O(N__8744),
            .I(N__8732));
    InMux I__684 (
            .O(N__8743),
            .I(N__8727));
    InMux I__683 (
            .O(N__8740),
            .I(N__8727));
    Span4Mux_v I__682 (
            .O(N__8735),
            .I(N__8720));
    Span4Mux_s3_h I__681 (
            .O(N__8732),
            .I(N__8720));
    LocalMux I__680 (
            .O(N__8727),
            .I(N__8720));
    Span4Mux_h I__679 (
            .O(N__8720),
            .I(N__8717));
    Odrv4 I__678 (
            .O(N__8717),
            .I(M_this_vram_read_data_3));
    InMux I__677 (
            .O(N__8714),
            .I(N__8711));
    LocalMux I__676 (
            .O(N__8711),
            .I(N__8708));
    Span4Mux_s3_h I__675 (
            .O(N__8708),
            .I(N__8700));
    InMux I__674 (
            .O(N__8707),
            .I(N__8697));
    InMux I__673 (
            .O(N__8706),
            .I(N__8690));
    InMux I__672 (
            .O(N__8705),
            .I(N__8690));
    InMux I__671 (
            .O(N__8704),
            .I(N__8690));
    InMux I__670 (
            .O(N__8703),
            .I(N__8687));
    Odrv4 I__669 (
            .O(N__8700),
            .I(\this_vga_ramdac.N_706_0 ));
    LocalMux I__668 (
            .O(N__8697),
            .I(\this_vga_ramdac.N_706_0 ));
    LocalMux I__667 (
            .O(N__8690),
            .I(\this_vga_ramdac.N_706_0 ));
    LocalMux I__666 (
            .O(N__8687),
            .I(\this_vga_ramdac.N_706_0 ));
    InMux I__665 (
            .O(N__8678),
            .I(N__8675));
    LocalMux I__664 (
            .O(N__8675),
            .I(\this_vga_ramdac.i2_mux_0 ));
    IoInMux I__663 (
            .O(N__8672),
            .I(N__8669));
    LocalMux I__662 (
            .O(N__8669),
            .I(N__8666));
    IoSpan4Mux I__661 (
            .O(N__8666),
            .I(N__8663));
    IoSpan4Mux I__660 (
            .O(N__8663),
            .I(N__8660));
    IoSpan4Mux I__659 (
            .O(N__8660),
            .I(N__8657));
    Span4Mux_s3_h I__658 (
            .O(N__8657),
            .I(N__8654));
    Odrv4 I__657 (
            .O(N__8654),
            .I(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_4 ));
    IoInMux I__656 (
            .O(N__8651),
            .I(N__8648));
    LocalMux I__655 (
            .O(N__8648),
            .I(N__8645));
    Span4Mux_s2_h I__654 (
            .O(N__8645),
            .I(N__8642));
    Span4Mux_h I__653 (
            .O(N__8642),
            .I(N__8639));
    Odrv4 I__652 (
            .O(N__8639),
            .I(N_94));
    IoInMux I__651 (
            .O(N__8636),
            .I(N__8633));
    LocalMux I__650 (
            .O(N__8633),
            .I(N__8630));
    Span4Mux_s3_v I__649 (
            .O(N__8630),
            .I(N__8627));
    Span4Mux_v I__648 (
            .O(N__8627),
            .I(N__8624));
    Span4Mux_v I__647 (
            .O(N__8624),
            .I(N__8621));
    Span4Mux_v I__646 (
            .O(N__8621),
            .I(N__8618));
    Odrv4 I__645 (
            .O(N__8618),
            .I(N_274_i));
    IoInMux I__644 (
            .O(N__8615),
            .I(N__8612));
    LocalMux I__643 (
            .O(N__8612),
            .I(\this_vga_signals.N_517_1 ));
    IoInMux I__642 (
            .O(N__8609),
            .I(N__8606));
    LocalMux I__641 (
            .O(N__8606),
            .I(N_205_i));
    IoInMux I__640 (
            .O(N__8603),
            .I(N__8600));
    LocalMux I__639 (
            .O(N__8600),
            .I(N__8597));
    IoSpan4Mux I__638 (
            .O(N__8597),
            .I(N__8594));
    Span4Mux_s0_h I__637 (
            .O(N__8594),
            .I(N__8591));
    Odrv4 I__636 (
            .O(N__8591),
            .I(\this_vga_ramdac.M_this_rgb_d_3_0_dreg ));
    CascadeMux I__635 (
            .O(N__8588),
            .I(\this_vga_ramdac.m5_cascade_ ));
    IoInMux I__634 (
            .O(N__8585),
            .I(N__8582));
    LocalMux I__633 (
            .O(N__8582),
            .I(N__8579));
    IoSpan4Mux I__632 (
            .O(N__8579),
            .I(N__8576));
    Span4Mux_s2_h I__631 (
            .O(N__8576),
            .I(N__8573));
    Odrv4 I__630 (
            .O(N__8573),
            .I(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_0 ));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_1_cry_8 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(un1_M_this_internal_address_q_cry_7),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_31_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_31_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_31_23_0_));
    defparam IN_MUX_bfv_31_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_31_24_0_ (
            .carryinitin(un1_M_this_external_address_q_cry_7),
            .carryinitout(bfn_31_24_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(un1_M_this_data_count_q_cry_7),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO),
            .carryinitout(bfn_15_25_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIIRV75_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__16529),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_684_g ));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI6RKH5_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__8615),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_517_1_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_3  (
            .USERSIGNALTOGLOBALBUFFER(N__19594),
            .GLOBALBUFFEROUTPUT(M_this_state_q_nss_g_0));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6RKH5_9_LC_1_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6RKH5_9_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6RKH5_9_LC_1_17_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI6RKH5_9_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__17143),
            .in2(_gnd_net_),
            .in3(N__15497),
            .lcout(\this_vga_signals.N_517_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_205_i_LC_1_22_1 .C_ON=1'b0;
    defparam \this_vga_signals.N_205_i_LC_1_22_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_205_i_LC_1_22_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_vga_signals.N_205_i_LC_1_22_1  (
            .in0(N__20214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20641),
            .lcout(N_205_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_0_LC_3_9_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_0_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_0_LC_3_9_4 .LUT_INIT=16'b0001110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_0_LC_3_9_4  (
            .in0(N__8822),
            .in1(N__8909),
            .in2(N__8771),
            .in3(N__8714),
            .lcout(\this_vga_ramdac.M_this_rgb_d_3_0_dreg ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m5_LC_3_12_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m5_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m5_LC_3_12_6 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m5_LC_3_12_6  (
            .in0(N__8863),
            .in1(N__8818),
            .in2(_gnd_net_),
            .in3(N__8905),
            .lcout(),
            .ltout(\this_vga_ramdac.m5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_1_LC_3_12_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_1_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_1_LC_3_12_7 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_1_LC_3_12_7  (
            .in0(N__8762),
            .in1(N__8864),
            .in2(N__8588),
            .in3(N__8707),
            .lcout(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_3_13_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_3_13_0 .LUT_INIT=16'b0010001110010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_3_13_0  (
            .in0(N__8861),
            .in1(N__8816),
            .in2(N__8766),
            .in3(N__8903),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_3_13_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_3_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_3_13_6 .LUT_INIT=16'b0110010100101011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_3_13_6  (
            .in0(N__8862),
            .in1(N__8815),
            .in2(N__8767),
            .in3(N__8904),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_3_LC_3_14_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_3_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_3_LC_3_14_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_3_LC_3_14_2  (
            .in0(N__8975),
            .in1(N__8705),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_4_LC_3_14_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_4_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_4_LC_3_14_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_4_LC_3_14_5  (
            .in0(N__8706),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8951),
            .lcout(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_2_LC_3_14_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_2_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_2_LC_3_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_2_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__8704),
            .in2(_gnd_net_),
            .in3(N__8915),
            .lcout(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_4_13_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_4_13_0 .LUT_INIT=16'b0001010100111101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_4_13_0  (
            .in0(N__8849),
            .in1(N__8808),
            .in2(N__8755),
            .in3(N__8890),
            .lcout(\this_vga_ramdac.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_250_LC_4_13_1 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_250_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_q_250_LC_4_13_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_250_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__23823),
            .in2(_gnd_net_),
            .in3(N__24787),
            .lcout(\this_vga_ramdac.N_706_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_13_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_13_5 .LUT_INIT=16'b0010010000111011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_4_13_5  (
            .in0(N__8891),
            .in1(N__8850),
            .in2(N__8817),
            .in3(N__8743),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_5_LC_4_14_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_5_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_5_LC_4_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNO_5_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__8703),
            .in2(_gnd_net_),
            .in3(N__8678),
            .lcout(\this_vga_ramdac.M_this_rgb_d_3_0_dregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNID8NA3_9_LC_7_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNID8NA3_9_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNID8NA3_9_LC_7_13_7 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNID8NA3_9_LC_7_13_7  (
            .in0(N__20218),
            .in1(N__9872),
            .in2(N__13485),
            .in3(N__16642),
            .lcout(N_94),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJVML2_9_LC_7_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJVML2_9_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIJVML2_9_LC_7_17_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIJVML2_9_LC_7_17_7  (
            .in0(N__16643),
            .in1(N__9868),
            .in2(_gnd_net_),
            .in3(N__13486),
            .lcout(N_274_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_9_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_9_9_0 .LUT_INIT=16'b1111101000110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_9_9_0  (
            .in0(N__9506),
            .in1(N__9629),
            .in2(N__14132),
            .in3(N__14572),
            .lcout(),
            .ltout(\this_vga_signals.if_N_6_mux_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNINGUT4R3_7_LC_9_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNINGUT4R3_7_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNINGUT4R3_7_LC_9_9_1 .LUT_INIT=16'b1000001000100010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNINGUT4R3_7_LC_9_9_1  (
            .in0(N__23853),
            .in1(N__8993),
            .in2(N__9014),
            .in3(N__9056),
            .lcout(M_this_vga_signals_address_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI6UL1Q3_7_LC_9_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI6UL1Q3_7_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI6UL1Q3_7_LC_9_9_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI6UL1Q3_7_LC_9_9_3  (
            .in0(N__23852),
            .in1(N__12095),
            .in2(_gnd_net_),
            .in3(N__12200),
            .lcout(M_this_vga_signals_address_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_a2_1_LC_9_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_a2_1_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_a2_1_LC_9_9_5 .LUT_INIT=16'b0001011111101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_a2_1_LC_9_9_5  (
            .in0(N__9584),
            .in1(N__14376),
            .in2(N__14582),
            .in3(N__9667),
            .lcout(\this_vga_signals.g0_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_LC_9_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_x2_LC_9_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_x2_LC_9_9_6  (
            .in0(N__13987),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14122),
            .lcout(\this_vga_signals.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIR4HAL91_7_LC_9_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIR4HAL91_7_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIR4HAL91_7_LC_9_10_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIR4HAL91_7_LC_9_10_0  (
            .in0(N__23851),
            .in1(N__9596),
            .in2(_gnd_net_),
            .in3(N__9080),
            .lcout(M_this_vga_signals_address_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_9_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_9_10_1 .LUT_INIT=16'b0001101001111010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_LC_9_10_1  (
            .in0(N__14375),
            .in1(N__9583),
            .in2(N__9668),
            .in3(N__14565),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_N_3_i_LC_9_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_N_3_i_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_N_3_i_LC_9_10_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_N_3_i_LC_9_10_3  (
            .in0(N__9038),
            .in1(N__11285),
            .in2(N__9032),
            .in3(N__12377),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_x1_LC_9_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_x1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_x1_LC_9_10_4 .LUT_INIT=16'b0010110101111000;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_x1_LC_9_10_4  (
            .in0(N__14564),
            .in1(N__9504),
            .in2(N__8978),
            .in3(N__9624),
            .lcout(\this_vga_signals.g2_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_5_LC_9_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_5_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_5_LC_9_10_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_5_LC_9_10_5  (
            .in0(N__15135),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12567),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_x0_LC_9_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_x0_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_x0_LC_9_10_6 .LUT_INIT=16'b1100101000110101;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_x0_LC_9_10_6  (
            .in0(N__9625),
            .in1(N__9505),
            .in2(N__14581),
            .in3(N__9079),
            .lcout(),
            .ltout(\this_vga_signals.g2_0_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_ns_LC_9_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_ns_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_ns_LC_9_10_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_ns_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__9071),
            .in2(N__9065),
            .in3(N__9062),
            .lcout(\this_vga_signals.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNINSNSM_7_LC_9_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNINSNSM_7_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNINSNSM_7_LC_9_11_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNINSNSM_7_LC_9_11_1  (
            .in0(N__12569),
            .in1(N__23860),
            .in2(_gnd_net_),
            .in3(N__12644),
            .lcout(M_this_vga_signals_address_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_9_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_9_11_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_9_11_4  (
            .in0(N__12089),
            .in1(N__12568),
            .in2(N__15155),
            .in3(N__12194),
            .lcout(\this_vga_signals.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_9_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_9_11_5 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_0_LC_9_11_5  (
            .in0(N__12193),
            .in1(N__14377),
            .in2(N__15449),
            .in3(N__12090),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_0_c_LC_9_12_0 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_0_c_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_0_c_LC_9_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_0_c_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__16343),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\this_vga_signals.mult1_un40_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_1_s_LC_9_12_1 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_1_s_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_1_s_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_1_s_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__9185),
            .in2(N__9239),
            .in3(N__9023),
            .lcout(\this_vga_signals.mult1_un40_sum_cry_1_s ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un40_sum_cry_0 ),
            .carryout(\this_vga_signals.mult1_un40_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.mult1_un40_sum_cry_1_THRU_LUT4_0_LC_9_12_2 .C_ON=1'b1;
    defparam \this_vga_signals.mult1_un40_sum_cry_1_THRU_LUT4_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.mult1_un40_sum_cry_1_THRU_LUT4_0_LC_9_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.mult1_un40_sum_cry_1_THRU_LUT4_0_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__9131),
            .in2(N__9149),
            .in3(N__9020),
            .lcout(\this_vga_signals.mult1_un40_sum_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un40_sum_cry_1 ),
            .carryout(\this_vga_signals.mult1_un40_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.mult1_un40_sum_cry_2_THRU_LUT4_0_LC_9_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.mult1_un40_sum_cry_2_THRU_LUT4_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.mult1_un40_sum_cry_2_THRU_LUT4_0_LC_9_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.mult1_un40_sum_cry_2_THRU_LUT4_0_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9017),
            .lcout(\this_vga_signals.mult1_un40_sum_cry_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_2_c_inv_LC_9_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_2_c_inv_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_2_c_inv_LC_9_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_cry_2_c_inv_LC_9_13_0  (
            .in0(N__9184),
            .in1(N__9144),
            .in2(_gnd_net_),
            .in3(N__9129),
            .lcout(N_70),
            .ltout(N_70_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_l_fx_LC_9_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_l_fx_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_l_fx_LC_9_13_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_l_fx_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9158),
            .in3(N__9245),
            .lcout(G_501),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_axb_3_LC_9_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_axb_3_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_axb_3_LC_9_13_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_axb_3_LC_9_13_4  (
            .in0(N__9155),
            .in1(N__9145),
            .in2(N__9222),
            .in3(N__9130),
            .lcout(\this_vga_signals.mult1_un47_sum_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_vram_write_en_i_0_i_0_LC_9_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_vram_write_en_i_0_i_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_vram_write_en_i_0_i_0_LC_9_13_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_this_vram_write_en_i_0_i_0_LC_9_13_7  (
            .in0(N__22385),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23552),
            .lcout(N_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_0_c_LC_9_14_0 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_0_c_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_0_c_LC_9_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_0_c_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__16220),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\this_vga_signals.mult1_un47_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_1_s_LC_9_14_1 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_1_s_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_1_s_LC_9_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_cry_1_s_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__9287),
            .in2(N__9203),
            .in3(N__9104),
            .lcout(\this_vga_signals.mult1_un47_sum_cry_1_s ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un47_sum_cry_0 ),
            .carryout(\this_vga_signals.mult1_un47_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_axb_3_LC_9_14_2 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_axb_3_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_axb_3_LC_9_14_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_axb_3_LC_9_14_2  (
            .in0(N__9265),
            .in1(N__9101),
            .in2(N__9227),
            .in3(N__9092),
            .lcout(\this_vga_signals.mult1_un54_sum_axb_3 ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un47_sum_cry_1 ),
            .carryout(\this_vga_signals.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_s_3_LC_9_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_s_3_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_s_3_LC_9_14_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_s_3_LC_9_14_3  (
            .in0(N__9089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9083),
            .lcout(\this_vga_signals.mult1_un47_sum_s_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_LC_9_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_LC_9_14_4 .LUT_INIT=16'b1110011110011110;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_2_LC_9_14_4  (
            .in0(N__15794),
            .in1(N__15890),
            .in2(N__16004),
            .in3(N__16101),
            .lcout(\this_vga_signals.mult1_un40_sum_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_1_l_fx_LC_9_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_1_l_fx_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_1_l_fx_LC_9_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_axb_1_l_fx_LC_9_14_6  (
            .in0(N__15793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9177),
            .lcout(\this_vga_signals.mult1_un40_sum_axb_1_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_s_3_LC_9_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_s_3_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_s_3_LC_9_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un40_sum_s_3_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9223),
            .lcout(\this_vga_signals.mult1_un40_sum_s_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_0_c_LC_9_15_0 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_0_c_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_0_c_LC_9_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_0_c_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__18106),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\this_vga_signals.mult1_un61_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_1_s_LC_9_15_1 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_1_s_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_1_s_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_cry_1_s_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__13841),
            .in2(N__9305),
            .in3(N__9194),
            .lcout(\this_vga_signals.mult1_un61_sum_cry_1_s ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un61_sum_cry_0 ),
            .carryout(\this_vga_signals.mult1_un61_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_axb_3_LC_9_15_2 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_axb_3_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_axb_3_LC_9_15_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_axb_3_LC_9_15_2  (
            .in0(N__12877),
            .in1(N__9164),
            .in2(N__9347),
            .in3(N__9191),
            .lcout(\this_vga_signals.mult1_un68_sum_axb_3 ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un61_sum_cry_1 ),
            .carryout(\this_vga_signals.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_s_3_LC_9_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_s_3_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_s_3_LC_9_15_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_s_3_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__9326),
            .in2(_gnd_net_),
            .in3(N__9188),
            .lcout(\this_vga_signals.mult1_un61_sum_s_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNITQQM_9_LC_9_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNITQQM_9_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNITQQM_9_LC_9_15_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNITQQM_9_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__16581),
            .in2(_gnd_net_),
            .in3(N__13804),
            .lcout(\this_vga_signals.CO1_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNICJJV_9_LC_9_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICJJV_9_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICJJV_9_LC_9_15_5 .LUT_INIT=16'b0111000110100111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNICJJV_9_LC_9_15_5  (
            .in0(N__15889),
            .in1(N__15792),
            .in2(N__16003),
            .in3(N__16100),
            .lcout(\this_vga_signals.N_70_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_3_LC_9_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_3_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_3_LC_9_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_3_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9301),
            .lcout(\this_vga_signals.mult1_un54_sum_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_0_c_LC_9_16_0 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_0_c_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_0_c_LC_9_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_0_c_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__17006),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\this_vga_signals.mult1_un54_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_1_s_LC_9_16_1 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_1_s_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_1_s_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_cry_1_s_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__11645),
            .in2(N__9275),
            .in3(N__9338),
            .lcout(\this_vga_signals.mult1_un54_sum_cry_1_s ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un54_sum_cry_0 ),
            .carryout(\this_vga_signals.mult1_un54_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_axb_3_LC_9_16_2 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_axb_3_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_axb_3_LC_9_16_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_axb_3_LC_9_16_2  (
            .in0(N__9300),
            .in1(N__9335),
            .in2(N__9254),
            .in3(N__9320),
            .lcout(\this_vga_signals.mult1_un61_sum_axb_3 ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un54_sum_cry_1 ),
            .carryout(\this_vga_signals.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_s_3_LC_9_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_s_3_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_s_3_LC_9_16_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_s_3_LC_9_16_3  (
            .in0(N__9317),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9308),
            .lcout(\this_vga_signals.mult1_un54_sum_s_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI54V41_5_LC_9_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI54V41_5_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI54V41_5_LC_9_16_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI54V41_5_LC_9_16_4  (
            .in0(N__14342),
            .in1(N__15423),
            .in2(_gnd_net_),
            .in3(N__15150),
            .lcout(\this_vga_signals.vsync_1_0_a2_6_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_sbtinv_5_LC_9_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_sbtinv_5_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_sbtinv_5_LC_9_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_sbtinv_5_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16338),
            .lcout(\this_vga_signals.M_hcounter_q_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_3_LC_9_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_3_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_3_LC_9_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_3_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9271),
            .lcout(\this_vga_signals.mult1_un47_sum_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m8_0_LC_9_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_m8_0_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m8_0_LC_9_17_0 .LUT_INIT=16'b0101001101010101;
    LogicCell40 \this_ppu.M_m8_0_LC_9_17_0  (
            .in0(N__9848),
            .in1(N__11849),
            .in2(N__13988),
            .in3(N__10598),
            .lcout(\this_ppu.M_N_13_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m9_i_x3_0_LC_9_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_m9_i_x3_0_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m9_i_x3_0_LC_9_17_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_ppu.M_m9_i_x3_0_LC_9_17_1  (
            .in0(N__14109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13985),
            .lcout(\this_ppu.M_m9_i_x3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_LC_9_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_LC_9_17_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_LC_9_17_4  (
            .in0(N__14498),
            .in1(N__14107),
            .in2(_gnd_net_),
            .in3(N__14335),
            .lcout(\this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m5_0_LC_9_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_m5_0_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m5_0_LC_9_17_5 .LUT_INIT=16'b0001111101010100;
    LogicCell40 \this_ppu.M_m5_0_LC_9_17_5  (
            .in0(N__10599),
            .in1(N__13981),
            .in2(N__11857),
            .in3(N__9847),
            .lcout(),
            .ltout(\this_ppu.M_N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m11_LC_9_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_m11_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m11_LC_9_17_6 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \this_ppu.M_m11_LC_9_17_6  (
            .in0(N__14144),
            .in1(N__14108),
            .in2(N__9374),
            .in3(N__9371),
            .lcout(),
            .ltout(\this_ppu.M_N_15_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_0_LC_9_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_0_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_0_LC_9_17_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_ppu.M_state_d_0_sqmuxa_i_0_0_o4_0_LC_9_17_7  (
            .in0(N__9365),
            .in1(N__15202),
            .in2(N__9359),
            .in3(N__15422),
            .lcout(\this_ppu.N_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m12_0_x3_s_0_1_0_LC_9_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_m12_0_x3_s_0_1_0_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m12_0_x3_s_0_1_0_LC_9_18_0 .LUT_INIT=16'b0001001011101101;
    LogicCell40 \this_ppu.M_m12_0_x3_s_0_1_0_LC_9_18_0  (
            .in0(N__14556),
            .in1(N__10499),
            .in2(N__14129),
            .in3(N__10492),
            .lcout(),
            .ltout(\this_ppu.M_m12_0_x3_s_0_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m12_0_x3_s_0_LC_9_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_m12_0_x3_s_0_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m12_0_x3_s_0_LC_9_18_1 .LUT_INIT=16'b1000011111100001;
    LogicCell40 \this_ppu.M_m12_0_x3_s_0_LC_9_18_1  (
            .in0(N__14118),
            .in1(N__14557),
            .in2(N__9356),
            .in3(N__9836),
            .lcout(\this_ppu.M_m12_0_x3_out_0 ),
            .ltout(\this_ppu.M_m12_0_x3_out_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_4_LC_9_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_4_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_4_LC_9_18_2 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \this_ppu.M_state_q_RNO_4_LC_9_18_2  (
            .in0(N__14114),
            .in1(N__13986),
            .in2(N__9353),
            .in3(N__9475),
            .lcout(\this_ppu.M_m1_e_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_m12_LC_9_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_m12_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_m12_LC_9_18_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_m12_LC_9_18_4  (
            .in0(N__15398),
            .in1(N__10518),
            .in2(_gnd_net_),
            .in3(N__10535),
            .lcout(),
            .ltout(\this_vga_signals.if_m12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_m14_0_LC_9_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_m14_0_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_m14_0_LC_9_18_5 .LUT_INIT=16'b1011101001010001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_m14_0_LC_9_18_5  (
            .in0(N__10493),
            .in1(N__14113),
            .in2(N__9350),
            .in3(N__14555),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0),
            .ltout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_c3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m1_LC_9_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_m1_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m1_LC_9_18_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_ppu.M_m1_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9479),
            .in3(N__10577),
            .lcout(\this_ppu.M_mZ0Z1 ),
            .ltout(\this_ppu.M_mZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIMJNMSC_LC_9_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIMJNMSC_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIMJNMSC_LC_9_18_7 .LUT_INIT=16'b0100000100000000;
    LogicCell40 \this_ppu.M_state_q_RNIMJNMSC_LC_9_18_7  (
            .in0(N__9476),
            .in1(N__9421),
            .in2(N__9467),
            .in3(N__10547),
            .lcout(\this_ppu.M_m1_e_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_9_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_9_19_1 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_9_19_1  (
            .in0(N__16103),
            .in1(N__15888),
            .in2(_gnd_net_),
            .in3(N__16002),
            .lcout(N_92),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_LC_9_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_LC_9_19_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_LC_9_19_2  (
            .in0(N__11858),
            .in1(N__10601),
            .in2(N__14580),
            .in3(N__9835),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1),
            .ltout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m12_0_o3_0_LC_9_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_m12_0_o3_0_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m12_0_o3_0_LC_9_19_3 .LUT_INIT=16'b0000111000001101;
    LogicCell40 \this_ppu.M_m12_0_o3_0_LC_9_19_3  (
            .in0(N__10576),
            .in1(N__14130),
            .in2(N__9443),
            .in3(N__9440),
            .lcout(\this_ppu.M_N_16_1 ),
            .ltout(\this_ppu.M_N_16_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_3_LC_9_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_3_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_3_LC_9_19_4 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \this_ppu.M_state_q_RNO_3_LC_9_19_4  (
            .in0(N__9434),
            .in1(N__9394),
            .in2(N__9428),
            .in3(N__10546),
            .lcout(),
            .ltout(\this_ppu.M_m1_e_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_2_LC_9_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_2_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_2_LC_9_19_5 .LUT_INIT=16'b1001000000000000;
    LogicCell40 \this_ppu.M_state_q_RNO_2_LC_9_19_5  (
            .in0(N__9425),
            .in1(N__9410),
            .in2(N__9404),
            .in3(N__9401),
            .lcout(\this_ppu.M_N_3_mux_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI8H768U_LC_9_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI8H768U_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI8H768U_LC_9_19_7 .LUT_INIT=16'b1111011011110000;
    LogicCell40 \this_ppu.M_state_q_RNI8H768U_LC_9_19_7  (
            .in0(N__9395),
            .in1(N__9386),
            .in2(N__24800),
            .in3(N__9380),
            .lcout(\this_ppu.N_256_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_current_q_0_LC_9_20_0 .C_ON=1'b1;
    defparam \this_ppu.M_current_q_0_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_current_q_0_LC_9_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.M_current_q_0_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__10995),
            .in2(N__22378),
            .in3(N__22386),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\this_ppu.un1_M_current_q_cry_0 ),
            .clk(N__25021),
            .ce(),
            .sr(N__9515));
    defparam \this_ppu.M_current_q_1_LC_9_20_1 .C_ON=1'b1;
    defparam \this_ppu.M_current_q_1_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_current_q_1_LC_9_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.M_current_q_1_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__10721),
            .in2(_gnd_net_),
            .in3(N__9533),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(\this_ppu.un1_M_current_q_cry_0 ),
            .carryout(\this_ppu.un1_M_current_q_cry_1 ),
            .clk(N__25021),
            .ce(),
            .sr(N__9515));
    defparam \this_ppu.M_current_q_2_LC_9_20_2 .C_ON=1'b1;
    defparam \this_ppu.M_current_q_2_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_current_q_2_LC_9_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.M_current_q_2_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__9936),
            .in2(_gnd_net_),
            .in3(N__9530),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(\this_ppu.un1_M_current_q_cry_1 ),
            .carryout(\this_ppu.un1_M_current_q_cry_2 ),
            .clk(N__25021),
            .ce(),
            .sr(N__9515));
    defparam \this_ppu.M_current_q_3_LC_9_20_3 .C_ON=1'b1;
    defparam \this_ppu.M_current_q_3_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_current_q_3_LC_9_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.M_current_q_3_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__10860),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(M_this_ppu_vram_addr_3),
            .ltout(),
            .carryin(\this_ppu.un1_M_current_q_cry_2 ),
            .carryout(\this_ppu.un1_M_current_q_cry_3 ),
            .clk(N__25021),
            .ce(),
            .sr(N__9515));
    defparam \this_ppu.M_current_q_4_LC_9_20_4 .C_ON=1'b1;
    defparam \this_ppu.M_current_q_4_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_current_q_4_LC_9_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.M_current_q_4_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__10223),
            .in2(_gnd_net_),
            .in3(N__9524),
            .lcout(M_this_ppu_vram_addr_4),
            .ltout(),
            .carryin(\this_ppu.un1_M_current_q_cry_3 ),
            .carryout(\this_ppu.un1_M_current_q_cry_4 ),
            .clk(N__25021),
            .ce(),
            .sr(N__9515));
    defparam \this_ppu.M_current_q_5_LC_9_20_5 .C_ON=1'b1;
    defparam \this_ppu.M_current_q_5_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_current_q_5_LC_9_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.M_current_q_5_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__10364),
            .in2(_gnd_net_),
            .in3(N__9521),
            .lcout(M_this_ppu_vram_addr_5),
            .ltout(),
            .carryin(\this_ppu.un1_M_current_q_cry_4 ),
            .carryout(\this_ppu.un1_M_current_q_cry_5 ),
            .clk(N__25021),
            .ce(),
            .sr(N__9515));
    defparam \this_ppu.M_current_q_6_LC_9_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_current_q_6_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_current_q_6_LC_9_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_current_q_6_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__10073),
            .in2(_gnd_net_),
            .in3(N__9518),
            .lcout(M_this_ppu_vram_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25021),
            .ce(),
            .sr(N__9515));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0_5_LC_10_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0_5_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0_5_LC_10_9_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0_5_LC_10_9_0  (
            .in0(N__12198),
            .in1(N__12466),
            .in2(N__11204),
            .in3(N__9649),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un68_sum_axb1_LC_10_9_1  (
            .in0(N__12364),
            .in1(N__11277),
            .in2(_gnd_net_),
            .in3(N__14373),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIN3CPT8_7_LC_10_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIN3CPT8_7_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIN3CPT8_7_LC_10_9_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIN3CPT8_7_LC_10_9_2  (
            .in0(N__23850),
            .in1(_gnd_net_),
            .in2(N__11288),
            .in3(N__12365),
            .lcout(M_this_vga_signals_address_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_10_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_10_9_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_LC_10_9_4  (
            .in0(N__11278),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12363),
            .lcout(\this_vga_signals.N_9_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_5_LC_10_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_5_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_5_LC_10_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIDB4TM3_5_LC_10_9_5  (
            .in0(N__12467),
            .in1(N__11200),
            .in2(N__9653),
            .in3(N__12199),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_esr_RNIDB4TM3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGU2FNB_5_LC_10_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGU2FNB_5_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGU2FNB_5_LC_10_9_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGU2FNB_5_LC_10_9_6  (
            .in0(N__11279),
            .in1(_gnd_net_),
            .in2(N__9572),
            .in3(N__9569),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_x2_0_0_a3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_10_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_10_9_7 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_14_LC_10_9_7  (
            .in0(N__9563),
            .in1(N__9704),
            .in2(N__9554),
            .in3(N__10610),
            .lcout(\this_vga_signals.N_5_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_10_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_10_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_10_10_0  (
            .in0(N__12069),
            .in1(N__15442),
            .in2(_gnd_net_),
            .in3(N__12166),
            .lcout(\this_vga_signals.N_9_i_0_0 ),
            .ltout(\this_vga_signals.N_9_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_x1_LC_10_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_x1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_x1_LC_10_10_1 .LUT_INIT=16'b1000001111100011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_x1_LC_10_10_1  (
            .in0(N__14541),
            .in1(N__14333),
            .in2(N__9551),
            .in3(N__12367),
            .lcout(\this_vga_signals.g0_2_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI6CQQNK_2_LC_10_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI6CQQNK_2_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI6CQQNK_2_LC_10_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI6CQQNK_2_LC_10_10_2  (
            .in0(N__9608),
            .in1(N__9590),
            .in2(_gnd_net_),
            .in3(N__11284),
            .lcout(\this_vga_signals.N_57_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_x0_LC_10_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_x0_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_x0_LC_10_10_3 .LUT_INIT=16'b1101100110010001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_x0_LC_10_10_3  (
            .in0(N__14374),
            .in1(N__9548),
            .in2(N__14576),
            .in3(N__12368),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_ns_LC_10_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_ns_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_ns_LC_10_10_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_ns_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__11283),
            .in2(N__9542),
            .in3(N__9539),
            .lcout(\this_vga_signals.N_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_10_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_10_10_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_0_a2_LC_10_10_5  (
            .in0(N__12167),
            .in1(_gnd_net_),
            .in2(N__15452),
            .in3(N__12070),
            .lcout(\this_vga_signals.N_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5RUBJ1_5_LC_10_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5RUBJ1_5_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5RUBJ1_5_LC_10_10_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5RUBJ1_5_LC_10_10_6  (
            .in0(N__15136),
            .in1(N__12560),
            .in2(N__14579),
            .in3(N__12165),
            .lcout(\this_vga_signals.m6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_10_7 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_LC_10_10_7  (
            .in0(N__12164),
            .in1(N__11339),
            .in2(N__9641),
            .in3(N__12068),
            .lcout(\this_vga_signals.mult1_un61_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_10_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_11_LC_10_11_0 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_11_LC_10_11_0  (
            .in0(N__9674),
            .in1(N__12280),
            .in2(N__9692),
            .in3(N__12268),
            .lcout(\this_vga_signals.if_i3_mux_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI820378_2_LC_10_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI820378_2_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI820378_2_LC_10_11_1 .LUT_INIT=16'b0110110000110110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI820378_2_LC_10_11_1  (
            .in0(N__14369),
            .in1(N__11381),
            .in2(N__14577),
            .in3(N__12373),
            .lcout(\this_vga_signals.M_vcounter_q_RNI820378Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_10_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_10_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_8_LC_10_11_2  (
            .in0(N__15362),
            .in1(N__12084),
            .in2(_gnd_net_),
            .in3(N__12191),
            .lcout(),
            .ltout(\this_vga_signals.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_LC_10_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_LC_10_11_3 .LUT_INIT=16'b1101101001111010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_LC_10_11_3  (
            .in0(N__14372),
            .in1(N__11287),
            .in2(N__9602),
            .in3(N__12375),
            .lcout(),
            .ltout(\this_vga_signals.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_10_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_10_11_4 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__14551),
            .in2(N__9599),
            .in3(N__9710),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI820378_0_2_LC_10_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI820378_0_2_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI820378_0_2_LC_10_11_5 .LUT_INIT=16'b0011011001101100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI820378_0_2_LC_10_11_5  (
            .in0(N__14370),
            .in1(N__11380),
            .in2(N__14578),
            .in3(N__12372),
            .lcout(\this_vga_signals.M_vcounter_q_RNI820378_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_2_LC_10_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_2_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_0_a3_2_LC_10_11_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_0_a3_2_LC_10_11_6  (
            .in0(N__14378),
            .in1(N__12083),
            .in2(N__15425),
            .in3(N__12190),
            .lcout(),
            .ltout(\this_vga_signals.g0_3_0_a3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_10_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_LC_10_11_7 .LUT_INIT=16'b1110011110111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_LC_10_11_7  (
            .in0(N__14371),
            .in1(N__11286),
            .in2(N__9713),
            .in3(N__12374),
            .lcout(\this_vga_signals.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_1_LC_10_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_1_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_1_LC_10_12_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_a4_1_1_LC_10_12_0  (
            .in0(N__12548),
            .in1(N__14303),
            .in2(N__15125),
            .in3(N__15414),
            .lcout(\this_vga_signals.if_m10_0_a4_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_10_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_10_12_1 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_1_LC_10_12_1  (
            .in0(N__14305),
            .in1(N__12082),
            .in2(N__15448),
            .in3(N__12189),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_10_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_10_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_10_12_2  (
            .in0(N__11620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12724),
            .lcout(\this_vga_signals.N_188_0 ),
            .ltout(\this_vga_signals.N_188_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC471_9_LC_10_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC471_9_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEC471_9_LC_10_12_3 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIEC471_9_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__15191),
            .in2(N__9695),
            .in3(N__16613),
            .lcout(\this_vga_signals.CO0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_0_0_0_LC_10_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_0_0_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_0_0_0_LC_10_12_4 .LUT_INIT=16'b0000000010000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_a4_0_0_0_LC_10_12_4  (
            .in0(N__12550),
            .in1(N__14304),
            .in2(N__15126),
            .in3(N__15415),
            .lcout(\this_vga_signals.if_m10_0_a4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_3_0_LC_10_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_3_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_3_0_LC_10_12_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_3_0_LC_10_12_5  (
            .in0(N__11324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12632),
            .lcout(),
            .ltout(\this_vga_signals.g1_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_10_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_10_12_6 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_LC_10_12_6  (
            .in0(N__12549),
            .in1(N__11398),
            .in2(N__9683),
            .in3(N__9680),
            .lcout(\this_vga_signals.if_N_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_10_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_10_12_7 .LUT_INIT=16'b1000000110110111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_c2_LC_10_12_7  (
            .in0(N__15044),
            .in1(N__13700),
            .in2(N__15447),
            .in3(N__12808),
            .lcout(\this_vga_signals.mult1_un47_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_ns_LC_10_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_ns_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_ns_LC_10_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_ns_LC_10_13_0  (
            .in0(N__11453),
            .in1(N__9722),
            .in2(_gnd_net_),
            .in3(N__11420),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_LC_10_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_LC_10_13_1 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_LC_10_13_1  (
            .in0(N__13805),
            .in1(N__13160),
            .in2(N__9728),
            .in3(N__11725),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_13_2 .LUT_INIT=16'b1010010110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_10_13_2  (
            .in0(N__13697),
            .in1(N__13912),
            .in2(N__9725),
            .in3(N__15029),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_10_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_10_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13038),
            .lcout(this_vga_signals_M_vcounter_q_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24981),
            .ce(N__15520),
            .sr(N__15493));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_0_LC_10_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_0_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_0_LC_10_13_4 .LUT_INIT=16'b0000110011001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_0_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__9803),
            .in2(N__9821),
            .in3(N__9784),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_13_6 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_13_6  (
            .in0(N__13315),
            .in1(N__13911),
            .in2(N__13705),
            .in3(N__12806),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13107),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24981),
            .ce(N__15520),
            .sr(N__15493));
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_14_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_10_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_10_14_0  (
            .in0(N__17144),
            .in1(N__13965),
            .in2(N__16682),
            .in3(N__16678),
            .lcout(this_vga_signals_M_vcounter_q_0),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__24986),
            .ce(),
            .sr(N__15492));
    defparam \this_vga_signals.M_vcounter_q_1_LC_10_14_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_10_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_10_14_1  (
            .in0(N__17146),
            .in1(N__14066),
            .in2(_gnd_net_),
            .in3(N__9716),
            .lcout(this_vga_signals_M_vcounter_q_1),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__24986),
            .ce(),
            .sr(N__15492));
    defparam \this_vga_signals.M_vcounter_q_2_LC_10_14_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_10_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_10_14_2  (
            .in0(N__17145),
            .in1(N__14470),
            .in2(_gnd_net_),
            .in3(N__9752),
            .lcout(this_vga_signals_M_vcounter_q_2),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__24986),
            .ce(),
            .sr(N__15492));
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_14_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_10_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_10_14_3  (
            .in0(N__17147),
            .in1(N__14254),
            .in2(_gnd_net_),
            .in3(N__9749),
            .lcout(this_vga_signals_M_vcounter_q_3),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__24986),
            .ce(),
            .sr(N__15492));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_14_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__15358),
            .in2(_gnd_net_),
            .in3(N__9746),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_14_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__15083),
            .in2(_gnd_net_),
            .in3(N__9743),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_14_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__13690),
            .in2(_gnd_net_),
            .in3(N__9740),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_14_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__13584),
            .in2(_gnd_net_),
            .in3(N__9737),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_15_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__13797),
            .in2(_gnd_net_),
            .in3(N__9734),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_10_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_10_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__16630),
            .in2(_gnd_net_),
            .in3(N__9731),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_10_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13173),
            .lcout(this_vga_signals_M_vcounter_q_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24994),
            .ce(N__15518),
            .sr(N__15490));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_9_LC_10_15_3  (
            .in0(N__13174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24994),
            .ce(N__15518),
            .sr(N__15490));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_15_4  (
            .in0(N__13081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24994),
            .ce(N__15518),
            .sr(N__15490));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13080),
            .lcout(this_vga_signals_M_vcounter_q_8_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24994),
            .ce(N__15518),
            .sr(N__15490));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_c2_LC_10_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_c2_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_c2_LC_10_16_0 .LUT_INIT=16'b0010001010111011;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_c2_LC_10_16_0  (
            .in0(N__13022),
            .in1(N__11767),
            .in2(_gnd_net_),
            .in3(N__12725),
            .lcout(\this_vga_signals.mult1_un40_sum_1_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_10_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_10_16_1 .LUT_INIT=16'b0011011100010011;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_ac0_3_0_LC_10_16_1  (
            .in0(N__13321),
            .in1(N__11674),
            .in2(N__11561),
            .in3(N__13021),
            .lcout(\this_vga_signals.mult1_un40_sum_0_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_0_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_3_LC_10_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_3_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_3_LC_10_16_2 .LUT_INIT=16'b0110001011000000;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_3_LC_10_16_2  (
            .in0(N__11569),
            .in1(N__9894),
            .in2(N__9824),
            .in3(N__11755),
            .lcout(\this_vga_signals.mult1_un40_sum_m_x0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_7_LC_10_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_7_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_7_LC_10_16_3 .LUT_INIT=16'b0100110110011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_7_LC_10_16_3  (
            .in0(N__9817),
            .in1(N__9802),
            .in2(N__11447),
            .in3(N__9788),
            .lcout(\this_vga_signals.N_81_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_3_LC_10_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_3_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_3_LC_10_16_4 .LUT_INIT=16'b1001011000010100;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_3_LC_10_16_4  (
            .in0(N__9895),
            .in1(N__11756),
            .in2(N__11573),
            .in3(N__9773),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_m_x1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_3_LC_10_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_3_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_3_LC_10_16_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_3_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__9767),
            .in2(N__9761),
            .in3(N__9758),
            .lcout(\this_vga_signals.mult1_un40_sum_m_ns_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m12_0_o2_381_10_1_LC_10_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_m12_0_o2_381_10_1_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m12_0_o2_381_10_1_LC_10_16_6 .LUT_INIT=16'b0011111101010101;
    LogicCell40 \this_ppu.M_m12_0_o2_381_10_1_LC_10_16_6  (
            .in0(N__15201),
            .in1(N__14301),
            .in2(N__13370),
            .in3(N__15127),
            .lcout(\this_ppu.M_m12_0_o2_381_10Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axbxc2_LC_10_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axbxc2_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axbxc2_LC_10_17_0 .LUT_INIT=16'b1011101111011101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axbxc2_LC_10_17_0  (
            .in0(N__13698),
            .in1(N__11557),
            .in2(_gnd_net_),
            .in3(N__13317),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_2_LC_10_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_2_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_2_LC_10_17_1 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_2_LC_10_17_1  (
            .in0(N__11738),
            .in1(N__9899),
            .in2(N__9878),
            .in3(N__11675),
            .lcout(\this_vga_signals.mult1_un40_sum_m_ns_2 ),
            .ltout(\this_vga_signals.mult1_un40_sum_m_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1_LC_10_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1_LC_10_17_2 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1_LC_10_17_2  (
            .in0(N__13929),
            .in1(_gnd_net_),
            .in2(N__9875),
            .in3(N__15093),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_10_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_10_17_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_6_LC_10_17_3  (
            .in0(N__12943),
            .in1(N__13369),
            .in2(_gnd_net_),
            .in3(N__13699),
            .lcout(\this_vga_signals.N_196_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_17_4 .LUT_INIT=16'b0111001100110001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_10_17_4  (
            .in0(N__13928),
            .in1(N__13211),
            .in2(N__13322),
            .in3(N__11879),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0),
            .ltout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un47_sum_c3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_LC_10_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_LC_10_17_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9851),
            .in3(N__13930),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1),
            .ltout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un54_sum_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m7_1_LC_10_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_m7_1_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m7_1_LC_10_17_6 .LUT_INIT=16'b1100111110000001;
    LogicCell40 \this_ppu.M_m7_1_LC_10_17_6  (
            .in0(N__13977),
            .in1(N__11835),
            .in2(N__9839),
            .in3(N__10600),
            .lcout(\this_ppu.M_m7Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_10_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_10_18_0 .LUT_INIT=16'b1011111100000000;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_LC_10_18_0  (
            .in0(N__11630),
            .in1(N__10491),
            .in2(N__14561),
            .in3(N__11975),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_c3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_m3_LC_10_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_m3_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_m3_LC_10_18_1 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_m3_LC_10_18_1  (
            .in0(N__14345),
            .in1(N__13931),
            .in2(_gnd_net_),
            .in3(N__11954),
            .lcout(this_vga_signals_un4_lcounter_if_i1_mux),
            .ltout(this_vga_signals_un4_lcounter_if_i1_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_10_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_10_18_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_10_18_2  (
            .in0(N__11955),
            .in1(_gnd_net_),
            .in2(N__10604),
            .in3(N__10519),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0),
            .ltout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_18_3 .LUT_INIT=16'b1000011111100001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_LC_10_18_3  (
            .in0(N__11933),
            .in1(N__11831),
            .in2(N__10580),
            .in3(N__11786),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un68_sum_axbxc3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m7_LC_10_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_m7_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m7_LC_10_18_4 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \this_ppu.M_m7_LC_10_18_4  (
            .in0(N__14512),
            .in1(N__14091),
            .in2(_gnd_net_),
            .in3(N__10565),
            .lcout(),
            .ltout(\this_ppu.M_N_11_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIFN38L2_LC_10_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIFN38L2_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIFN38L2_LC_10_18_5 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \this_ppu.M_state_q_RNIFN38L2_LC_10_18_5  (
            .in0(N__10559),
            .in1(N__14699),
            .in2(N__10550),
            .in3(N__15094),
            .lcout(\this_ppu.M_m12_0_o2_381_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam d_m1_0_LC_10_18_6.C_ON=1'b0;
    defparam d_m1_0_LC_10_18_6.SEQ_MODE=4'b0000;
    defparam d_m1_0_LC_10_18_6.LUT_INIT=16'b1001011001101001;
    LogicCell40 d_m1_0_LC_10_18_6 (
            .in0(N__11956),
            .in1(N__10534),
            .in2(N__10523),
            .in3(N__11844),
            .lcout(this_vga_signals_un4_lcounter_if_generate_plus_mult1_un61_sum_axbxc3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_m14_0_x3_LC_10_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_m14_0_x3_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_m14_0_x3_LC_10_18_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_m14_0_x3_LC_10_18_7  (
            .in0(N__14346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11830),
            .lcout(this_vga_signals_un4_lcounter_if_N_7_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_LC_10_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_LC_10_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_state_q_RNO_0_LC_10_19_0  (
            .in0(N__10365),
            .in1(N__10224),
            .in2(N__10083),
            .in3(N__9935),
            .lcout(),
            .ltout(\this_ppu.un1_M_state_d8_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_LC_10_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_LC_10_19_1 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \this_ppu.M_state_q_LC_10_19_1  (
            .in0(N__22365),
            .in1(N__10691),
            .in2(N__9908),
            .in3(N__9905),
            .lcout(M_this_ppu_vram_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25012),
            .ce(),
            .sr(N__24743));
    defparam \this_ppu.M_state_q_RNO_1_LC_10_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_1_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_1_LC_10_19_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_state_q_RNO_1_LC_10_19_2  (
            .in0(N__10994),
            .in1(N__10859),
            .in2(N__10728),
            .in3(N__22363),
            .lcout(\this_ppu.un1_M_state_d8_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_10_19_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_10_19_5 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_0_11_LC_10_19_5  (
            .in0(N__22811),
            .in1(N__22085),
            .in2(N__22301),
            .in3(N__21818),
            .lcout(),
            .ltout(M_this_sprites_ram_read_data_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_vram_write_data_0_i_0_LC_10_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_0_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_0_LC_10_19_6 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \this_vga_signals.M_this_vram_write_data_0_i_0_LC_10_19_6  (
            .in0(N__20882),
            .in1(N__23501),
            .in2(N__10685),
            .in3(N__22364),
            .lcout(M_this_vram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_10_20_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_10_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_10_20_3  (
            .in0(N__10670),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25016),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_10_20_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_10_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10619),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25016),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_10_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_10_20_6 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIOLTE3_6_LC_10_20_6  (
            .in0(N__10658),
            .in1(N__14513),
            .in2(N__11663),
            .in3(N__13706),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_10_20_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_10_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10625),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25016),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_x0_LC_11_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_x0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_x0_LC_11_9_0 .LUT_INIT=16'b0100011001101110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_x0_LC_11_9_0  (
            .in0(N__11996),
            .in1(N__14384),
            .in2(N__12376),
            .in3(N__14574),
            .lcout(),
            .ltout(\this_vga_signals.g0_16_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_ns_LC_11_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_ns_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_ns_LC_11_9_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_ns_LC_11_9_1  (
            .in0(N__11273),
            .in1(_gnd_net_),
            .in2(N__10613),
            .in3(N__12305),
            .lcout(\this_vga_signals.g3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_a2_0_LC_11_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_a2_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_a2_0_LC_11_9_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_a2_0_LC_11_9_2  (
            .in0(N__12091),
            .in1(N__11271),
            .in2(N__14387),
            .in3(N__11213),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_11_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_11_9_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_1_LC_11_9_3  (
            .in0(N__11274),
            .in1(N__14126),
            .in2(_gnd_net_),
            .in3(N__12362),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_11_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_11_9_4 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_11_9_4  (
            .in0(N__14383),
            .in1(N__11174),
            .in2(N__11168),
            .in3(N__11165),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI5DK9PN1_7_LC_11_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI5DK9PN1_7_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI5DK9PN1_7_LC_11_9_5 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI5DK9PN1_7_LC_11_9_5  (
            .in0(N__23854),
            .in1(N__12206),
            .in2(N__11159),
            .in3(N__11138),
            .lcout(this_vga_signals_address_0_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_11_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_11_9_6 .LUT_INIT=16'b1011011100100001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_11_9_6  (
            .in0(N__11144),
            .in1(N__14127),
            .in2(N__11132),
            .in3(N__14575),
            .lcout(\this_vga_signals.mult1_un75_sum_c2_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_0_LC_11_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_0_LC_11_9_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_0_LC_11_9_7  (
            .in0(N__11272),
            .in1(N__11219),
            .in2(N__11123),
            .in3(N__12361),
            .lcout(\this_vga_signals.g3_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_1_0_LC_11_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_1_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_1_0_LC_11_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_1_0_LC_11_10_0  (
            .in0(N__12171),
            .in1(N__12065),
            .in2(N__15153),
            .in3(N__12561),
            .lcout(\this_vga_signals.g3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_LC_11_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_LC_11_10_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_N_4_i_0_LC_11_10_1  (
            .in0(N__12456),
            .in1(N__11193),
            .in2(N__12088),
            .in3(N__12169),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_i ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_11_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_2_LC_11_10_2 .LUT_INIT=16'b1000111011101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_2_LC_11_10_2  (
            .in0(N__14540),
            .in1(N__14365),
            .in2(N__11114),
            .in3(N__11275),
            .lcout(\this_vga_signals.g1_2 ),
            .ltout(\this_vga_signals.g1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_11_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_m2_LC_11_10_3 .LUT_INIT=16'b1011011100010010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_m2_LC_11_10_3  (
            .in0(N__14366),
            .in1(N__15446),
            .in2(N__11291),
            .in3(N__12298),
            .lcout(\this_vga_signals.N_57_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_10_4 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_LC_11_10_4  (
            .in0(N__12172),
            .in1(N__15429),
            .in2(N__14386),
            .in3(N__12067),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOH6PPC_5_LC_11_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOH6PPC_5_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOH6PPC_5_LC_11_10_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIOH6PPC_5_LC_11_10_5  (
            .in0(N__11276),
            .in1(N__12575),
            .in2(N__11222),
            .in3(N__12366),
            .lcout(\this_vga_signals.m48_i_x4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_11_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_11_10_6 .LUT_INIT=16'b1110100011010100;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_LC_11_10_6  (
            .in0(N__12170),
            .in1(N__15430),
            .in2(N__14385),
            .in3(N__12066),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_x_LC_11_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_x_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_x_LC_11_10_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_N_4_i_0_x_LC_11_10_7  (
            .in0(N__12457),
            .in1(N__11194),
            .in2(_gnd_net_),
            .in3(N__12168),
            .lcout(\this_vga_signals.N_4_i_0_x ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_1_LC_11_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_N_4_i_0_1_LC_11_11_0 .LUT_INIT=16'b0001110011011110;
    LogicCell40 \this_vga_signals.un5_vaddress_N_4_i_0_1_LC_11_11_0  (
            .in0(N__12533),
            .in1(N__15105),
            .in2(N__15450),
            .in3(N__12383),
            .lcout(\this_vga_signals.N_4_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_1_LC_11_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_1_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_1_LC_11_11_1 .LUT_INIT=16'b0100000100011010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_1_LC_11_11_1  (
            .in0(N__15104),
            .in1(N__12532),
            .in2(N__15424),
            .in3(N__12639),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_11_2 .LUT_INIT=16'b1111110001000101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_11_2  (
            .in0(N__11330),
            .in1(N__12660),
            .in2(N__11180),
            .in3(N__11465),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.g0_0_i_o3_LC_11_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.g0_0_i_o3_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.g0_0_i_o3_LC_11_11_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.g0_0_i_o3_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11177),
            .in3(N__12175),
            .lcout(\this_vga_signals.N_81_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_x2_0_0_LC_11_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_x2_0_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_x2_0_0_LC_11_11_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_x2_0_0_LC_11_11_4  (
            .in0(N__12534),
            .in1(N__14306),
            .in2(N__15451),
            .in3(N__15106),
            .lcout(),
            .ltout(\this_vga_signals.if_m10_0_x2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_LC_11_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_LC_11_11_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_a4_LC_11_11_5  (
            .in0(N__11405),
            .in1(N__12071),
            .in2(N__11357),
            .in3(N__12174),
            .lcout(\this_vga_signals.if_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_11_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_11_11_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_11_11_6  (
            .in0(N__12817),
            .in1(N__11495),
            .in2(N__11354),
            .in3(N__11464),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_x2_LC_11_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_x2_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_x2_LC_11_11_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_x2_LC_11_11_7  (
            .in0(N__12661),
            .in1(N__11399),
            .in2(N__11345),
            .in3(N__12072),
            .lcout(\this_vga_signals.if_N_7_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_11_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_11_12_0 .LUT_INIT=16'b0000011100000001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_0_LC_11_12_0  (
            .in0(N__11494),
            .in1(N__11540),
            .in2(N__11524),
            .in3(N__12807),
            .lcout(\this_vga_signals.mult1_un47_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_12_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__11314),
            .in2(N__11342),
            .in3(N__12628),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_11_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m2_1_LC_11_12_2 .LUT_INIT=16'b1000000100100100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m2_1_LC_11_12_2  (
            .in0(N__14302),
            .in1(N__15064),
            .in2(N__15427),
            .in3(N__12538),
            .lcout(\this_vga_signals.if_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x1_LC_11_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x1_LC_11_12_3 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x1_LC_11_12_3  (
            .in0(N__12536),
            .in1(N__15369),
            .in2(N__11329),
            .in3(N__12630),
            .lcout(\this_vga_signals.if_m10_0_a4_1_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x0_LC_11_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x0_LC_11_12_4 .LUT_INIT=16'b0100100010000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_x0_LC_11_12_4  (
            .in0(N__12631),
            .in1(N__15432),
            .in2(N__11325),
            .in3(N__12537),
            .lcout(),
            .ltout(\this_vga_signals.if_m10_0_a4_1_0_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_ns_LC_11_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_ns_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_ns_LC_11_12_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m10_0_a4_1_0_ns_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__11414),
            .in2(N__11408),
            .in3(N__11397),
            .lcout(\this_vga_signals.if_m10_0_a4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_11_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_11_12_6 .LUT_INIT=16'b0111000110111100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_11_12_6  (
            .in0(N__12629),
            .in1(N__15063),
            .in2(N__15426),
            .in3(N__12535),
            .lcout(\this_vga_signals.mult1_un54_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIK5K7M3_4_LC_11_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIK5K7M3_4_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIK5K7M3_4_LC_11_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIK5K7M3_4_LC_11_12_7  (
            .in0(N__15433),
            .in1(N__12073),
            .in2(_gnd_net_),
            .in3(N__12173),
            .lcout(\this_vga_signals.g0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x1_LC_11_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x1_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x1_LC_11_13_0 .LUT_INIT=16'b0110100111100001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x1_LC_11_13_0  (
            .in0(N__13066),
            .in1(N__12851),
            .in2(N__12816),
            .in3(N__12967),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_11_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_11_13_1 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_LC_11_13_1  (
            .in0(N__11616),
            .in1(N__13187),
            .in2(N__12723),
            .in3(N__13651),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNISGOS_4_LC_11_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNISGOS_4_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNISGOS_4_LC_11_13_2 .LUT_INIT=16'b1111111000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNISGOS_4_LC_11_13_2  (
            .in0(N__13583),
            .in1(N__12999),
            .in2(N__11621),
            .in3(N__13799),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_fast_esr_RNISGOSZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIP2HP1_5_LC_11_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIP2HP1_5_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIP2HP1_5_LC_11_13_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIP2HP1_5_LC_11_13_3  (
            .in0(N__12713),
            .in1(_gnd_net_),
            .in2(N__11372),
            .in3(N__12731),
            .lcout(\this_vga_signals.vaddress_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x0_LC_11_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x0_LC_11_13_4 .LUT_INIT=16'b0001111001111000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_x0_LC_11_13_4  (
            .in0(N__13067),
            .in1(N__12852),
            .in2(N__12815),
            .in3(N__12968),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_ns_LC_11_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_ns_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_ns_LC_11_13_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_1_ns_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__12404),
            .in2(N__11369),
            .in3(N__11366),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_11_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_11_13_6 .LUT_INIT=16'b0010110100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_11_13_6  (
            .in0(N__12804),
            .in1(N__11520),
            .in2(N__11360),
            .in3(N__11538),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_11_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_11_13_7 .LUT_INIT=16'b0000010011111011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_11_13_7  (
            .in0(N__11539),
            .in1(N__12805),
            .in2(N__11525),
            .in3(N__12624),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_a2_1_LC_11_14_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_a2_1_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_a2_1_LC_11_14_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_state_d_0_sqmuxa_i_0_0_a2_1_LC_11_14_0  (
            .in0(N__11439),
            .in1(N__11715),
            .in2(_gnd_net_),
            .in3(N__11695),
            .lcout(N_475),
            .ltout(N_475_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m1_e_LC_11_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_e_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_e_LC_11_14_1 .LUT_INIT=16'b1000101000001010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_e_LC_11_14_1  (
            .in0(N__13146),
            .in1(N__12706),
            .in2(N__11501),
            .in3(N__11609),
            .lcout(\this_vga_signals.if_N_3_mux ),
            .ltout(\this_vga_signals.if_N_3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axbxc1_LC_11_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axbxc1_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axbxc1_LC_11_14_2 .LUT_INIT=16'b0110110010010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axbxc1_LC_11_14_2  (
            .in0(N__13065),
            .in1(N__12961),
            .in2(N__11498),
            .in3(N__12405),
            .lcout(\this_vga_signals.mult1_un47_sum_axb2_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axb2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_11_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_11_14_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__11480),
            .in2(N__11474),
            .in3(N__11471),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13111),
            .lcout(this_vga_signals_M_vcounter_q_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24982),
            .ce(N__15521),
            .sr(N__15491));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_11_14_5  (
            .in0(N__12673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_M_vcounter_q_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24982),
            .ce(N__15521),
            .sr(N__15491));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x1_LC_11_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x1_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x1_LC_11_14_6 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x1_LC_11_14_6  (
            .in0(N__12705),
            .in1(N__11596),
            .in2(N__11443),
            .in3(N__11694),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0_1_0_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x0_LC_11_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x0_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x0_LC_11_14_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c3_0_1_0_x0_LC_11_14_7  (
            .in0(N__11595),
            .in1(N__12704),
            .in2(_gnd_net_),
            .in3(N__11435),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0_1_0_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axb2_LC_11_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axb2_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axb2_LC_11_15_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_axb2_LC_11_15_2  (
            .in0(N__14623),
            .in1(N__11848),
            .in2(_gnd_net_),
            .in3(N__11960),
            .lcout(\this_vga_signals.mult1_un61_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15537),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24987),
            .ce(N__15519),
            .sr(N__15488));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15538),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24987),
            .ce(N__15519),
            .sr(N__15488));
    defparam \this_vga_signals.un4_lcounter_if_m5_0_1_LC_11_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_m5_0_1_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_m5_0_1_LC_11_16_0 .LUT_INIT=16'b0110110111111001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_m5_0_1_LC_11_16_0  (
            .in0(N__11699),
            .in1(N__13145),
            .in2(N__11732),
            .in3(N__13019),
            .lcout(\this_vga_signals.if_m5_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_1_LC_11_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_1_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_1_LC_11_16_1 .LUT_INIT=16'b0000110011100001;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_1_LC_11_16_1  (
            .in0(N__13018),
            .in1(N__11727),
            .in2(N__13154),
            .in3(N__11697),
            .lcout(\this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axb1_LC_11_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axb1_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axb1_LC_11_16_2 .LUT_INIT=16'b0001100010010110;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axb1_LC_11_16_2  (
            .in0(N__13791),
            .in1(N__13674),
            .in2(N__16615),
            .in3(N__13556),
            .lcout(\this_vga_signals.mult1_un40_sum_1_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_LC_11_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_LC_11_16_3 .LUT_INIT=16'b1001010101101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_LC_11_16_3  (
            .in0(N__13017),
            .in1(N__11728),
            .in2(N__13155),
            .in3(N__11698),
            .lcout(\this_vga_signals.N_370_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axb1_LC_11_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axb1_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axb1_LC_11_16_4 .LUT_INIT=16'b0101100010110110;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_0_axb1_LC_11_16_4  (
            .in0(N__13790),
            .in1(N__13555),
            .in2(N__16614),
            .in3(N__13020),
            .lcout(\this_vga_signals.mult1_un40_sum_0_axb1_i ),
            .ltout(\this_vga_signals.mult1_un40_sum_0_axb1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_1_LC_11_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_1_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_1_LC_11_16_5 .LUT_INIT=16'b0101010110010101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x1_1_LC_11_16_5  (
            .in0(N__13293),
            .in1(N__16588),
            .in2(N__11543),
            .in3(N__13792),
            .lcout(\this_vga_signals.mult1_un40_sum_m_x1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axbxc2_LC_11_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axbxc2_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axbxc2_LC_11_16_6 .LUT_INIT=16'b1100011010011100;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_1_axbxc2_LC_11_16_6  (
            .in0(N__11768),
            .in1(N__11754),
            .in2(N__13314),
            .in3(N__13675),
            .lcout(\this_vga_signals.mult1_un40_sum1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_0_LC_11_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_0_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_0_LC_11_16_7 .LUT_INIT=16'b0110010110011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIELM41_0_LC_11_16_7  (
            .in0(N__13016),
            .in1(N__11726),
            .in2(N__13153),
            .in3(N__11696),
            .lcout(\this_vga_signals.N_330_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8MCG1_9_LC_11_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8MCG1_9_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI8MCG1_9_LC_11_17_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI8MCG1_9_LC_11_17_0  (
            .in0(N__13354),
            .in1(N__16612),
            .in2(_gnd_net_),
            .in3(N__14128),
            .lcout(\this_vga_signals.vsync_1_0_a2_6_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_m11_1_LC_11_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_m11_1_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_m11_1_LC_11_17_1 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \this_vga_signals.un4_lcounter_if_m11_1_LC_11_17_1  (
            .in0(N__14270),
            .in1(N__13925),
            .in2(_gnd_net_),
            .in3(N__13207),
            .lcout(),
            .ltout(\this_vga_signals.if_m11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_m11_LC_11_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_m11_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_m11_LC_11_17_2 .LUT_INIT=16'b1011100011100010;
    LogicCell40 \this_vga_signals.un4_lcounter_if_m11_LC_11_17_2  (
            .in0(N__13926),
            .in1(N__13310),
            .in2(N__11648),
            .in3(N__11880),
            .lcout(this_vga_signals_un4_lcounter_if_i3_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_11_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_11_17_4 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_11_17_4  (
            .in0(N__16611),
            .in1(N__13800),
            .in2(_gnd_net_),
            .in3(N__13585),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16215),
            .lcout(\this_vga_signals.mult1_un47_sum_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_LC_11_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_LC_11_18_1 .LUT_INIT=16'b0101010001000001;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_LC_11_18_1  (
            .in0(N__14344),
            .in1(N__11916),
            .in2(N__15440),
            .in3(N__11969),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_x1_LC_11_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_x1_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_x1_LC_11_18_2 .LUT_INIT=16'b0100110000001100;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_x1_LC_11_18_2  (
            .in0(N__11899),
            .in1(N__11829),
            .in2(N__11633),
            .in3(N__11887),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_1_0_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_ns_LC_11_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_ns_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_ns_LC_11_18_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_3_1_0_ns_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__17434),
            .in2(N__11978),
            .in3(N__11929),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_1_LC_11_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_1_LC_11_18_4 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_2_1_LC_11_18_4  (
            .in0(N__15137),
            .in1(N__13924),
            .in2(_gnd_net_),
            .in3(N__13206),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_2_2_1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_2_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_sx_LC_11_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_sx_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_sx_LC_11_18_5 .LUT_INIT=16'b1010101110111110;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_sx_LC_11_18_5  (
            .in0(N__14343),
            .in1(N__15397),
            .in2(N__11963),
            .in3(N__11918),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__14624),
            .in2(_gnd_net_),
            .in3(N__11953),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_4_tz_LC_11_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_4_tz_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_4_tz_LC_11_18_7 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_4_tz_LC_11_18_7  (
            .in0(N__12942),
            .in1(N__11917),
            .in2(_gnd_net_),
            .in3(N__13847),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_2_4_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_LC_11_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_LC_11_19_2 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_LC_11_19_2  (
            .in0(N__11906),
            .in1(N__11900),
            .in2(_gnd_net_),
            .in3(N__11888),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_c2_LC_11_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_c2_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_c2_LC_11_19_3 .LUT_INIT=16'b0000011100001101;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_c2_LC_11_19_3  (
            .in0(N__14531),
            .in1(N__14347),
            .in2(N__11861),
            .in3(N__11853),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_11_20_4 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_11_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11774),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25013),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_11_20_7 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_11_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11780),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25013),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_x1_LC_12_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_x1_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_x1_LC_12_9_7 .LUT_INIT=16'b0111110000011100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_x1_LC_12_9_7  (
            .in0(N__14573),
            .in1(N__14379),
            .in2(N__11995),
            .in3(N__12357),
            .lcout(\this_vga_signals.g0_16_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIU9QNGC_4_LC_12_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIU9QNGC_4_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIU9QNGC_4_LC_12_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIU9QNGC_4_LC_12_10_1  (
            .in0(N__15431),
            .in1(N__12299),
            .in2(_gnd_net_),
            .in3(N__12287),
            .lcout(\this_vga_signals.N_57_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_12_10_2 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_12_10_2  (
            .in0(N__12587),
            .in1(N__12281),
            .in2(N__12476),
            .in3(N__12269),
            .lcout(\this_vga_signals.if_i3_mux_0_1 ),
            .ltout(\this_vga_signals.if_i3_mux_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_12_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_12_10_3 .LUT_INIT=16'b1110111000011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_12_10_3  (
            .in0(N__12235),
            .in1(N__14131),
            .in2(N__12257),
            .in3(N__14562),
            .lcout(\this_vga_signals.if_N_6_mux_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_2_LC_12_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_2_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_2_LC_12_10_4 .LUT_INIT=16'b0011011010011100;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_2_LC_12_10_4  (
            .in0(N__14563),
            .in1(N__12254),
            .in2(N__12248),
            .in3(N__12236),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_12_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_12_10_5 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_18_LC_12_10_5  (
            .in0(N__12227),
            .in1(N__12221),
            .in2(N__12215),
            .in3(N__12212),
            .lcout(\this_vga_signals.g2_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_i_LC_12_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_i_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_i_LC_12_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_i_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__15428),
            .in2(N__12192),
            .in3(N__12061),
            .lcout(\this_vga_signals.N_5_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_1_LC_12_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_1_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_1_LC_12_11_2 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_1_LC_12_11_2  (
            .in0(N__14367),
            .in1(N__15141),
            .in2(N__15441),
            .in3(N__12551),
            .lcout(),
            .ltout(\this_vga_signals.g0_10_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_12_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_12_11_3 .LUT_INIT=16'b1001000011000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_LC_12_11_3  (
            .in0(N__15143),
            .in1(N__12662),
            .in2(N__12647),
            .in3(N__12640),
            .lcout(\this_vga_signals.if_N_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_0_5_LC_12_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_0_5_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_0_5_LC_12_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI9OGF9_0_5_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__15142),
            .in2(_gnd_net_),
            .in3(N__12552),
            .lcout(\this_vga_signals.m48_i_x4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g4_1_0_LC_12_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g4_1_0_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g4_1_0_LC_12_11_5 .LUT_INIT=16'b1101111011111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g4_1_0_LC_12_11_5  (
            .in0(N__12553),
            .in1(N__15402),
            .in2(N__15154),
            .in3(N__14368),
            .lcout(\this_vga_signals.g4_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_12_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_12_11_6 .LUT_INIT=16'b0101101000111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_LC_12_11_6  (
            .in0(N__12833),
            .in1(N__12902),
            .in2(N__12743),
            .in3(N__12410),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_0_c_LC_12_12_0 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_0_c_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_0_c_LC_12_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_0_c_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__17903),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\this_vga_signals.mult1_un68_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_1_s_LC_12_12_1 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_1_s_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_1_s_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_cry_1_s_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__14630),
            .in2(N__12890),
            .in3(N__12443),
            .lcout(\this_vga_signals.mult1_un68_sum_cry_1_s ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un68_sum_cry_0 ),
            .carryout(\this_vga_signals.mult1_un68_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_axb_3_LC_12_12_2 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_axb_3_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_axb_3_LC_12_12_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_axb_3_LC_12_12_2  (
            .in0(N__15639),
            .in1(N__12440),
            .in2(N__12866),
            .in3(N__12428),
            .lcout(\this_vga_signals.mult1_un75_sum_axb_3 ),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un68_sum_cry_1 ),
            .carryout(\this_vga_signals.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_s_3_LC_12_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_s_3_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_s_3_LC_12_12_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un68_sum_s_3_LC_12_12_3  (
            .in0(N__12425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12413),
            .lcout(\this_vga_signals.mult1_un68_sum_s_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_12_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_12_12_4 .LUT_INIT=16'b0010110101111000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_12_12_4  (
            .in0(N__12406),
            .in1(N__12829),
            .in2(N__13382),
            .in3(N__12901),
            .lcout(\this_vga_signals.N_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_12_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_12_12_6 .LUT_INIT=16'b0001001001111110;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_4_LC_12_12_6  (
            .in0(N__13683),
            .in1(N__13578),
            .in2(N__13423),
            .in3(N__12857),
            .lcout(\this_vga_signals.g1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_3_LC_12_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_3_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_3_LC_12_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_3_LC_12_12_7  (
            .in0(N__12886),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un61_sum_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g6_0_LC_12_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g6_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g6_0_LC_12_13_0 .LUT_INIT=16'b0111111011001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g6_0_LC_12_13_0  (
            .in0(N__13655),
            .in1(N__13568),
            .in2(N__13424),
            .in3(N__12856),
            .lcout(\this_vga_signals.g6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI1K2D4_7_LC_12_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI1K2D4_7_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI1K2D4_7_LC_12_13_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI1K2D4_7_LC_12_13_2  (
            .in0(N__12914),
            .in1(N__14723),
            .in2(_gnd_net_),
            .in3(N__12818),
            .lcout(M_this_vga_signals_address_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_12_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_12_13_3 .LUT_INIT=16'b0011001101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_27_LC_12_13_3  (
            .in0(N__15092),
            .in1(N__13656),
            .in2(_gnd_net_),
            .in3(N__13927),
            .lcout(\this_vga_signals.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_12_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_12_13_6 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_12_13_6  (
            .in0(N__13798),
            .in1(N__12993),
            .in2(_gnd_net_),
            .in3(N__13567),
            .lcout(\this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0ASZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_12_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_12_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13045),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24977),
            .ce(N__15523),
            .sr(N__15489));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12679),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24977),
            .ce(N__15523),
            .sr(N__15489));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_12_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_12_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12680),
            .lcout(this_vga_signals_M_vcounter_q_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24977),
            .ce(N__15523),
            .sr(N__15489));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_12_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_12_15_1 .LUT_INIT=16'b0110011010111011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_c_0_1_LC_12_15_1  (
            .in0(N__13773),
            .in1(N__13545),
            .in2(_gnd_net_),
            .in3(N__13159),
            .lcout(\this_vga_signals.mult1_un47_sum_ac0_3_c_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_12_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13178),
            .lcout(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24983),
            .ce(N__15522),
            .sr(N__15487));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13112),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24983),
            .ce(N__15522),
            .sr(N__15487));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13085),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24983),
            .ce(N__15522),
            .sr(N__15487));
    defparam \this_vga_signals.un5_vaddress_if_m1_0_0_LC_12_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_0_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_0_LC_12_15_5 .LUT_INIT=16'b1100110010010011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_0_0_LC_12_15_5  (
            .in0(N__13885),
            .in1(N__13544),
            .in2(N__13297),
            .in3(N__12992),
            .lcout(\this_vga_signals.vaddress_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_12_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_12_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13049),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24983),
            .ce(N__15522),
            .sr(N__15487));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_12_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_12_15_7 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_12_15_7  (
            .in0(N__13271),
            .in1(N__13884),
            .in2(_gnd_net_),
            .in3(N__12991),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNINLU91_7_LC_12_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNINLU91_7_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNINLU91_7_LC_12_16_0 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNINLU91_7_LC_12_16_0  (
            .in0(N__12947),
            .in1(N__15984),
            .in2(N__13359),
            .in3(N__16085),
            .lcout(\this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0 ),
            .ltout(\this_vga_signals.M_this_vga_ramdac_en_i_o2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIC1F54_7_LC_12_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIC1F54_7_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIC1F54_7_LC_12_16_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIC1F54_7_LC_12_16_1  (
            .in0(N__14716),
            .in1(_gnd_net_),
            .in2(N__12905),
            .in3(N__13481),
            .lcout(N_192_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_16_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__13554),
            .in2(_gnd_net_),
            .in3(N__13788),
            .lcout(N_183_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_12_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_12_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__13292),
            .in2(_gnd_net_),
            .in3(N__13886),
            .lcout(\this_vga_signals.N_188_0_0_0 ),
            .ltout(\this_vga_signals.N_188_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_12_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_25_LC_12_16_4 .LUT_INIT=16'b1011110110111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_25_LC_12_16_4  (
            .in0(N__13394),
            .in1(N__13676),
            .in2(N__13388),
            .in3(N__13789),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_1_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_12_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_12_16_5 .LUT_INIT=16'b1101000010110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_3_LC_12_16_5  (
            .in0(N__16638),
            .in1(N__13793),
            .in2(N__13385),
            .in3(N__13557),
            .lcout(\this_vga_signals.g1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_LC_12_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_LC_12_16_6 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_LC_12_16_6  (
            .in0(N__13677),
            .in1(N__16637),
            .in2(N__13358),
            .in3(N__15878),
            .lcout(N_190_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGBLD1_7_LC_12_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGBLD1_7_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIGBLD1_7_LC_12_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIGBLD1_7_LC_12_17_2  (
            .in0(N__13802),
            .in1(N__15152),
            .in2(N__13586),
            .in3(N__15339),
            .lcout(N_275),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_1_LC_12_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_1_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_1_LC_12_17_3 .LUT_INIT=16'b1111000011010010;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_x0_1_LC_12_17_3  (
            .in0(N__16639),
            .in1(N__13801),
            .in2(N__13316),
            .in3(N__13232),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_m_x0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_1_LC_12_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_1_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_1_LC_12_17_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un40_sum_m_ns_1_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__13226),
            .in2(N__13220),
            .in3(N__13217),
            .lcout(\this_vga_signals.mult1_un40_sum_m_ns_1 ),
            .ltout(\this_vga_signals.mult1_un40_sum_m_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_a3_1_LC_12_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_a3_1_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_a3_1_LC_12_17_5 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un61_sum_ac0_2_a3_1_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__15151),
            .in2(N__13190),
            .in3(N__13923),
            .lcout(\this_vga_signals.if_N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_LC_12_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_LC_12_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un54_sum_sbtinv_LC_12_17_6  (
            .in0(N__16992),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un54_sum_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIL9AC2_7_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIL9AC2_7_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIL9AC2_7_LC_12_18_0 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIL9AC2_7_LC_12_18_0  (
            .in0(N__13433),
            .in1(N__14957),
            .in2(N__16102),
            .in3(N__14828),
            .lcout(N_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_12_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_12_18_3 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIMHLD1_7_LC_12_18_3  (
            .in0(N__16640),
            .in1(N__13803),
            .in2(N__13701),
            .in3(N__13582),
            .lcout(),
            .ltout(\this_vga_signals.N_177_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0T225_9_LC_12_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0T225_9_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0T225_9_LC_12_18_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI0T225_9_LC_12_18_4  (
            .in0(N__13439),
            .in1(N__14740),
            .in2(N__13490),
            .in3(N__13487),
            .lcout(N_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNICJJV_0_9_LC_12_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICJJV_0_9_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICJJV_0_9_LC_12_18_5 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNICJJV_0_9_LC_12_18_5  (
            .in0(N__15877),
            .in1(N__15992),
            .in2(N__15791),
            .in3(N__16093),
            .lcout(\this_vga_signals.N_269_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNILVSO_6_LC_12_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNILVSO_6_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNILVSO_6_LC_12_18_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNILVSO_6_LC_12_18_7  (
            .in0(N__15781),
            .in1(_gnd_net_),
            .in2(N__16342),
            .in3(N__16216),
            .lcout(\this_vga_signals.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_12_19_1  (
            .in0(N__17002),
            .in1(N__14918),
            .in2(_gnd_net_),
            .in3(N__14909),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1),
            .ltout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_a0_2_9_LC_12_19_2 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_a0_2_9_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_a0_2_9_LC_12_19_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_ppu.sprites_addr_1_i_a0_2_9_LC_12_19_2  (
            .in0(N__17799),
            .in1(N__17888),
            .in2(N__13427),
            .in3(N__18099),
            .lcout(\this_ppu.sprites_addr_1_i_a0_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o2_4_LC_12_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o2_4_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o2_4_LC_12_19_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_o2_4_LC_12_19_3  (
            .in0(N__14687),
            .in1(N__14670),
            .in2(_gnd_net_),
            .in3(N__14645),
            .lcout(\this_vga_signals.N_185_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_o2_LC_12_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_o2_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_o2_LC_12_20_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_o2_LC_12_20_2  (
            .in0(N__14672),
            .in1(N__14641),
            .in2(_gnd_net_),
            .in3(N__14685),
            .lcout(N_175_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_12_20_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_12_20_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_12_20_3  (
            .in0(N__14686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14671),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25006),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_LC_13_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_LC_13_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un61_sum_sbtinv_LC_13_13_4  (
            .in0(N__18100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un61_sum_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_0_LC_13_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_0_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_0_LC_13_13_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \this_vga_signals.un4_lcounter_if_generate_plus_mult1_un54_sum_axbxc1_0_LC_13_13_7  (
            .in0(N__14334),
            .in1(N__15236),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vram_addr_1_i_7_LC_13_14_0 .C_ON=1'b0;
    defparam \this_ppu.vram_addr_1_i_7_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vram_addr_1_i_7_LC_13_14_0 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \this_ppu.vram_addr_1_i_7_LC_13_14_0  (
            .in0(N__15790),
            .in1(N__15991),
            .in2(N__23843),
            .in3(N__16092),
            .lcout(N_90_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m11_0_LC_13_14_5 .C_ON=1'b0;
    defparam \this_ppu.M_m11_0_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m11_0_LC_13_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_m11_0_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__14471),
            .in2(_gnd_net_),
            .in3(N__14255),
            .lcout(N_184_0),
            .ltout(N_184_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_13_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_13_14_6 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(N__14067),
            .in2(N__13991),
            .in3(N__13966),
            .lcout(\this_vga_signals.N_272_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_0_c_LC_13_15_0 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_0_c_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_0_c_LC_13_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_0_c_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__17803),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\this_vga_signals.mult1_un75_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_1_c_inv_LC_13_15_1 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_1_c_inv_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_1_c_inv_LC_13_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_1_c_inv_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__14783),
            .in2(N__15661),
            .in3(N__17901),
            .lcout(G_504),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un75_sum_cry_0 ),
            .carryout(\this_vga_signals.mult1_un75_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_13_15_2 .C_ON=1'b1;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_13_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__14762),
            .in2(N__14777),
            .in3(N__15657),
            .lcout(G_503),
            .ltout(),
            .carryin(\this_vga_signals.mult1_un75_sum_cry_1 ),
            .carryout(\this_vga_signals.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_s_3_LC_13_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_s_3_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_s_3_LC_13_15_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un4_pcounter_if_generate_plus_mult1_un75_sum_s_3_LC_13_15_3  (
            .in0(N__14756),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14747),
            .lcout(\this_vga_signals.N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_m12_0_o2_381_4_LC_13_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_m12_0_o2_381_4_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_m12_0_o2_381_4_LC_13_16_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_m12_0_o2_381_4_LC_13_16_5  (
            .in0(N__17897),
            .in1(N__16967),
            .in2(N__17807),
            .in3(N__16197),
            .lcout(),
            .ltout(\this_ppu.M_m12_0_o2_381Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI38322_LC_13_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI38322_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI38322_LC_13_16_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_ppu.M_state_q_RNI38322_LC_13_16_6  (
            .in0(N__22384),
            .in1(N__18066),
            .in2(N__14744),
            .in3(N__15959),
            .lcout(),
            .ltout(\this_ppu.M_m12_0_o2_381_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIIL1T5_LC_13_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIIL1T5_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIIL1T5_LC_13_16_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_ppu.M_state_q_RNIIL1T5_LC_13_16_7  (
            .in0(N__14945),
            .in1(N__14741),
            .in2(N__14726),
            .in3(N__14715),
            .lcout(\this_ppu.M_m12_0_o2_381_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_0_6_LC_13_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_0_6_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_0_6_LC_13_17_3 .LUT_INIT=16'b1001010111010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_0_6_LC_13_17_3  (
            .in0(N__15938),
            .in1(N__15844),
            .in2(N__16063),
            .in3(N__14843),
            .lcout(\this_vga_signals.SUM_7_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_13_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_6_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_6_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15806),
            .lcout(\this_vga_signals.M_hcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24988),
            .ce(N__15706),
            .sr(N__17057));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_6_LC_13_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_6_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_6_LC_13_17_5 .LUT_INIT=16'b1100100101101100;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNIPK611_6_LC_13_17_5  (
            .in0(N__15845),
            .in1(N__14844),
            .in2(N__16064),
            .in3(N__15939),
            .lcout(\this_vga_signals.N_336_0 ),
            .ltout(\this_vga_signals.N_336_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_17_6 .LUT_INIT=16'b0111010000100010;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_17_6  (
            .in0(N__14845),
            .in1(N__16284),
            .in2(N__14849),
            .in3(N__14801),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI21GQ_6_LC_13_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI21GQ_6_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_fast_esr_RNI21GQ_6_LC_13_18_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \this_vga_signals.M_hcounter_q_fast_esr_RNI21GQ_6_LC_13_18_0  (
            .in0(N__16168),
            .in1(_gnd_net_),
            .in2(N__16314),
            .in3(N__14846),
            .lcout(\this_vga_signals.N_287 ),
            .ltout(\this_vga_signals.N_287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_18_1 .LUT_INIT=16'b0100111001010101;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_18_1  (
            .in0(N__14804),
            .in1(N__16170),
            .in2(N__14822),
            .in3(N__14819),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_13_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_13_18_2 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__14890),
            .in2(N__14813),
            .in3(N__14863),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3),
            .ltout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un61_sum_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_c3_LC_13_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_c3_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_c3_LC_13_18_3 .LUT_INIT=16'b0000010011011111;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_c3_LC_13_18_3  (
            .in0(N__16955),
            .in1(N__16171),
            .in2(N__14810),
            .in3(N__15685),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x0_LC_13_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x0_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x0_LC_13_18_4 .LUT_INIT=16'b1101001001001011;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x0_LC_13_18_4  (
            .in0(N__16291),
            .in1(N__16207),
            .in2(N__14807),
            .in3(N__16867),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_13_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_13_18_5 .LUT_INIT=16'b0011010011111100;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_13_18_5  (
            .in0(N__14803),
            .in1(N__16285),
            .in2(N__15766),
            .in3(N__16167),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_c3_LC_13_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_c3_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_c3_LC_13_18_6 .LUT_INIT=16'b0111001100110001;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_c3_LC_13_18_6  (
            .in0(N__16286),
            .in1(N__14862),
            .in2(N__15767),
            .in3(N__14802),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_18_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__16290),
            .in2(N__14786),
            .in3(N__16169),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_2_1_9_LC_13_19_0 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_2_1_9_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_2_1_9_LC_13_19_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.sprites_addr_1_i_2_1_9_LC_13_19_0  (
            .in0(N__16816),
            .in1(N__17979),
            .in2(_gnd_net_),
            .in3(N__18098),
            .lcout(\this_ppu.sprites_addr_1_i_2_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_1 .LUT_INIT=16'b1000011101100000;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un54_sum_axb1_LC_13_19_1  (
            .in0(N__16065),
            .in1(N__15846),
            .in2(N__15983),
            .in3(N__15768),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_19_2 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x1_LC_13_19_2  (
            .in0(N__16202),
            .in1(N__16853),
            .in2(N__14930),
            .in3(N__16315),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_19_3 .LUT_INIT=16'b1001110000111001;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_x0_LC_13_19_3  (
            .in0(N__16316),
            .in1(N__16233),
            .in2(N__16868),
            .in3(N__16203),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_19_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_ns_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__14927),
            .in2(N__14921),
            .in3(N__16762),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1 ),
            .ltout(\this_vga_signals.mult1_un68_sum_axbxc3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_13_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_13_19_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_ac0_1_LC_13_19_5  (
            .in0(N__18097),
            .in1(N__16987),
            .in2(N__14912),
            .in3(N__14908),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_13_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_13_19_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_13_19_6  (
            .in0(N__16860),
            .in1(N__16318),
            .in2(N__16240),
            .in3(N__16763),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x1_LC_13_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x1_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x1_LC_13_19_7 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_x1_LC_13_19_7  (
            .in0(N__16317),
            .in1(N__16204),
            .in2(N__16869),
            .in3(N__14907),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_m1_0_LC_13_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_m1_0_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_m1_0_LC_13_20_4 .LUT_INIT=16'b0101101010011010;
    LogicCell40 \this_vga_signals.un3_haddress_if_m1_0_LC_13_20_4  (
            .in0(N__16205),
            .in1(N__14894),
            .in2(N__14879),
            .in3(N__14867),
            .lcout(\this_vga_signals.mult1_un68_sum_axb1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.pixel_clk_inferred_clock_RNO_LC_13_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.pixel_clk_inferred_clock_RNO_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.pixel_clk_inferred_clock_RNO_LC_13_20_6 .LUT_INIT=16'b0010010001000010;
    LogicCell40 \this_vga_signals.pixel_clk_inferred_clock_RNO_LC_13_20_6  (
            .in0(N__17801),
            .in1(N__15674),
            .in2(N__15665),
            .in3(N__17896),
            .lcout(M_this_vga_signals_pixel_clk_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_14_14_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__15542),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_M_vcounter_q_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24969),
            .ce(N__15524),
            .sr(N__15486));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFF6A3_5_LC_14_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFF6A3_5_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFF6A3_5_LC_14_15_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIFF6A3_5_LC_14_15_4  (
            .in0(N__15458),
            .in1(N__15264),
            .in2(N__15203),
            .in3(N__15128),
            .lcout(\this_vga_signals.N_455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGUM81_9_LC_14_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGUM81_9_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGUM81_9_LC_14_15_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGUM81_9_LC_14_15_6  (
            .in0(N__14944),
            .in1(N__15875),
            .in2(_gnd_net_),
            .in3(N__15976),
            .lcout(\this_vga_signals.N_459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_14_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_14_16_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIORPF_9_LC_14_16_1  (
            .in0(N__15876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15961),
            .lcout(\this_vga_signals.N_404_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_0_LC_14_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_0_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_0_LC_14_16_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_state_d_0_sqmuxa_i_0_0_o2_0_LC_14_16_3  (
            .in0(N__15774),
            .in1(N__16309),
            .in2(_gnd_net_),
            .in3(N__16056),
            .lcout(N_204_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIOT0S1_9_LC_14_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIOT0S1_9_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIOT0S1_9_LC_14_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIOT0S1_9_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__17029),
            .in2(_gnd_net_),
            .in3(N__17086),
            .lcout(\this_vga_signals.N_517_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_a3_1_9_LC_14_17_0 .C_ON=1'b1;
    defparam \this_ppu.sprites_addr_1_i_a3_1_9_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_a3_1_9_LC_14_17_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \this_ppu.sprites_addr_1_i_a3_1_9_LC_14_17_0  (
            .in0(N__17788),
            .in1(N__17881),
            .in2(N__17802),
            .in3(_gnd_net_),
            .lcout(\this_ppu.N_4_0_1 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_14_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_14_17_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_14_17_1  (
            .in0(N__17148),
            .in1(N__18067),
            .in2(_gnd_net_),
            .in3(N__14933),
            .lcout(this_vga_signals_M_hcounter_q_2),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_1_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_2 ),
            .clk(N__24984),
            .ce(),
            .sr(N__17056));
    defparam \this_vga_signals.M_hcounter_q_3_LC_14_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_14_17_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_14_17_2  (
            .in0(N__17140),
            .in1(N__16996),
            .in2(_gnd_net_),
            .in3(N__16115),
            .lcout(this_vga_signals_M_hcounter_q_3),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_1_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_3 ),
            .clk(N__24984),
            .ce(),
            .sr(N__17056));
    defparam \this_vga_signals.M_hcounter_q_4_LC_14_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_14_17_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_14_17_3  (
            .in0(N__17149),
            .in1(N__16198),
            .in2(_gnd_net_),
            .in3(N__16112),
            .lcout(this_vga_signals_M_hcounter_q_4),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_1_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_4 ),
            .clk(N__24984),
            .ce(),
            .sr(N__17056));
    defparam \this_vga_signals.M_hcounter_q_5_LC_14_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_14_17_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_14_17_4  (
            .in0(N__17141),
            .in1(N__16310),
            .in2(_gnd_net_),
            .in3(N__16109),
            .lcout(this_vga_signals_M_hcounter_q_5),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_1_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_5 ),
            .clk(N__24984),
            .ce(),
            .sr(N__17056));
    defparam \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUF_LC_14_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUF_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUF_LC_14_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUF_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__15765),
            .in2(_gnd_net_),
            .in3(N__16106),
            .lcout(\this_vga_signals.un1_M_hcounter_d_1_cry_5_c_RNIUHUFZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_1_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_7_LC_14_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_14_17_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_14_17_6  (
            .in0(N__17142),
            .in1(N__16062),
            .in2(_gnd_net_),
            .in3(N__16007),
            .lcout(this_vga_signals_M_hcounter_q_7),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_1_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_7 ),
            .clk(N__24984),
            .ce(),
            .sr(N__17056));
    defparam \this_vga_signals.M_hcounter_q_8_LC_14_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_14_17_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_14_17_7  (
            .in0(N__17150),
            .in1(N__15960),
            .in2(_gnd_net_),
            .in3(N__15896),
            .lcout(this_vga_signals_M_hcounter_q_8),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_1_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_1_cry_8 ),
            .clk(N__24984),
            .ce(),
            .sr(N__17056));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_14_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_14_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__15863),
            .in2(_gnd_net_),
            .in3(N__15893),
            .lcout(this_vga_signals_M_hcounter_q_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24989),
            .ce(N__15707),
            .sr(N__17055));
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_14_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_6_LC_14_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_6_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15805),
            .lcout(this_vga_signals_M_hcounter_q_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24989),
            .ce(N__15707),
            .sr(N__17055));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_14_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_14_19_0 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_14_19_0  (
            .in0(N__16214),
            .in1(N__16764),
            .in2(N__17000),
            .in3(N__15686),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_0_0_9_LC_14_19_1 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_0_0_9_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_0_0_9_LC_14_19_1 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \this_ppu.sprites_addr_1_i_0_0_9_LC_14_19_1  (
            .in0(N__23842),
            .in1(N__17953),
            .in2(N__16820),
            .in3(N__17928),
            .lcout(),
            .ltout(\this_ppu.sprites_addr_1_i_0_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_0_2_9_LC_14_19_2 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_0_2_9_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_0_2_9_LC_14_19_2 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \this_ppu.sprites_addr_1_i_0_2_9_LC_14_19_2  (
            .in0(N__17929),
            .in1(N__16508),
            .in2(N__16499),
            .in3(N__16496),
            .lcout(),
            .ltout(\this_ppu.sprites_addr_1_i_0_2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_0_9_LC_14_19_3 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_0_9_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_0_9_LC_14_19_3 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \this_ppu.sprites_addr_1_i_0_9_LC_14_19_3  (
            .in0(N__16787),
            .in1(N__17954),
            .in2(N__16484),
            .in3(N__16793),
            .lcout(N_138_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_ns_LC_14_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_ns_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_ns_LC_14_19_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un68_sum_axbxc3_ns_LC_14_19_4  (
            .in0(N__16373),
            .in1(N__16367),
            .in2(_gnd_net_),
            .in3(N__16361),
            .lcout(if_generate_plus_mult1_un68_sum_axbxc3_ns),
            .ltout(if_generate_plus_mult1_un68_sum_axbxc3_ns_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_14_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_14_19_5 .LUT_INIT=16'b1000011001111001;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_14_19_5  (
            .in0(N__16355),
            .in1(N__16986),
            .in2(N__16349),
            .in3(N__16727),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0),
            .ltout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m1_0_x1_LC_14_19_6 .C_ON=1'b0;
    defparam \this_ppu.sprites_m1_0_x1_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m1_0_x1_LC_14_19_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_ppu.sprites_m1_0_x1_LC_14_19_6  (
            .in0(N__18245),
            .in1(N__17190),
            .in2(N__16346),
            .in3(N__17172),
            .lcout(\this_ppu.sprites_m1_0_xZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m1_0_x0_LC_14_19_7 .C_ON=1'b0;
    defparam \this_ppu.sprites_m1_0_x0_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m1_0_x0_LC_14_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_ppu.sprites_m1_0_x0_LC_14_19_7  (
            .in0(N__17171),
            .in1(N__18244),
            .in2(N__17194),
            .in3(N__17927),
            .lcout(\this_ppu.sprites_m1_0_xZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_m7_0_x4_0_LC_14_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_m7_0_x4_0_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_m7_0_x4_0_LC_14_20_3 .LUT_INIT=16'b0100101111010010;
    LogicCell40 \this_vga_signals.un3_haddress_if_m7_0_x4_0_LC_14_20_3  (
            .in0(N__16870),
            .in1(N__16319),
            .in2(N__16241),
            .in3(N__16206),
            .lcout(),
            .ltout(\this_vga_signals.if_N_8_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_m7_0_m2_0_LC_14_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_m7_0_m2_0_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_m7_0_m2_0_LC_14_20_4 .LUT_INIT=16'b0011001110001110;
    LogicCell40 \this_vga_signals.un3_haddress_if_m7_0_m2_0_LC_14_20_4  (
            .in0(N__18082),
            .in1(N__16988),
            .in2(N__16730),
            .in3(N__16725),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un75_sum_c3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_m7_0_o4_LC_14_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_m7_0_o4_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_m7_0_o4_LC_14_20_6 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un3_haddress_if_m7_0_o4_LC_14_20_6  (
            .in0(N__18083),
            .in1(N__16726),
            .in2(N__17902),
            .in3(N__17170),
            .lcout(\this_vga_signals.if_N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_13_LC_14_21_1.C_ON=1'b0;
    defparam M_this_internal_address_q_13_LC_14_21_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_13_LC_14_21_1.LUT_INIT=16'b0011010100110000;
    LogicCell40 M_this_internal_address_q_13_LC_14_21_1 (
            .in0(N__25212),
            .in1(N__21242),
            .in2(N__21637),
            .in3(N__18911),
            .lcout(M_this_internal_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25002),
            .ce(),
            .sr(N__24739));
    defparam M_this_internal_address_q_7_LC_14_23_1.C_ON=1'b0;
    defparam M_this_internal_address_q_7_LC_14_23_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_7_LC_14_23_1.LUT_INIT=16'b0011010100110000;
    LogicCell40 M_this_internal_address_q_7_LC_14_23_1 (
            .in0(N__25213),
            .in1(N__18776),
            .in2(N__21638),
            .in3(N__18305),
            .lcout(M_this_internal_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25014),
            .ce(),
            .sr(N__24734));
    defparam CONSTANT_ONE_LUT4_LC_14_24_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_14_24_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_14_24_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_14_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4UBI1_9_LC_15_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4UBI1_9_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4UBI1_9_LC_15_15_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI4UBI1_9_LC_15_15_0  (
            .in0(N__16662),
            .in1(N__16712),
            .in2(_gnd_net_),
            .in3(N__16702),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI4UBI1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_15_15_1 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_15_15_1 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_15_15_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_15_15_1  (
            .in0(N__16703),
            .in1(N__16888),
            .in2(_gnd_net_),
            .in3(N__24785),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24970),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_RNIFKS8_0_LC_15_15_5 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_RNIFKS8_0_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \this_pixel_clk.M_counter_q_RNIFKS8_0_LC_15_15_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_RNIFKS8_0_LC_15_15_5  (
            .in0(N__16700),
            .in1(N__16887),
            .in2(_gnd_net_),
            .in3(N__24784),
            .lcout(M_counter_q_RNIFKS8_0),
            .ltout(M_counter_q_RNIFKS8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.G_210_LC_15_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.G_210_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.G_210_LC_15_15_6 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \this_vga_signals.G_210_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16706),
            .in3(N__16701),
            .lcout(\this_vga_signals.GZ0Z_210 ),
            .ltout(\this_vga_signals.GZ0Z_210_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIRV75_9_LC_15_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIRV75_9_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIRV75_9_LC_15_15_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIRV75_9_LC_15_15_7  (
            .in0(N__16688),
            .in1(N__16661),
            .in2(N__16646),
            .in3(N__16641),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNIIRV75Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_15_16_5 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_15_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16889),
            .lcout(\this_pixel_clk.M_counter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24974),
            .ce(),
            .sr(N__24742));
    defparam \this_sprites_ram.mem_radreg_11_LC_15_17_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_11_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_11_LC_15_17_0 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \this_sprites_ram.mem_radreg_11_LC_15_17_0  (
            .in0(N__23858),
            .in1(N__16778),
            .in2(N__16739),
            .in3(N__18287),
            .lcout(\this_sprites_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24978),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIG0MN6_7_LC_15_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIG0MN6_7_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIG0MN6_7_LC_15_17_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIG0MN6_7_LC_15_17_6  (
            .in0(N__23857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16874),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_15_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_15_18_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_15_18_0  (
            .in0(N__17200),
            .in1(N__17173),
            .in2(_gnd_net_),
            .in3(N__18247),
            .lcout(if_generate_plus_mult1_un75_sum_axbxc3),
            .ltout(if_generate_plus_mult1_un75_sum_axbxc3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un5_sprites_addr_1_ac0_1_LC_15_18_1 .C_ON=1'b0;
    defparam \this_ppu.un5_sprites_addr_1_ac0_1_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un5_sprites_addr_1_ac0_1_LC_15_18_1 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \this_ppu.un5_sprites_addr_1_ac0_1_LC_15_18_1  (
            .in0(N__23830),
            .in1(N__17966),
            .in2(N__16826),
            .in3(N__17933),
            .lcout(\this_ppu.un5_sprites_addr_1_c2 ),
            .ltout(\this_ppu.un5_sprites_addr_1_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un5_sprites_addr_1_ac0_5_LC_15_18_2 .C_ON=1'b0;
    defparam \this_ppu.un5_sprites_addr_1_ac0_5_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un5_sprites_addr_1_ac0_5_LC_15_18_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \this_ppu.un5_sprites_addr_1_ac0_5_LC_15_18_2  (
            .in0(N__16773),
            .in1(_gnd_net_),
            .in2(N__16823),
            .in3(N__18249),
            .lcout(\this_ppu.un5_sprites_addr_1_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_8_tz_9_LC_15_18_3 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_8_tz_9_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_8_tz_9_LC_15_18_3 .LUT_INIT=16'b0000111010101110;
    LogicCell40 \this_ppu.sprites_addr_1_i_8_tz_9_LC_15_18_3  (
            .in0(N__17996),
            .in1(N__16815),
            .in2(N__18093),
            .in3(N__17935),
            .lcout(\this_ppu.sprites_addr_1_i_7_tz_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_a7_9_LC_15_18_4 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_a7_9_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_a7_9_LC_15_18_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.sprites_addr_1_i_a7_9_LC_15_18_4  (
            .in0(N__17934),
            .in1(N__18062),
            .in2(_gnd_net_),
            .in3(N__17995),
            .lcout(\this_ppu.sprites_addr_1_i_a7Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un5_sprites_addr_1_axbxc3_LC_15_18_5 .C_ON=1'b0;
    defparam \this_ppu.un5_sprites_addr_1_axbxc3_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un5_sprites_addr_1_axbxc3_LC_15_18_5 .LUT_INIT=16'b1011000001000000;
    LogicCell40 \this_ppu.un5_sprites_addr_1_axbxc3_LC_15_18_5  (
            .in0(N__18250),
            .in1(N__18268),
            .in2(N__23856),
            .in3(N__16774),
            .lcout(\this_ppu.un5_sprites_addr1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_15_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_15_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un82_sum_axb1_LC_15_18_6  (
            .in0(N__17201),
            .in1(N__17174),
            .in2(N__18107),
            .in3(N__18248),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_axb1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_15_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_15_19_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_15_19_3  (
            .in0(N__17775),
            .in1(N__17119),
            .in2(_gnd_net_),
            .in3(N__17871),
            .lcout(this_vga_signals_M_hcounter_q_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24990),
            .ce(),
            .sr(N__17054));
    defparam \this_vga_signals.M_hcounter_q_0_LC_15_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_15_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_15_19_4  (
            .in0(N__17118),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17774),
            .lcout(this_vga_signals_M_hcounter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24990),
            .ce(),
            .sr(N__17054));
    defparam \this_vga_signals.un3_haddress_if_m7_0_m2_LC_15_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_m7_0_m2_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_m7_0_m2_LC_15_19_6 .LUT_INIT=16'b0001101100100111;
    LogicCell40 \this_vga_signals.un3_haddress_if_m7_0_m2_LC_15_19_6  (
            .in0(N__17001),
            .in1(N__16916),
            .in2(N__18101),
            .in3(N__18246),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3),
            .ltout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un82_sum_c3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m1_0_ns_LC_15_19_7 .C_ON=1'b0;
    defparam \this_ppu.sprites_m1_0_ns_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m1_0_ns_LC_15_19_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \this_ppu.sprites_m1_0_ns_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__16910),
            .in2(N__16904),
            .in3(N__16901),
            .lcout(this_ppu_sprites_N_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_2_LC_15_20_3.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_2_LC_15_20_3.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_2_LC_15_20_3.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_internal_address_q_RNO_0_2_LC_15_20_3 (
            .in0(N__21212),
            .in1(N__18471),
            .in2(N__22759),
            .in3(N__21975),
            .lcout(M_this_internal_address_q_3_ns_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_9_LC_15_20_4.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_9_LC_15_20_4.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_9_LC_15_20_4.LUT_INIT=16'b0000111100100111;
    LogicCell40 M_this_internal_address_q_RNO_0_9_LC_15_20_4 (
            .in0(N__21977),
            .in1(N__22754),
            .in2(N__19093),
            .in3(N__21214),
            .lcout(M_this_internal_address_q_3_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_8_LC_15_20_6.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_8_LC_15_20_6.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_8_LC_15_20_6.LUT_INIT=16'b0000001011011111;
    LogicCell40 M_this_internal_address_q_RNO_0_8_LC_15_20_6 (
            .in0(N__21976),
            .in1(N__21213),
            .in2(N__21035),
            .in3(N__19215),
            .lcout(M_this_internal_address_q_3_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_2_LC_15_21_1.C_ON=1'b0;
    defparam M_this_internal_address_q_2_LC_15_21_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_2_LC_15_21_1.LUT_INIT=16'b0100011101000100;
    LogicCell40 M_this_internal_address_q_2_LC_15_21_1 (
            .in0(N__16895),
            .in1(N__21601),
            .in2(N__25252),
            .in3(N__18452),
            .lcout(M_this_internal_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24997),
            .ce(),
            .sr(N__24737));
    defparam M_this_internal_address_q_9_LC_15_21_3.C_ON=1'b0;
    defparam M_this_internal_address_q_9_LC_15_21_3.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_9_LC_15_21_3.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_9_LC_15_21_3 (
            .in0(N__17225),
            .in1(N__25215),
            .in2(N__21626),
            .in3(N__19067),
            .lcout(M_this_internal_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24997),
            .ce(),
            .sr(N__24737));
    defparam M_this_internal_address_q_RNO_0_3_LC_15_21_4.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_3_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_3_LC_15_21_4.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_internal_address_q_RNO_0_3_LC_15_21_4 (
            .in0(N__21224),
            .in1(N__18342),
            .in2(N__23198),
            .in3(N__22021),
            .lcout(),
            .ltout(M_this_internal_address_q_3_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_3_LC_15_21_5.C_ON=1'b0;
    defparam M_this_internal_address_q_3_LC_15_21_5.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_3_LC_15_21_5.LUT_INIT=16'b0001101100001010;
    LogicCell40 M_this_internal_address_q_3_LC_15_21_5 (
            .in0(N__21602),
            .in1(N__25214),
            .in2(N__17219),
            .in3(N__18323),
            .lcout(M_this_internal_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24997),
            .ce(),
            .sr(N__24737));
    defparam M_this_internal_address_q_8_LC_15_21_6.C_ON=1'b0;
    defparam M_this_internal_address_q_8_LC_15_21_6.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_8_LC_15_21_6.LUT_INIT=16'b0011101000110000;
    LogicCell40 M_this_internal_address_q_8_LC_15_21_6 (
            .in0(N__21225),
            .in1(N__17216),
            .in2(N__21625),
            .in3(N__19196),
            .lcout(M_this_internal_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24997),
            .ce(),
            .sr(N__24737));
    defparam M_this_state_q_RNI20CE_0_LC_15_22_2.C_ON=1'b0;
    defparam M_this_state_q_RNI20CE_0_LC_15_22_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI20CE_0_LC_15_22_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 M_this_state_q_RNI20CE_0_LC_15_22_2 (
            .in0(_gnd_net_),
            .in1(N__25197),
            .in2(_gnd_net_),
            .in3(N__24798),
            .lcout(M_this_state_q_RNI20CEZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_15_23_0.C_ON=1'b1;
    defparam M_this_data_count_q_0_LC_15_23_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_15_23_0.LUT_INIT=16'b0011110000111100;
    LogicCell40 M_this_data_count_q_0_LC_15_23_0 (
            .in0(_gnd_net_),
            .in1(N__19556),
            .in2(N__23545),
            .in3(_gnd_net_),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(un1_M_this_data_count_q_cry_0),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_1_LC_15_23_1.C_ON=1'b1;
    defparam M_this_data_count_q_1_LC_15_23_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_15_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_1_LC_15_23_1 (
            .in0(_gnd_net_),
            .in1(N__23522),
            .in2(N__19388),
            .in3(N__17210),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_0),
            .carryout(un1_M_this_data_count_q_cry_1),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_2_LC_15_23_2.C_ON=1'b1;
    defparam M_this_data_count_q_2_LC_15_23_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_15_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_2_LC_15_23_2 (
            .in0(_gnd_net_),
            .in1(N__19415),
            .in2(N__23546),
            .in3(N__17207),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_1),
            .carryout(un1_M_this_data_count_q_cry_2),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_3_LC_15_23_3.C_ON=1'b1;
    defparam M_this_data_count_q_3_LC_15_23_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_15_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_3_LC_15_23_3 (
            .in0(_gnd_net_),
            .in1(N__23526),
            .in2(N__19430),
            .in3(N__17204),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_2),
            .carryout(un1_M_this_data_count_q_cry_3),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_4_LC_15_23_4.C_ON=1'b1;
    defparam M_this_data_count_q_4_LC_15_23_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_15_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_4_LC_15_23_4 (
            .in0(_gnd_net_),
            .in1(N__19442),
            .in2(N__23547),
            .in3(N__17252),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_3),
            .carryout(un1_M_this_data_count_q_cry_4),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_5_LC_15_23_5.C_ON=1'b1;
    defparam M_this_data_count_q_5_LC_15_23_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_15_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_5_LC_15_23_5 (
            .in0(_gnd_net_),
            .in1(N__23530),
            .in2(N__19475),
            .in3(N__17249),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_4),
            .carryout(un1_M_this_data_count_q_cry_5),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_6_LC_15_23_6.C_ON=1'b1;
    defparam M_this_data_count_q_6_LC_15_23_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_15_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_6_LC_15_23_6 (
            .in0(_gnd_net_),
            .in1(N__19487),
            .in2(N__23548),
            .in3(N__17246),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_5),
            .carryout(un1_M_this_data_count_q_cry_6),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_7_LC_15_23_7.C_ON=1'b1;
    defparam M_this_data_count_q_7_LC_15_23_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_15_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_7_LC_15_23_7 (
            .in0(_gnd_net_),
            .in1(N__23534),
            .in2(N__19460),
            .in3(N__17243),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_6),
            .carryout(un1_M_this_data_count_q_cry_7),
            .clk(N__25007),
            .ce(),
            .sr(N__17696));
    defparam M_this_data_count_q_8_LC_15_24_0.C_ON=1'b1;
    defparam M_this_data_count_q_8_LC_15_24_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_15_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_8_LC_15_24_0 (
            .in0(_gnd_net_),
            .in1(N__19513),
            .in2(N__23540),
            .in3(N__17240),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(un1_M_this_data_count_q_cry_8),
            .clk(N__25015),
            .ce(),
            .sr(N__17695));
    defparam M_this_data_count_q_9_LC_15_24_1.C_ON=1'b1;
    defparam M_this_data_count_q_9_LC_15_24_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_15_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_9_LC_15_24_1 (
            .in0(_gnd_net_),
            .in1(N__23505),
            .in2(N__19529),
            .in3(N__17237),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_8),
            .carryout(un1_M_this_data_count_q_cry_9),
            .clk(N__25015),
            .ce(),
            .sr(N__17695));
    defparam M_this_data_count_q_10_LC_15_24_2.C_ON=1'b1;
    defparam M_this_data_count_q_10_LC_15_24_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_15_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_10_LC_15_24_2 (
            .in0(_gnd_net_),
            .in1(N__19402),
            .in2(N__23541),
            .in3(N__17234),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_9),
            .carryout(un1_M_this_data_count_q_cry_10),
            .clk(N__25015),
            .ce(),
            .sr(N__17695));
    defparam M_this_data_count_q_11_LC_15_24_3.C_ON=1'b1;
    defparam M_this_data_count_q_11_LC_15_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_15_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_11_LC_15_24_3 (
            .in0(_gnd_net_),
            .in1(N__23509),
            .in2(N__19544),
            .in3(N__17231),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_10),
            .carryout(un1_M_this_data_count_q_cry_11),
            .clk(N__25015),
            .ce(),
            .sr(N__17695));
    defparam M_this_data_count_q_12_LC_15_24_4.C_ON=1'b1;
    defparam M_this_data_count_q_12_LC_15_24_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_15_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_12_LC_15_24_4 (
            .in0(_gnd_net_),
            .in1(N__19499),
            .in2(N__23542),
            .in3(N__17228),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_11),
            .carryout(un1_M_this_data_count_q_cry_12),
            .clk(N__25015),
            .ce(),
            .sr(N__17695));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_15_24_5.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_15_24_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_15_24_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_0_LC_15_24_5 (
            .in0(_gnd_net_),
            .in1(N__17346),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_15_24_6.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_15_24_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_15_24_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_1_LC_15_24_6 (
            .in0(_gnd_net_),
            .in1(N__17348),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12_THRU_CRY_0_THRU_CO),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_15_24_7.C_ON=1'b1;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_15_24_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_15_24_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_data_count_q_cry_12_c_THRU_CRY_2_LC_15_24_7 (
            .in0(_gnd_net_),
            .in1(N__17347),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_M_this_data_count_q_cry_12_THRU_CRY_1_THRU_CO),
            .carryout(un1_M_this_data_count_q_cry_12_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_15_25_0.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_15_25_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_15_25_0.LUT_INIT=16'b1110101110111110;
    LogicCell40 M_this_data_count_q_13_LC_15_25_0 (
            .in0(N__25251),
            .in1(N__23543),
            .in2(N__19571),
            .in3(N__17318),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25017),
            .ce(),
            .sr(N__24731));
    defparam \this_reset_cond.M_stage_q_3_LC_16_13_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_16_13_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_16_13_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_16_13_0  (
            .in0(N__19352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17315),
            .lcout(M_this_state_q_nss_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24965),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_16_13_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_16_13_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_16_13_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__19351),
            .in2(_gnd_net_),
            .in3(N__19319),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24965),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_13_LC_16_17_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_13_LC_16_17_1 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_13_LC_16_17_1 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \this_sprites_ram.mem_radreg_13_LC_16_17_1  (
            .in0(N__18286),
            .in1(N__17273),
            .in2(N__17302),
            .in3(N__17264),
            .lcout(\this_sprites_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24973),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_12_LC_16_17_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_12_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \this_sprites_ram.mem_radreg_12_LC_16_17_4 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \this_sprites_ram.mem_radreg_12_LC_16_17_4  (
            .in0(N__17272),
            .in1(N__17263),
            .in2(_gnd_net_),
            .in3(N__18285),
            .lcout(\this_sprites_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24973),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_16_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_16_18_3 .LUT_INIT=16'b1001101110001001;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_ac0_3_0_LC_16_18_3  (
            .in0(N__17870),
            .in1(N__17714),
            .in2(N__17795),
            .in3(N__19755),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0),
            .ltout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_c3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_LC_16_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_LC_16_18_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_LC_16_18_4  (
            .in0(N__19756),
            .in1(_gnd_net_),
            .in2(N__18290),
            .in3(N__23691),
            .lcout(if_generate_plus_mult1_un89_sum_axbxc3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m6_0_LC_16_19_0 .C_ON=1'b0;
    defparam \this_ppu.sprites_m6_0_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m6_0_LC_16_19_0 .LUT_INIT=16'b1001101101110110;
    LogicCell40 \this_ppu.sprites_m6_0_LC_16_19_0  (
            .in0(N__17869),
            .in1(N__17712),
            .in2(N__17800),
            .in3(N__19754),
            .lcout(),
            .ltout(\this_ppu.sprites_N_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m7_0_LC_16_19_1 .C_ON=1'b0;
    defparam \this_ppu.sprites_m7_0_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m7_0_LC_16_19_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \this_ppu.sprites_m7_0_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18272),
            .in3(N__23690),
            .lcout(),
            .ltout(\this_ppu.sprites_m7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.N_140_i_LC_16_19_2 .C_ON=1'b0;
    defparam \this_ppu.N_140_i_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.N_140_i_LC_16_19_2 .LUT_INIT=16'b0000100010100010;
    LogicCell40 \this_ppu.N_140_i_LC_16_19_2  (
            .in0(N__23859),
            .in1(N__18269),
            .in2(N__18257),
            .in3(N__18254),
            .lcout(N_140_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_16_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_16_19_4 .LUT_INIT=16'b1101010000101011;
    LogicCell40 \this_vga_signals.un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_16_19_4  (
            .in0(N__17952),
            .in1(N__18105),
            .in2(N__17889),
            .in3(N__17994),
            .lcout(this_vga_signals_un3_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m1_LC_16_19_5 .C_ON=1'b0;
    defparam \this_ppu.sprites_m1_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m1_LC_16_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_ppu.sprites_m1_LC_16_19_5  (
            .in0(N__17965),
            .in1(N__17951),
            .in2(_gnd_net_),
            .in3(N__17936),
            .lcout(),
            .ltout(\this_ppu.sprites_mZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m5_LC_16_19_6 .C_ON=1'b0;
    defparam \this_ppu.sprites_m5_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m5_LC_16_19_6 .LUT_INIT=16'b0101010111101000;
    LogicCell40 \this_ppu.sprites_m5_LC_16_19_6  (
            .in0(N__17865),
            .in1(N__17773),
            .in2(N__17717),
            .in3(N__17713),
            .lcout(\this_ppu.sprites_N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_10_LC_16_20_0.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_10_LC_16_20_0.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_10_LC_16_20_0.LUT_INIT=16'b0100011101010101;
    LogicCell40 M_this_internal_address_q_RNO_0_10_LC_16_20_0 (
            .in0(N__18951),
            .in1(N__21215),
            .in2(N__23194),
            .in3(N__22003),
            .lcout(),
            .ltout(M_this_internal_address_q_3_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_10_LC_16_20_1.C_ON=1'b0;
    defparam M_this_internal_address_q_10_LC_16_20_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_10_LC_16_20_1.LUT_INIT=16'b0001110100001100;
    LogicCell40 M_this_internal_address_q_10_LC_16_20_1 (
            .in0(N__25152),
            .in1(N__21583),
            .in2(N__17699),
            .in3(N__18932),
            .lcout(M_this_internal_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24985),
            .ce(),
            .sr(N__24736));
    defparam M_this_internal_address_q_RNO_1_0_LC_16_21_0.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_0_LC_16_21_0.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_0_LC_16_21_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_0_LC_16_21_0 (
            .in0(_gnd_net_),
            .in1(N__20011),
            .in2(N__20141),
            .in3(N__20140),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_0),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(un1_M_this_internal_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_1_LC_16_21_1.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_1_LC_16_21_1.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_1_LC_16_21_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_1_LC_16_21_1 (
            .in0(_gnd_net_),
            .in1(N__19861),
            .in2(_gnd_net_),
            .in3(N__18578),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_1),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_0),
            .carryout(un1_M_this_internal_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_2_LC_16_21_2.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_2_LC_16_21_2.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_2_LC_16_21_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_2_LC_16_21_2 (
            .in0(_gnd_net_),
            .in1(N__18472),
            .in2(_gnd_net_),
            .in3(N__18446),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_2),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_1),
            .carryout(un1_M_this_internal_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_3_LC_16_21_3.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_3_LC_16_21_3.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_3_LC_16_21_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_3_LC_16_21_3 (
            .in0(_gnd_net_),
            .in1(N__18346),
            .in2(_gnd_net_),
            .in3(N__18317),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_3),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_2),
            .carryout(un1_M_this_internal_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_4_LC_16_21_4.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_4_LC_16_21_4.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_4_LC_16_21_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_4_LC_16_21_4 (
            .in0(_gnd_net_),
            .in1(N__20269),
            .in2(_gnd_net_),
            .in3(N__18314),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_4),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_3),
            .carryout(un1_M_this_internal_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_5_LC_16_21_5.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_5_LC_16_21_5.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_5_LC_16_21_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_5_LC_16_21_5 (
            .in0(_gnd_net_),
            .in1(N__21406),
            .in2(_gnd_net_),
            .in3(N__18311),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_5),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_4),
            .carryout(un1_M_this_internal_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_6_LC_16_21_6.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_6_LC_16_21_6.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_6_LC_16_21_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_6_LC_16_21_6 (
            .in0(_gnd_net_),
            .in1(N__21279),
            .in2(_gnd_net_),
            .in3(N__18308),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_6),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_5),
            .carryout(un1_M_this_internal_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_7_LC_16_21_7.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_7_LC_16_21_7.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_7_LC_16_21_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_7_LC_16_21_7 (
            .in0(_gnd_net_),
            .in1(N__18808),
            .in2(_gnd_net_),
            .in3(N__18293),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_7),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_6),
            .carryout(un1_M_this_internal_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_8_LC_16_22_0.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_8_LC_16_22_0.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_8_LC_16_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_8_LC_16_22_0 (
            .in0(_gnd_net_),
            .in1(N__19216),
            .in2(_gnd_net_),
            .in3(N__19190),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_8),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(un1_M_this_internal_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_9_LC_16_22_1.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_9_LC_16_22_1.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_9_LC_16_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_9_LC_16_22_1 (
            .in0(_gnd_net_),
            .in1(N__19086),
            .in2(_gnd_net_),
            .in3(N__19061),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_9),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_8),
            .carryout(un1_M_this_internal_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_10_LC_16_22_2.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_10_LC_16_22_2.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_10_LC_16_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_10_LC_16_22_2 (
            .in0(_gnd_net_),
            .in1(N__18958),
            .in2(_gnd_net_),
            .in3(N__18923),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_10),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_9),
            .carryout(un1_M_this_internal_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_11_LC_16_22_3.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_11_LC_16_22_3.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_11_LC_16_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_11_LC_16_22_3 (
            .in0(_gnd_net_),
            .in1(N__24079),
            .in2(_gnd_net_),
            .in3(N__18920),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_11),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_10),
            .carryout(un1_M_this_internal_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_12_LC_16_22_4.C_ON=1'b1;
    defparam M_this_internal_address_q_RNO_1_12_LC_16_22_4.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_12_LC_16_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_internal_address_q_RNO_1_12_LC_16_22_4 (
            .in0(_gnd_net_),
            .in1(N__24169),
            .in2(_gnd_net_),
            .in3(N__18917),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_12),
            .ltout(),
            .carryin(un1_M_this_internal_address_q_cry_11),
            .carryout(un1_M_this_internal_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_1_13_LC_16_22_5.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_1_13_LC_16_22_5.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_1_13_LC_16_22_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_this_internal_address_q_RNO_1_13_LC_16_22_5 (
            .in0(_gnd_net_),
            .in1(N__24030),
            .in2(_gnd_net_),
            .in3(N__18914),
            .lcout(M_this_internal_address_q_RNO_1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_7_LC_16_23_0.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_7_LC_16_23_0.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_7_LC_16_23_0.LUT_INIT=16'b0010011100110011;
    LogicCell40 M_this_internal_address_q_RNO_0_7_LC_16_23_0 (
            .in0(N__21233),
            .in1(N__18801),
            .in2(N__20874),
            .in3(N__22028),
            .lcout(M_this_internal_address_q_3_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_0_LC_16_23_2.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_0_LC_16_23_2.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_0_LC_16_23_2.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_internal_address_q_RNO_0_0_LC_16_23_2 (
            .in0(N__21232),
            .in1(N__20004),
            .in2(N__20873),
            .in3(N__22027),
            .lcout(M_this_internal_address_q_3_ns_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam N_235_0_sbtinv_LC_16_23_4.C_ON=1'b0;
    defparam N_235_0_sbtinv_LC_16_23_4.SEQ_MODE=4'b0000;
    defparam N_235_0_sbtinv_LC_16_23_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 N_235_0_sbtinv_LC_16_23_4 (
            .in0(N__20192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_235_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIEOD9_13_LC_16_24_1.C_ON=1'b0;
    defparam M_this_data_count_q_RNIEOD9_13_LC_16_24_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIEOD9_13_LC_16_24_1.LUT_INIT=16'b0000000001010101;
    LogicCell40 M_this_data_count_q_RNIEOD9_13_LC_16_24_1 (
            .in0(N__19567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19555),
            .lcout(M_this_state_q_srsts_0_a2_1_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIAVRI_11_LC_16_24_2.C_ON=1'b0;
    defparam M_this_data_count_q_RNIAVRI_11_LC_16_24_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIAVRI_11_LC_16_24_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIAVRI_11_LC_16_24_2 (
            .in0(N__19540),
            .in1(N__19525),
            .in2(N__19514),
            .in3(N__19498),
            .lcout(M_this_state_q_srsts_0_a2_1_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIAQQL_4_LC_16_24_4.C_ON=1'b0;
    defparam M_this_data_count_q_RNIAQQL_4_LC_16_24_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIAQQL_4_LC_16_24_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIAQQL_4_LC_16_24_4 (
            .in0(N__19486),
            .in1(N__19471),
            .in2(N__19459),
            .in3(N__19441),
            .lcout(M_this_state_q_srsts_0_a2_1_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIBTAK_10_LC_16_24_5.C_ON=1'b0;
    defparam M_this_data_count_q_RNIBTAK_10_LC_16_24_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIBTAK_10_LC_16_24_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 M_this_data_count_q_RNIBTAK_10_LC_16_24_5 (
            .in0(N__19426),
            .in1(N__19414),
            .in2(N__19403),
            .in3(N__19384),
            .lcout(),
            .ltout(M_this_state_q_srsts_0_a2_1_8_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNIDFF62_10_LC_16_24_6.C_ON=1'b0;
    defparam M_this_data_count_q_RNIDFF62_10_LC_16_24_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNIDFF62_10_LC_16_24_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_data_count_q_RNIDFF62_10_LC_16_24_6 (
            .in0(N__19373),
            .in1(N__19367),
            .in2(N__19361),
            .in3(N__19358),
            .lcout(N_240),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_17_12_6  (
            .in0(N__19344),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24966),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_17_12_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_17_12_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__19345),
            .in2(_gnd_net_),
            .in3(N__19325),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24966),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_i_a2_0_3_LC_17_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_i_a2_0_3_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_i_a2_0_3_LC_17_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_i_i_a2_0_3_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(N__20448),
            .in2(_gnd_net_),
            .in3(N__22022),
            .lcout(N_476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o4_1_LC_17_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o4_1_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_o4_1_LC_17_19_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_i_o4_1_LC_17_19_0  (
            .in0(N__19799),
            .in1(N__20626),
            .in2(_gnd_net_),
            .in3(N__19828),
            .lcout(\this_vga_signals.N_224_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_addr_1_i_7_LC_17_19_3 .C_ON=1'b0;
    defparam \this_ppu.sprites_addr_1_i_7_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_addr_1_i_7_LC_17_19_3 .LUT_INIT=16'b1001000001100000;
    LogicCell40 \this_ppu.sprites_addr_1_i_7_LC_17_19_3  (
            .in0(N__23692),
            .in1(N__19766),
            .in2(N__23861),
            .in3(N__19760),
            .lcout(N_134_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_1_4_LC_17_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_1_4_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_1_4_LC_17_19_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_1_4_LC_17_19_4  (
            .in0(N__20487),
            .in1(N__19628),
            .in2(N__20549),
            .in3(N__19613),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_1_4_LC_17_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_1_4_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_1_4_LC_17_19_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_a2_0_1_4_LC_17_19_5  (
            .in0(N__23430),
            .in1(N__20449),
            .in2(N__20589),
            .in3(N__24790),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4 ),
            .ltout(\this_vga_signals.M_this_state_q_srsts_0_i_a2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_17_19_6.C_ON=1'b0;
    defparam M_this_state_q_4_LC_17_19_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_17_19_6.LUT_INIT=16'b0111000011111111;
    LogicCell40 M_this_state_q_4_LC_17_19_6 (
            .in0(N__24599),
            .in1(N__20600),
            .in2(N__19622),
            .in3(N__19619),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24991),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_4_LC_17_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_4_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_4_LC_17_20_2 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_0_4_LC_17_20_2  (
            .in0(N__19821),
            .in1(N__20147),
            .in2(N__19802),
            .in3(N__24788),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_17_20_3.C_ON=1'b0;
    defparam M_this_state_q_1_LC_17_20_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_17_20_3.LUT_INIT=16'b0101010101010100;
    LogicCell40 M_this_state_q_1_LC_17_20_3 (
            .in0(N__24789),
            .in1(N__25153),
            .in2(N__19607),
            .in3(N__23431),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24995),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_17_20_4.C_ON=1'b0;
    defparam M_this_state_q_0_LC_17_20_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_17_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_state_q_0_LC_17_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19598),
            .lcout(M_this_state_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24995),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.port_nmib_i_o2_LC_17_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.port_nmib_i_o2_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.port_nmib_i_o2_LC_17_20_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.port_nmib_i_o2_LC_17_20_7  (
            .in0(N__23407),
            .in1(N__19794),
            .in2(_gnd_net_),
            .in3(N__20447),
            .lcout(N_235_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_1_LC_17_21_0.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_1_LC_17_21_0.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_1_LC_17_21_0.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_internal_address_q_RNO_0_1_LC_17_21_0 (
            .in0(N__21223),
            .in1(N__19860),
            .in2(N__21043),
            .in3(N__22042),
            .lcout(M_this_internal_address_q_3_ns_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_2_4_LC_17_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_2_4_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_a2_2_4_LC_17_21_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_a2_2_4_LC_17_21_1  (
            .in0(N__22041),
            .in1(N__20167),
            .in2(N__25196),
            .in3(N__24786),
            .lcout(\this_vga_signals.N_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un19_i_i_i_a2_LC_17_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un19_i_i_i_a2_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un19_i_i_i_a2_LC_17_21_2 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \this_vga_signals.un19_i_i_i_a2_LC_17_21_2  (
            .in0(N__19798),
            .in1(N__22072),
            .in2(N__20591),
            .in3(N__22040),
            .lcout(un19_i_i_i_a2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_11_LC_17_22_7.C_ON=1'b0;
    defparam M_this_internal_address_q_11_LC_17_22_7.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_11_LC_17_22_7.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_11_LC_17_22_7 (
            .in0(N__20390),
            .in1(N__25159),
            .in2(N__21636),
            .in3(N__20126),
            .lcout(M_this_internal_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25003),
            .ce(),
            .sr(N__24735));
    defparam M_this_internal_address_q_0_LC_17_23_0.C_ON=1'b0;
    defparam M_this_internal_address_q_0_LC_17_23_0.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_0_LC_17_23_0.LUT_INIT=16'b0101000001011100;
    LogicCell40 M_this_internal_address_q_0_LC_17_23_0 (
            .in0(N__20120),
            .in1(N__20114),
            .in2(N__21633),
            .in3(N__25161),
            .lcout(M_this_internal_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25008),
            .ce(),
            .sr(N__24732));
    defparam M_this_internal_address_q_1_LC_17_23_6.C_ON=1'b0;
    defparam M_this_internal_address_q_1_LC_17_23_6.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_1_LC_17_23_6.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_1_LC_17_23_6 (
            .in0(N__19985),
            .in1(N__25160),
            .in2(N__21634),
            .in3(N__19976),
            .lcout(M_this_internal_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25008),
            .ce(),
            .sr(N__24732));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_a2_1_0_LC_18_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_a2_1_0_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_a2_1_0_LC_18_18_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_a2_1_0_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__19835),
            .in2(_gnd_net_),
            .in3(N__21114),
            .lcout(\this_vga_signals.N_479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_a2_2_LC_18_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_a2_2_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_i_a2_2_LC_18_19_0 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_i_a2_2_LC_18_19_0  (
            .in0(N__20446),
            .in1(N__19800),
            .in2(N__20630),
            .in3(N__19829),
            .lcout(),
            .ltout(\this_vga_signals.N_343_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_18_19_1.C_ON=1'b0;
    defparam M_this_state_q_2_LC_18_19_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_18_19_1.LUT_INIT=16'b0000000000001011;
    LogicCell40 M_this_state_q_2_LC_18_19_1 (
            .in0(N__19801),
            .in1(N__22053),
            .in2(N__19769),
            .in3(N__24799),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24996),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_a4_LC_18_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_a4_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_a4_LC_18_19_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_a4_LC_18_19_7  (
            .in0(N__21113),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20445),
            .lcout(\this_vga_signals.N_483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_18_20_3.C_ON=1'b0;
    defparam M_this_state_q_3_LC_18_20_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_18_20_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 M_this_state_q_3_LC_18_20_3 (
            .in0(_gnd_net_),
            .in1(N__20450),
            .in2(_gnd_net_),
            .in3(N__22031),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24998),
            .ce(),
            .sr(N__24741));
    defparam M_this_internal_address_q_5_LC_18_21_2.C_ON=1'b0;
    defparam M_this_internal_address_q_5_LC_18_21_2.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_5_LC_18_21_2.LUT_INIT=16'b0011101000110000;
    LogicCell40 M_this_internal_address_q_5_LC_18_21_2 (
            .in0(N__21196),
            .in1(N__21380),
            .in2(N__21566),
            .in3(N__20417),
            .lcout(M_this_internal_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25004),
            .ce(),
            .sr(N__24740));
    defparam M_this_internal_address_q_6_LC_18_21_3.C_ON=1'b0;
    defparam M_this_internal_address_q_6_LC_18_21_3.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_6_LC_18_21_3.LUT_INIT=16'b0010111000001100;
    LogicCell40 M_this_internal_address_q_6_LC_18_21_3 (
            .in0(N__21197),
            .in1(N__21541),
            .in2(N__21251),
            .in3(N__20408),
            .lcout(M_this_internal_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25004),
            .ce(),
            .sr(N__24740));
    defparam M_this_internal_address_q_12_LC_18_22_1.C_ON=1'b0;
    defparam M_this_internal_address_q_12_LC_18_22_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_12_LC_18_22_1.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_12_LC_18_22_1 (
            .in0(N__21122),
            .in1(N__25220),
            .in2(N__21612),
            .in3(N__20399),
            .lcout(M_this_internal_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25009),
            .ce(),
            .sr(N__24738));
    defparam M_this_internal_address_q_RNO_0_4_LC_18_23_2.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_4_LC_18_23_2.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_4_LC_18_23_2.LUT_INIT=16'b0001001110110011;
    LogicCell40 M_this_internal_address_q_RNO_0_4_LC_18_23_2 (
            .in0(N__22036),
            .in1(N__20259),
            .in2(N__21231),
            .in3(N__20823),
            .lcout(M_this_internal_address_q_3_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_11_LC_18_23_5.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_11_LC_18_23_5.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_11_LC_18_23_5.LUT_INIT=16'b0100011101010101;
    LogicCell40 M_this_internal_address_q_RNO_0_11_LC_18_23_5 (
            .in0(N__24080),
            .in1(N__21219),
            .in2(N__20827),
            .in3(N__22035),
            .lcout(M_this_internal_address_q_3_ns_1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_4_LC_18_24_1.C_ON=1'b0;
    defparam M_this_internal_address_q_4_LC_18_24_1.SEQ_MODE=4'b1000;
    defparam M_this_internal_address_q_4_LC_18_24_1.LUT_INIT=16'b0101001101010000;
    LogicCell40 M_this_internal_address_q_4_LC_18_24_1 (
            .in0(N__20384),
            .in1(N__25219),
            .in2(N__21635),
            .in3(N__20378),
            .lcout(M_this_internal_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25018),
            .ce(),
            .sr(N__24733));
    defparam \this_vga_signals.M_this_vram_write_data_0_i_1_LC_19_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_1_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_1_LC_19_14_3 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \this_vga_signals.M_this_vram_write_data_0_i_1_LC_19_14_3  (
            .in0(N__23500),
            .in1(N__21752),
            .in2(N__21042),
            .in3(N__22404),
            .lcout(M_this_vram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o4_4_4_LC_19_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o4_4_4_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o4_4_4_LC_19_19_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_o4_4_4_LC_19_19_4  (
            .in0(N__20699),
            .in1(N__20678),
            .in2(N__20660),
            .in3(N__20625),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4 ),
            .ltout(\this_vga_signals.M_this_state_q_srsts_0_i_o4_4Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_2_7_LC_19_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_2_7_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_2_7_LC_19_19_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_2_7_LC_19_19_5  (
            .in0(N__24595),
            .in1(N__20590),
            .in2(N__20561),
            .in3(N__24791),
            .lcout(\this_vga_signals.N_490 ),
            .ltout(\this_vga_signals.N_490_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_0_7_LC_19_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_0_7_LC_19_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_0_7_LC_19_19_6 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_0_7_LC_19_19_6  (
            .in0(N__20545),
            .in1(N__20507),
            .in2(N__20558),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_vga_signals.N_386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_19_19_7.C_ON=1'b0;
    defparam M_this_state_q_7_LC_19_19_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_19_19_7.LUT_INIT=16'b1111000011110010;
    LogicCell40 M_this_state_q_7_LC_19_19_7 (
            .in0(N__21116),
            .in1(N__22052),
            .in2(N__20555),
            .in3(N__24792),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24999),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_internal_address_q_3_ss0_i_a3_0_a2_LC_19_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_internal_address_q_3_ss0_i_a3_0_a2_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_internal_address_q_3_ss0_i_a3_0_a2_LC_19_20_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_internal_address_q_3_ss0_i_a3_0_a2_LC_19_20_0  (
            .in0(_gnd_net_),
            .in1(N__21660),
            .in2(_gnd_net_),
            .in3(N__25154),
            .lcout(N_355),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_6_LC_19_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_6_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_6_LC_19_20_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_6_LC_19_20_2  (
            .in0(N__24794),
            .in1(N__21649),
            .in2(_gnd_net_),
            .in3(N__22030),
            .lcout(),
            .ltout(\this_vga_signals.N_387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_19_20_3.C_ON=1'b0;
    defparam M_this_state_q_6_LC_19_20_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_19_20_3.LUT_INIT=16'b1111000011111000;
    LogicCell40 M_this_state_q_6_LC_19_20_3 (
            .in0(N__20459),
            .in1(N__20506),
            .in2(N__20552),
            .in3(N__20544),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25005),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_5_LC_19_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_5_LC_19_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_5_LC_19_20_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_0_a2_5_LC_19_20_5  (
            .in0(N__21661),
            .in1(N__22029),
            .in2(_gnd_net_),
            .in3(N__24793),
            .lcout(),
            .ltout(\this_vga_signals.N_391_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_19_20_6.C_ON=1'b0;
    defparam M_this_state_q_5_LC_19_20_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_19_20_6.LUT_INIT=16'b1111000111110000;
    LogicCell40 M_this_state_q_5_LC_19_20_6 (
            .in0(N__20543),
            .in1(N__20505),
            .in2(N__20462),
            .in3(N__20458),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25005),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_internal_address_q_3s2_i_0_LC_19_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_internal_address_q_3s2_i_0_LC_19_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_internal_address_q_3s2_i_0_LC_19_20_7 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \this_vga_signals.M_this_internal_address_q_3s2_i_0_LC_19_20_7  (
            .in0(N__25155),
            .in1(_gnd_net_),
            .in2(N__21665),
            .in3(N__21650),
            .lcout(N_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_5_LC_19_21_0.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_5_LC_19_21_0.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_5_LC_19_21_0.LUT_INIT=16'b0001101100110011;
    LogicCell40 M_this_internal_address_q_RNO_0_5_LC_19_21_0 (
            .in0(N__21170),
            .in1(N__21399),
            .in2(N__21091),
            .in3(N__22044),
            .lcout(M_this_internal_address_q_3_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_6_LC_19_21_3.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_6_LC_19_21_3.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_6_LC_19_21_3.LUT_INIT=16'b0000011110001111;
    LogicCell40 M_this_internal_address_q_RNO_0_6_LC_19_21_3 (
            .in0(N__22045),
            .in1(N__21171),
            .in2(N__21280),
            .in3(N__22711),
            .lcout(M_this_internal_address_q_3_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_13_LC_19_21_6.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_13_LC_19_21_6.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_13_LC_19_21_6.LUT_INIT=16'b0100011101010101;
    LogicCell40 M_this_internal_address_q_RNO_0_13_LC_19_21_6 (
            .in0(N__23988),
            .in1(N__21169),
            .in2(N__22712),
            .in3(N__22043),
            .lcout(M_this_internal_address_q_3_ns_1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_internal_address_q_RNO_0_12_LC_19_22_1.C_ON=1'b0;
    defparam M_this_internal_address_q_RNO_0_12_LC_19_22_1.SEQ_MODE=4'b0000;
    defparam M_this_internal_address_q_RNO_0_12_LC_19_22_1.LUT_INIT=16'b0000001011011111;
    LogicCell40 M_this_internal_address_q_RNO_0_12_LC_19_22_1 (
            .in0(N__22054),
            .in1(N__21198),
            .in2(N__21092),
            .in3(N__24160),
            .lcout(M_this_internal_address_q_3_ns_1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_a2_2_0_LC_20_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_a2_2_0_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_a2_2_0_LC_20_18_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_a2_2_0_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(N__22026),
            .in2(_gnd_net_),
            .in3(N__21115),
            .lcout(\this_vga_signals.N_481 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_1_LC_21_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_1_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_1_LC_21_18_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_i_1_LC_21_18_7  (
            .in0(N__21078),
            .in1(N__22779),
            .in2(N__21047),
            .in3(N__24344),
            .lcout(M_this_sprites_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_0_LC_21_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_0_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_0_LC_21_20_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_i_0_LC_21_20_5  (
            .in0(N__20881),
            .in1(N__22788),
            .in2(N__20831),
            .in3(N__24354),
            .lcout(M_this_sprites_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_vram_write_data_0_i_2_LC_22_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_2_LC_22_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_2_LC_22_13_7 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \this_vga_signals.M_this_vram_write_data_0_i_2_LC_22_13_7  (
            .in0(N__23536),
            .in1(N__21761),
            .in2(N__22766),
            .in3(N__22411),
            .lcout(M_this_vram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_22_18_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_22_18_5 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_0_12_LC_22_18_5  (
            .in0(N__22270),
            .in1(N__22124),
            .in2(N__22212),
            .in3(N__21671),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_23_13_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_23_13_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_23_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_LC_23_13_4  (
            .in0(N__22910),
            .in1(N__21800),
            .in2(_gnd_net_),
            .in3(N__21779),
            .lcout(),
            .ltout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_23_13_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_23_13_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_23_13_5 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_0_12_LC_23_13_5  (
            .in0(N__22211),
            .in1(N__22268),
            .in2(N__21767),
            .in3(N__22544),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_23_13_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_23_13_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_23_13_6 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_0_11_LC_23_13_6  (
            .in0(N__22484),
            .in1(N__22269),
            .in2(N__21764),
            .in3(N__22610),
            .lcout(M_this_sprites_ram_read_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_23_14_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_23_14_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_23_14_5 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI1MK12_12_LC_23_14_5  (
            .in0(N__22298),
            .in1(N__22421),
            .in2(N__22217),
            .in3(N__22577),
            .lcout(),
            .ltout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_23_14_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_23_14_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIAJNR3_11_LC_23_14_6  (
            .in0(N__22299),
            .in1(N__22454),
            .in2(N__21755),
            .in3(N__21710),
            .lcout(M_this_sprites_ram_read_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_23_14_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_23_14_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_23_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_0_LC_23_14_7  (
            .in0(N__22907),
            .in1(N__21743),
            .in2(_gnd_net_),
            .in3(N__21728),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_23_17_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_23_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_LC_23_17_1  (
            .in0(N__22855),
            .in1(N__21704),
            .in2(_gnd_net_),
            .in3(N__21692),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_23_17_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_23_17_3 .LUT_INIT=16'b1110001100100011;
    LogicCell40 \this_sprites_ram.mem_radreg_RNIIJNR3_11_LC_23_17_3  (
            .in0(N__23219),
            .in1(N__22157),
            .in2(N__22300),
            .in3(N__23009),
            .lcout(),
            .ltout(M_this_sprites_ram_read_data_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_vram_write_data_0_i_3_LC_23_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_3_LC_23_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_vram_write_data_0_i_3_LC_23_17_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \this_vga_signals.M_this_vram_write_data_0_i_3_LC_23_17_4  (
            .in0(N__23193),
            .in1(N__23470),
            .in2(N__22415),
            .in3(N__22412),
            .lcout(M_this_vram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_23_18_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_23_18_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_sprites_ram.mem_radreg_RNI5MK12_12_LC_23_18_0  (
            .in0(N__22285),
            .in1(N__22949),
            .in2(N__22213),
            .in3(N__22982),
            .lcout(\this_sprites_ram.mem_DOUT_7_i_m2_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_18_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_LC_23_18_3  (
            .in0(N__22895),
            .in1(N__22151),
            .in2(_gnd_net_),
            .in3(N__22139),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_23_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_23_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_RNILA4P_LC_23_19_2  (
            .in0(N__22118),
            .in1(N__22106),
            .in2(_gnd_net_),
            .in3(N__22898),
            .lcout(\this_sprites_ram.mem_mem_1_0_RNILA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_LC_23_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_LC_23_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_LC_23_19_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_sn_m2_0_LC_23_19_7  (
            .in0(_gnd_net_),
            .in1(N__22073),
            .in2(_gnd_net_),
            .in3(N__22055),
            .lcout(N_24_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_22_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_7_0_wclke_3_LC_23_22_2  (
            .in0(N__24173),
            .in1(N__24094),
            .in2(N__24041),
            .in3(N__23918),
            .lcout(\this_sprites_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_11_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_11_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_11_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_wclke_3_LC_24_11_6  (
            .in0(N__24207),
            .in1(N__24130),
            .in2(N__24051),
            .in3(N__23941),
            .lcout(\this_sprites_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_11_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_11_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_11_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_wclke_3_LC_24_11_7  (
            .in0(N__23942),
            .in1(N__24034),
            .in2(N__24134),
            .in3(N__24208),
            .lcout(\this_sprites_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_12_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_12_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_12_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_sprites_ram.mem_mem_1_0_wclke_3_LC_24_12_1  (
            .in0(N__24129),
            .in1(N__24209),
            .in2(N__24052),
            .in3(N__23940),
            .lcout(\this_sprites_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_24_12_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_24_12_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_24_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_LC_24_12_3  (
            .in0(N__22637),
            .in1(N__22622),
            .in2(_gnd_net_),
            .in3(N__22916),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_24_13_1 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_24_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_0_RNIJ62P_0_LC_24_13_1  (
            .in0(N__22914),
            .in1(N__22604),
            .in2(_gnd_net_),
            .in3(N__22592),
            .lcout(\this_sprites_ram.mem_mem_0_0_RNIJ62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_24_13_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_24_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_LC_24_13_3  (
            .in0(N__22915),
            .in1(N__22571),
            .in2(_gnd_net_),
            .in3(N__22559),
            .lcout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_wclke_3_LC_24_13_6  (
            .in0(N__24206),
            .in1(N__24120),
            .in2(N__24053),
            .in3(N__23931),
            .lcout(\this_sprites_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_24_14_0 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_24_14_0 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_24_14_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_LC_24_14_0  (
            .in0(N__22906),
            .in1(N__22514),
            .in2(_gnd_net_),
            .in3(N__22496),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_24_14_5 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_24_14_5 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_24_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_0_LC_24_14_5  (
            .in0(N__22478),
            .in1(N__22460),
            .in2(_gnd_net_),
            .in3(N__22905),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_24_14_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_24_14_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_24_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_0_RNINE6P_0_LC_24_14_6  (
            .in0(N__22904),
            .in1(N__22448),
            .in2(_gnd_net_),
            .in3(N__22433),
            .lcout(\this_sprites_ram.mem_mem_2_0_RNINE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_24_17_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_24_17_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_24_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_3_1_RNIRI8P_0_LC_24_17_2  (
            .in0(N__22909),
            .in1(N__23246),
            .in2(_gnd_net_),
            .in3(N__23228),
            .lcout(\this_sprites_ram.mem_mem_3_1_RNIRI8PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_4_0_wclke_3_LC_24_17_3  (
            .in0(N__24194),
            .in1(N__24103),
            .in2(N__24056),
            .in3(N__23919),
            .lcout(\this_sprites_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_3_LC_24_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_3_LC_24_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_3_LC_24_17_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_i_3_LC_24_17_6  (
            .in0(N__23192),
            .in1(N__22795),
            .in2(N__23129),
            .in3(N__24359),
            .lcout(M_this_sprites_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_17_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_17_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_17_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_1_1_RNINA4P_0_LC_24_17_7  (
            .in0(N__23036),
            .in1(N__23024),
            .in2(_gnd_net_),
            .in3(N__22908),
            .lcout(\this_sprites_ram.mem_mem_1_1_RNINA4PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_7 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_7 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_sprites_ram.mem_mem_0_1_RNIL62P_0_LC_24_18_7  (
            .in0(N__23003),
            .in1(N__22894),
            .in2(_gnd_net_),
            .in3(N__22988),
            .lcout(\this_sprites_ram.mem_mem_0_1_RNIL62PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_19_2 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_19_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_sprites_ram.mem_mem_2_1_RNIPE6P_0_LC_24_19_2  (
            .in0(N__22896),
            .in1(N__22976),
            .in2(_gnd_net_),
            .in3(N__22964),
            .lcout(\this_sprites_ram.mem_mem_2_1_RNIPE6PZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_19_3 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_19_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_sprites_ram.mem_mem_3_0_RNIPI8P_LC_24_19_3  (
            .in0(N__22943),
            .in1(N__22928),
            .in2(_gnd_net_),
            .in3(N__22897),
            .lcout(\this_sprites_ram.mem_mem_3_0_RNIPI8PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_2_LC_24_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_2_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_sprites_ram_write_data_1_i_2_LC_24_20_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \this_vga_signals.M_this_sprites_ram_write_data_1_i_2_LC_24_20_2  (
            .in0(N__22799),
            .in1(N__22755),
            .in2(N__22699),
            .in3(N__24358),
            .lcout(M_this_sprites_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_22_4 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_22_4 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_22_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_5_0_wclke_3_LC_24_22_4  (
            .in0(N__24174),
            .in1(N__24095),
            .in2(N__24055),
            .in3(N__23929),
            .lcout(\this_sprites_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_22_6 .C_ON=1'b0;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_22_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_sprites_ram.mem_mem_6_0_wclke_3_LC_24_22_6  (
            .in0(N__24175),
            .in1(N__24096),
            .in2(N__24054),
            .in3(N__23930),
            .lcout(\this_sprites_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.sprites_m7_LC_24_31_7 .C_ON=1'b0;
    defparam \this_ppu.sprites_m7_LC_24_31_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.sprites_m7_LC_24_31_7 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \this_ppu.sprites_m7_LC_24_31_7  (
            .in0(N__23855),
            .in1(N__23702),
            .in2(_gnd_net_),
            .in3(N__23669),
            .lcout(sprites_m7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_external_address_q_0_LC_31_23_0.C_ON=1'b1;
    defparam M_this_external_address_q_0_LC_31_23_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_0_LC_31_23_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_0_LC_31_23_0 (
            .in0(N__25253),
            .in1(N__23347),
            .in2(N__23544),
            .in3(N__23535),
            .lcout(M_this_external_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_31_23_0_),
            .carryout(un1_M_this_external_address_q_cry_0),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_1_LC_31_23_1.C_ON=1'b1;
    defparam M_this_external_address_q_1_LC_31_23_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_1_LC_31_23_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_1_LC_31_23_1 (
            .in0(N__25261),
            .in1(N__23329),
            .in2(_gnd_net_),
            .in3(N__23318),
            .lcout(M_this_external_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_0),
            .carryout(un1_M_this_external_address_q_cry_1),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_2_LC_31_23_2.C_ON=1'b1;
    defparam M_this_external_address_q_2_LC_31_23_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_2_LC_31_23_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_2_LC_31_23_2 (
            .in0(N__25254),
            .in1(N__23299),
            .in2(_gnd_net_),
            .in3(N__23288),
            .lcout(M_this_external_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_1),
            .carryout(un1_M_this_external_address_q_cry_2),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_3_LC_31_23_3.C_ON=1'b1;
    defparam M_this_external_address_q_3_LC_31_23_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_3_LC_31_23_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_3_LC_31_23_3 (
            .in0(N__25262),
            .in1(N__23275),
            .in2(_gnd_net_),
            .in3(N__23264),
            .lcout(M_this_external_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_2),
            .carryout(un1_M_this_external_address_q_cry_3),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_4_LC_31_23_4.C_ON=1'b1;
    defparam M_this_external_address_q_4_LC_31_23_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_4_LC_31_23_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_4_LC_31_23_4 (
            .in0(N__25255),
            .in1(N__23257),
            .in2(_gnd_net_),
            .in3(N__24566),
            .lcout(M_this_external_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_3),
            .carryout(un1_M_this_external_address_q_cry_4),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_5_LC_31_23_5.C_ON=1'b1;
    defparam M_this_external_address_q_5_LC_31_23_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_5_LC_31_23_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_5_LC_31_23_5 (
            .in0(N__25263),
            .in1(N__24556),
            .in2(_gnd_net_),
            .in3(N__24545),
            .lcout(M_this_external_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_4),
            .carryout(un1_M_this_external_address_q_cry_5),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_6_LC_31_23_6.C_ON=1'b1;
    defparam M_this_external_address_q_6_LC_31_23_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_6_LC_31_23_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_6_LC_31_23_6 (
            .in0(N__25256),
            .in1(N__24535),
            .in2(_gnd_net_),
            .in3(N__24524),
            .lcout(M_this_external_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_5),
            .carryout(un1_M_this_external_address_q_cry_6),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_7_LC_31_23_7.C_ON=1'b1;
    defparam M_this_external_address_q_7_LC_31_23_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_7_LC_31_23_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_7_LC_31_23_7 (
            .in0(N__25264),
            .in1(N__24508),
            .in2(_gnd_net_),
            .in3(N__24497),
            .lcout(M_this_external_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_6),
            .carryout(un1_M_this_external_address_q_cry_7),
            .clk(N__25034),
            .ce(),
            .sr(N__24745));
    defparam M_this_external_address_q_8_LC_31_24_0.C_ON=1'b1;
    defparam M_this_external_address_q_8_LC_31_24_0.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_8_LC_31_24_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_8_LC_31_24_0 (
            .in0(N__25260),
            .in1(N__24478),
            .in2(_gnd_net_),
            .in3(N__24467),
            .lcout(M_this_external_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_31_24_0_),
            .carryout(un1_M_this_external_address_q_cry_8),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam M_this_external_address_q_9_LC_31_24_1.C_ON=1'b1;
    defparam M_this_external_address_q_9_LC_31_24_1.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_9_LC_31_24_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_9_LC_31_24_1 (
            .in0(N__25276),
            .in1(N__24448),
            .in2(_gnd_net_),
            .in3(N__24437),
            .lcout(M_this_external_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_8),
            .carryout(un1_M_this_external_address_q_cry_9),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam M_this_external_address_q_10_LC_31_24_2.C_ON=1'b1;
    defparam M_this_external_address_q_10_LC_31_24_2.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_10_LC_31_24_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_10_LC_31_24_2 (
            .in0(N__25257),
            .in1(N__24418),
            .in2(_gnd_net_),
            .in3(N__24407),
            .lcout(M_this_external_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_9),
            .carryout(un1_M_this_external_address_q_cry_10),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam M_this_external_address_q_11_LC_31_24_3.C_ON=1'b1;
    defparam M_this_external_address_q_11_LC_31_24_3.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_11_LC_31_24_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_11_LC_31_24_3 (
            .in0(N__25274),
            .in1(N__24391),
            .in2(_gnd_net_),
            .in3(N__24380),
            .lcout(M_this_external_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_10),
            .carryout(un1_M_this_external_address_q_cry_11),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam M_this_external_address_q_12_LC_31_24_4.C_ON=1'b1;
    defparam M_this_external_address_q_12_LC_31_24_4.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_12_LC_31_24_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_12_LC_31_24_4 (
            .in0(N__25258),
            .in1(N__24373),
            .in2(_gnd_net_),
            .in3(N__24362),
            .lcout(M_this_external_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_11),
            .carryout(un1_M_this_external_address_q_cry_12),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam M_this_external_address_q_13_LC_31_24_5.C_ON=1'b1;
    defparam M_this_external_address_q_13_LC_31_24_5.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_13_LC_31_24_5.LUT_INIT=16'b1011101111101110;
    LogicCell40 M_this_external_address_q_13_LC_31_24_5 (
            .in0(N__25275),
            .in1(N__25315),
            .in2(_gnd_net_),
            .in3(N__25304),
            .lcout(M_this_external_address_qZ0Z_13),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_12),
            .carryout(un1_M_this_external_address_q_cry_13),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam M_this_external_address_q_14_LC_31_24_6.C_ON=1'b1;
    defparam M_this_external_address_q_14_LC_31_24_6.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_14_LC_31_24_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_external_address_q_14_LC_31_24_6 (
            .in0(N__25259),
            .in1(N__25291),
            .in2(_gnd_net_),
            .in3(N__25280),
            .lcout(M_this_external_address_qZ0Z_14),
            .ltout(),
            .carryin(un1_M_this_external_address_q_cry_13),
            .carryout(un1_M_this_external_address_q_cry_14),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam M_this_external_address_q_15_LC_31_24_7.C_ON=1'b0;
    defparam M_this_external_address_q_15_LC_31_24_7.SEQ_MODE=4'b1000;
    defparam M_this_external_address_q_15_LC_31_24_7.LUT_INIT=16'b1011101111101110;
    LogicCell40 M_this_external_address_q_15_LC_31_24_7 (
            .in0(N__25277),
            .in1(N__25048),
            .in2(_gnd_net_),
            .in3(N__25064),
            .lcout(M_this_external_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__25035),
            .ce(),
            .sr(N__24744));
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o4_5_4_LC_32_23_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o4_5_4_LC_32_23_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_0_i_o4_5_4_LC_32_23_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_0_i_o4_5_4_LC_32_23_3  (
            .in0(N__24644),
            .in1(N__24632),
            .in2(N__24620),
            .in3(N__24611),
            .lcout(\this_vga_signals.M_this_state_q_srsts_0_i_o4_5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
