-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     May 9 2022 09:54:28

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : in std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : in std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    debug : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_clk_c : std_logic;
signal \this_vga_signals.N_469_0\ : std_logic;
signal port_rw_c_i : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \N_33\ : std_logic;
signal \N_11\ : std_logic;
signal rgb_c_0 : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1Z0Z_9\ : std_logic;
signal \this_vga_signals.rgb_cnst_i_1Z0Z_3_cascade_\ : std_logic;
signal \this_vga_signals.rgb_cnst_i_1Z0Z_5\ : std_logic;
signal rgb_c_5 : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIAV48E1Z0Z_9\ : std_logic;
signal rgb_c_3 : std_logic;
signal \this_vga_signals.N_379_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIA99QRZ0Z_9_cascade_\ : std_logic;
signal rgb_c_1 : std_logic;
signal \this_vga_signals.rgb_cnst_i_0_5\ : std_logic;
signal \N_11_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \this_vga_signals.if_i3_mux_2_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m2_8_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m8_0_ns_1\ : std_logic;
signal \this_vga_signals.if_m8_0_ns_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_3_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_3\ : std_logic;
signal \this_vga_signals.if_N_4_2\ : std_logic;
signal \this_vga_signals.if_i4_mux_0_1_cascade_\ : std_logic;
signal \this_vga_signals.vsync_1_0_a3_5_cascade_\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \this_vga_signals.if_m13_0_ns_1_cascade_\ : std_logic;
signal \this_vga_signals.if_i3_mux_0_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m13_0_ns_1\ : std_logic;
signal \this_vga_signals.if_i3_mux_0_0_0\ : std_logic;
signal \this_vga_signals.g2_1_cascade_\ : std_logic;
signal \this_vga_signals.g2_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1_1_0\ : std_logic;
signal \this_vga_signals.g0_5_0_1\ : std_logic;
signal \this_vga_signals.g3_0_2_0\ : std_logic;
signal \this_vga_signals.g2_cascade_\ : std_logic;
signal \this_vga_signals.g0_3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_2_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_1_cascade_\ : std_logic;
signal \this_vga_signals.rgb_1_2_cascade_\ : std_logic;
signal \this_vga_signals.if_i3_mux_0_0\ : std_logic;
signal \this_vga_signals.if_i3_mux_2\ : std_logic;
signal \this_vga_signals.g1\ : std_logic;
signal \this_vga_signals.g3_0_2_cascade_\ : std_logic;
signal \this_vga_signals.if_N_3_0_i_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_c_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_1\ : std_logic;
signal \this_vga_signals.if_N_15_mux\ : std_logic;
signal \this_vga_signals.if_m13_ns_1_cascade_\ : std_logic;
signal \this_vga_signals.if_m13_ns\ : std_logic;
signal \this_vga_signals.if_N_7\ : std_logic;
signal \this_vga_signals.d_N_9_0\ : std_logic;
signal \this_vga_signals.rgb_1_4_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIETZ0Z844\ : std_logic;
signal \this_vga_signals.d_N_5_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_i_x1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_2_N_2L1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.un11_address_0_5\ : std_logic;
signal \this_vga_signals.vsync_1_0_a3_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.d_N_8_0\ : std_logic;
signal \this_vga_signals.un11_address_1_5_cascade_\ : std_logic;
signal \this_vga_signals.g0_11_1\ : std_logic;
signal \this_vga_signals.g0_6_0\ : std_logic;
signal \this_vga_signals.g2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g3_cascade_\ : std_logic;
signal \this_vga_signals.g2_4_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_i_1_cascade_\ : std_logic;
signal \this_vga_signals.un11_address_2_5_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_i_x0_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3\ : std_logic;
signal \this_vga_signals.if_N_3_0_i\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_c_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_3_c\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_ac0_1_0\ : std_logic;
signal \this_vga_signals.if_N_3_0_i_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_2\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb2_0\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_0\ : std_logic;
signal \this_vga_signals.g0_5_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_x1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_x0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_1\ : std_logic;
signal \this_vga_signals.un11_address_c4_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_5_4_1_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_5_4_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.un11_address_c4_i\ : std_logic;
signal \this_vga_signals.SUM_2_i_a4_1_0_3_cascade_\ : std_logic;
signal \this_vga_signals.un11_address_c5_a0_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_9_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_8_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_7_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.SUM_2_i_a4_0_a0_2_3_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2_i_a4_a0_2_3\ : std_logic;
signal \this_vga_signals.SUM_2_i_1_0_3\ : std_logic;
signal \this_vga_signals.SUM_2_i_0_1_3\ : std_logic;
signal \this_vga_signals.SUM_2_i_0_3\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\ : std_logic;
signal \N_18\ : std_logic;
signal \this_vga_signals.hsync_1_i_0_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.N_469_0_g\ : std_logic;
signal \this_vga_signals.N_608_g\ : std_logic;
signal \this_vga_signals.N_381_0\ : std_logic;
signal \this_vga_signals.N_390_cascade_\ : std_logic;
signal \this_vga_signals.rgb_cnst_i_0_2_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIO6OD01Z0Z_9_cascade_\ : std_logic;
signal rgb_c_2 : std_logic;
signal \this_vga_signals.g0_i_x2_1_0\ : std_logic;
signal \this_vga_signals.N_10_i\ : std_logic;
signal \this_vga_signals.N_10_i_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x2_5_1\ : std_logic;
signal \this_vga_signals.if_N_13_i_i_1\ : std_logic;
signal \this_vga_signals.g4_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_0_N_3L3\ : std_logic;
signal \this_vga_signals.N_3_1_0_1\ : std_logic;
signal \this_vga_signals.g0_i_x2_1_1_cascade_\ : std_logic;
signal \this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x2_1_1\ : std_logic;
signal \this_vga_signals.g0_i_x1\ : std_logic;
signal \this_vga_signals.g0_i_x0_cascade_\ : std_logic;
signal \this_vga_signals_un16_address_if_i1_mux_0_cascade_\ : std_logic;
signal \this_vga_signals.N_6_i_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_0\ : std_logic;
signal \this_vga_signals.N_11_i\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_axb1\ : std_logic;
signal \this_vga_signals.g0_5_0_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_5_4\ : std_logic;
signal \this_vga_signals.g0_25_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_c\ : std_logic;
signal \this_vga_signals.if_N_13_i_i_1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g2_0_0_0\ : std_logic;
signal \this_vga_signals.N_371_0\ : std_logic;
signal rgb_c_4 : std_logic;
signal \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0\ : std_logic;
signal \this_vga_signals.un11_address_0_7_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2\ : std_logic;
signal \this_vga_signals.g0_3_0\ : std_logic;
signal \this_vga_signals.N_28_0_cascade_\ : std_logic;
signal \this_vga_signals.N_42_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNIVV6F6Z0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.rgb297_i_a3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.SUM_2_i_a4_0_a0_2_3\ : std_logic;
signal \this_vga_signals.N_33_0\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.N_49\ : std_logic;
signal \this_vga_signals.N_33_0_cascade_\ : std_logic;
signal \this_vga_signals.CO0_i_i\ : std_logic;
signal \this_vga_signals.N_45_cascade_\ : std_logic;
signal \N_23_0\ : std_logic;
signal \N_23_0_cascade_\ : std_logic;
signal \this_pixel_clock.M_counter_q_i_1\ : std_logic;
signal \bfn_12_24_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_12_25_0_\ : std_logic;
signal \this_vga_signals.N_22\ : std_logic;
signal \this_vga_signals.g1_0_0_2_cascade_\ : std_logic;
signal \this_vga_signals.N_21\ : std_logic;
signal \this_vga_signals.g0_i_x2_1\ : std_logic;
signal \this_vga_signals.g4_1\ : std_logic;
signal \this_vga_signals.g0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x2_5\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_9_1_0\ : std_logic;
signal \this_vga_signals.g1_5\ : std_logic;
signal \this_vga_signals.N_6\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_0_0_1_cascade_\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.g2_0_1_0\ : std_logic;
signal \this_vga_signals.g0_i_x2_2\ : std_logic;
signal \this_vga_signals.g0_i_0_N_4L5_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_0_N_5L7\ : std_logic;
signal \this_vga_signals.if_i4_mux_0_0_0_1\ : std_logic;
signal \this_vga_signals.N_6_i\ : std_logic;
signal \this_vga_signals.g1_1_2\ : std_logic;
signal \this_vga_signals.g1_4_1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.g0_i_0_N_2L1\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_vcounter_d_1_sqmuxa_i_a3_1\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.if_N_8_i_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_2\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c2_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_9_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb1\ : std_logic;
signal \this_vga_signals.SUM_3_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.N_34\ : std_logic;
signal \this_vga_signals.N_34_cascade_\ : std_logic;
signal \this_vga_signals.SUM_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c2_0\ : std_logic;
signal \this_vga_signals.N_469_1\ : std_logic;
signal debug_0_i : std_logic;
signal \this_vga_signals.rgb_cnst_i_a5_0_0Z0Z_3\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1\ : std_logic;
signal \this_vga_signals.if_m3_5_cascade_\ : std_logic;
signal \this_vga_signals.if_N_3_i\ : std_logic;
signal \this_vga_signals.if_m5_4_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb2_0_1_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_1\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.g0_1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.g4_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_3_d_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_ac0_4\ : std_logic;
signal \this_vga_signals.g0_i_o2_0_0_x2_0_cascade_\ : std_logic;
signal \this_vga_signals.N_16\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_i_1\ : std_logic;
signal \this_vga_signals.if_N_1_i_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0\ : std_logic;
signal \N_401\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_2\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \M_counter_q_RNIJR071_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \M_counter_q_RNIQR4I2_1\ : std_logic;
signal \this_vga_signals.rgb_bmZ0Z_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.if_N_13_i_i_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_0\ : std_logic;
signal \this_vga_signals.if_N_16_i_0\ : std_logic;
signal \this_vga_signals.g0_1_N_5L8\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_0_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_ac0_3_d\ : std_logic;
signal \this_vga_signals.g0_1_N_3L3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.g0_1_N_6L11_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0\ : std_logic;
signal \this_vga_signals.g0_1_N_7L13\ : std_logic;
signal \this_vga_signals.g0_1_N_8L15_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axb2_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.if_N_6_3_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_8\ : std_logic;
signal \N_349_0_cascade_\ : std_logic;
signal port_enb_c : std_logic;
signal \this_delay_clk.M_this_delay_clk_out_0\ : std_logic;
signal debug_0 : std_logic;
signal port_rw_c : std_logic;
signal port_address_c_7 : std_logic;
signal \debug_0_cascade_\ : std_logic;
signal \this_start_data_delay_M_last_q\ : std_logic;
signal \M_current_address_qZ0Z_0\ : std_logic;
signal \N_312_0\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_0\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \un1_M_current_address_q_cry_0\ : std_logic;
signal \un1_M_current_address_q_cry_1\ : std_logic;
signal \un1_M_current_address_q_cry_2\ : std_logic;
signal \un1_M_current_address_q_cry_3\ : std_logic;
signal \un1_M_current_address_q_cry_4\ : std_logic;
signal \un1_M_current_address_q_cry_5\ : std_logic;
signal \un1_M_current_address_q_cry_6\ : std_logic;
signal \un1_M_current_address_q_cry_7\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \un1_M_current_address_q_cry_8\ : std_logic;
signal \un1_M_current_address_q_cry_9\ : std_logic;
signal \un1_M_current_address_q_cry_10\ : std_logic;
signal \un1_M_current_address_q_cry_11\ : std_logic;
signal \un1_M_current_address_q_cry_12\ : std_logic;
signal \this_pixel_clock.M_counter_qZ0Z_0\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \this_vga_signals.rgb_bmZ0Z_0\ : std_logic;
signal \this_vga_signals.rgb_bmZ0Z_2\ : std_logic;
signal \m7_am_cascade_\ : std_logic;
signal m7_ns : std_logic;
signal \m28_cascade_\ : std_logic;
signal \m32_am_cascade_\ : std_logic;
signal m7_bm : std_logic;
signal m32_bm : std_logic;
signal m32_ns : std_logic;
signal rgb_2_4 : std_logic;
signal m29 : std_logic;
signal \this_vga_signals.rgb_bmZ0Z_3\ : std_logic;
signal port_data_c_5 : std_logic;
signal \N_413_cascade_\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_12\ : std_logic;
signal \N_411\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_10\ : std_logic;
signal \M_current_address_qZ0Z_10\ : std_logic;
signal \N_404\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_3\ : std_logic;
signal \M_current_address_qZ0Z_3\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_5\ : std_logic;
signal \N_406\ : std_logic;
signal \M_current_address_qZ0Z_5\ : std_logic;
signal \N_402_cascade_\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_1\ : std_logic;
signal \M_current_address_qZ0Z_1\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_8\ : std_logic;
signal \N_409\ : std_logic;
signal \M_current_address_qZ0Z_8\ : std_logic;
signal \N_412\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_11\ : std_logic;
signal port_data_c_4 : std_logic;
signal \M_current_address_q_RNO_1Z0Z_9\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal rgb291_cry_0 : std_logic;
signal rgb291_cry_1 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal rgb291_cry_2 : std_logic;
signal rgb291 : std_logic;
signal \this_vga_signals.rgb_1_sqmuxa\ : std_logic;
signal \mem_radreg_RNIMTEJ4_0_11\ : std_logic;
signal \mem_radreg_RNIETEJ4_0_11\ : std_logic;
signal \m44_cascade_\ : std_logic;
signal \m22_am_cascade_\ : std_logic;
signal m22_ns : std_logic;
signal m22_bm : std_logic;
signal m24 : std_logic;
signal \m40_cascade_\ : std_logic;
signal m41 : std_logic;
signal m10 : std_logic;
signal \rgb_1_axb_0_cascade_\ : std_logic;
signal m15 : std_logic;
signal rgb_1_0 : std_logic;
signal m37 : std_logic;
signal m19 : std_logic;
signal rgb_1_axb_0 : std_logic;
signal a0_b_0 : std_logic;
signal \m46_am_cascade_\ : std_logic;
signal m46_bm : std_logic;
signal rgb_2_5 : std_logic;
signal \N_352\ : std_logic;
signal \N_408_cascade_\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_7\ : std_logic;
signal \M_current_address_qZ0Z_7\ : std_logic;
signal \N_405\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_4\ : std_logic;
signal \M_current_address_qZ0Z_4\ : std_logic;
signal \M_state_q_ns_0_a3_0_2_0\ : std_logic;
signal \N_351\ : std_logic;
signal \N_403_cascade_\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_2\ : std_logic;
signal \M_current_address_qZ0Z_2\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_13\ : std_logic;
signal \M_state_qZ0Z_1\ : std_logic;
signal \N_407_cascade_\ : std_logic;
signal \M_current_address_q_RNO_1Z0Z_6\ : std_logic;
signal \M_current_address_qZ0Z_6\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal \M_current_address_qZ0Z_9\ : std_logic;
signal \N_410\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_0\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \mem_radreg_RNIETEJ4_11\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal this_vram_mem_radreg_11 : std_logic;
signal \mem_radreg_RNIMTEJ4_11\ : std_logic;
signal m14 : std_logic;
signal \rgb_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \M_vcounter_q_esr_RNIB9J4TN_9\ : std_logic;
signal \M_vcounter_q_esr_RNICJRF0D_9\ : std_logic;
signal rgb_1_cry_0 : std_logic;
signal rgb_1_cry_1 : std_logic;
signal rgb_1_cry_2 : std_logic;
signal rgb_1_6 : std_logic;
signal this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3 : std_logic;
signal \rgb_1_cry_0_0_c_RNOZ0Z_0\ : std_logic;
signal \M_vcounter_q_esr_RNI1H9RHL_9\ : std_logic;
signal rgb_1_3 : std_logic;
signal rgb_1_4 : std_logic;
signal rgb_1_5 : std_logic;
signal \rgb_1_6_THRU_CO\ : std_logic;
signal m36 : std_logic;
signal port_address_c_0 : std_logic;
signal port_address_c_1 : std_logic;
signal \M_state_q_ns_0_a3_0_1_1\ : std_logic;
signal port_data_c_1 : std_logic;
signal \M_this_vram_write_data_1\ : std_logic;
signal \N_349_0\ : std_logic;
signal port_data_c_6 : std_logic;
signal \M_state_qZ0Z_0\ : std_logic;
signal \N_414\ : std_logic;
signal this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1 : std_logic;
signal this_vga_signals_un16_address_if_i1_mux_0 : std_logic;
signal \M_this_vga_signals_address_10\ : std_logic;
signal \rgbZ0Z_1_cascade_\ : std_logic;
signal \M_vcounter_q_esr_RNI2RH6LA_9\ : std_logic;
signal \rgbZ0Z_1\ : std_logic;
signal \M_vcounter_q_esr_RNIVLNKSA_9\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_axbxc3\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal port_data_c_0 : std_logic;
signal \M_this_vram_write_data_0\ : std_logic;
signal \this_vga_signals.SUM_3_1\ : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vram.mem_WE_12\ : std_logic;
signal \this_vga_signals.rgb_1_2\ : std_logic;
signal \this_vram.mem_WE_8\ : std_logic;
signal \this_vram.mem_out_bus0_3\ : std_logic;
signal \this_vram.mem_out_bus4_3\ : std_logic;
signal \this_vram.mem_N_88\ : std_logic;
signal \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\ : std_logic;
signal \this_vram.mem_N_105\ : std_logic;
signal \this_vram.mem_WE_10\ : std_logic;
signal \this_vram.mem_WE_14\ : std_logic;
signal \this_vram_mem_N_112\ : std_logic;
signal \this_vga_signals.rgb_1_4\ : std_logic;
signal clk_0_c_g : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_vram_write_data_3\ : std_logic;
signal \this_vram.mem_out_bus4_1\ : std_logic;
signal \this_vram.mem_out_bus0_1\ : std_logic;
signal \this_vram.mem_out_bus2_1\ : std_logic;
signal \this_vram.mem_out_bus6_1\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_N_91\ : std_logic;
signal \this_vram.mem_out_bus5_1\ : std_logic;
signal \this_vram.mem_out_bus1_1\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus3_1\ : std_logic;
signal \this_vram.mem_out_bus7_1\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus1_0\ : std_logic;
signal \this_vram.mem_out_bus5_0\ : std_logic;
signal \this_vram.mem_out_bus2_3\ : std_logic;
signal \this_vram.mem_out_bus6_3\ : std_logic;
signal \this_vram.mem_mem_2_1_RNI01N11Z0Z_0\ : std_logic;
signal \this_vram.mem_out_bus0_2\ : std_logic;
signal \this_vram.mem_out_bus4_2\ : std_logic;
signal \this_vram.mem_out_bus1_2\ : std_logic;
signal \this_vram.mem_out_bus5_2\ : std_logic;
signal \this_vram.mem_out_bus2_2\ : std_logic;
signal \this_vram.mem_out_bus6_2\ : std_logic;
signal \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_mem_0_1_RNISOIZ0Z11\ : std_logic;
signal \this_vram.mem_N_98\ : std_logic;
signal \this_vram.mem_out_bus1_3\ : std_logic;
signal \this_vram.mem_out_bus5_3\ : std_logic;
signal \this_vram.mem_out_bus3_3\ : std_logic;
signal \this_vram.mem_out_bus7_3\ : std_logic;
signal \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_\ : std_logic;
signal \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0\ : std_logic;
signal \this_vram.mem_N_102\ : std_logic;
signal \this_vram.mem_mem_1_0_RNISSKZ0Z11\ : std_logic;
signal \this_vram_mem_N_109\ : std_logic;
signal \this_vram.mem_out_bus3_2\ : std_logic;
signal \this_vram.mem_out_bus7_2\ : std_logic;
signal \this_vram.mem_mem_1_1_RNIUSKZ0Z11\ : std_logic;
signal \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_\ : std_logic;
signal \this_vram.mem_radregZ0Z_12\ : std_logic;
signal \this_vram.mem_N_95\ : std_logic;
signal \this_vram.mem_out_bus6_0\ : std_logic;
signal \this_vram.mem_out_bus2_0\ : std_logic;
signal \this_vram.mem_mem_2_0_RNIU0NZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus7_0\ : std_logic;
signal \this_vram.mem_out_bus3_0\ : std_logic;
signal \this_vram.mem_mem_3_0_RNI05PZ0Z11\ : std_logic;
signal \this_vram.mem_out_bus0_0\ : std_logic;
signal \this_vram.mem_out_bus4_0\ : std_logic;
signal \this_vram.mem_radregZ0Z_13\ : std_logic;
signal \this_vram.mem_mem_0_0_RNIQOIZ0Z11\ : std_logic;
signal \this_vram.mem_WE_6\ : std_logic;
signal port_data_c_2 : std_logic;
signal \M_this_vram_write_data_2\ : std_logic;
signal \this_vram.mem_WE_4\ : std_logic;
signal \this_vram.mem_WE_0\ : std_logic;
signal \M_current_address_qZ0Z_12\ : std_logic;
signal \M_current_address_qZ0Z_13\ : std_logic;
signal \M_current_address_qZ0Z_11\ : std_logic;
signal \M_this_vram_write_en_0_sqmuxa\ : std_logic;
signal \this_vram.mem_WE_2\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \this_vga_signals.if_m2_5_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0\ : std_logic;
signal \M_this_vga_signals_address_9\ : std_logic;
signal \this_vga_signals.N_9_0\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal port_address_c_5 : std_logic;
signal port_address_c_6 : std_logic;
signal port_address_c_2 : std_logic;
signal port_address_c_3 : std_logic;
signal port_address_c_4 : std_logic;
signal \M_state_q_ns_0_a3_0_0_1_0\ : std_logic;
signal \M_state_q_ns_0_a3_0_0_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic;
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal port_address_wire : std_logic_vector(15 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal port_rw_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    port_address_wire <= port_address;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    port_rw_wire <= port_rw;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \this_vram.mem_out_bus0_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= \N__16019\&\N__20438\&\N__12020\&\N__10076\&\N__17483\&\N__15089\&\N__11852\&\N__17747\&\N__19205\&\N__20123\&\N__10259\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= \N__13640\&\N__15224\&\N__13973\&\N__14816\&\N__15458\&\N__13367\&\N__14675\&\N__13508\&\N__15710\&\N__13241\&\N__12731\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16574\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17582\&'0'&'0'&'0';
    \this_vram.mem_out_bus0_3\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus0_2\ <= \this_vram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_0_1_physical_RADDR_wire\ <= \N__16013\&\N__20432\&\N__12014\&\N__10070\&\N__17477\&\N__15083\&\N__11846\&\N__17741\&\N__19199\&\N__20117\&\N__10253\;
    \this_vram.mem_mem_0_1_physical_WADDR_wire\ <= \N__13634\&\N__15218\&\N__13967\&\N__14810\&\N__15452\&\N__13361\&\N__14669\&\N__13502\&\N__15704\&\N__13235\&\N__12725\;
    \this_vram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18008\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19727\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_1\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_0\ <= \this_vram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_0_physical_RADDR_wire\ <= \N__16007\&\N__20426\&\N__12008\&\N__10064\&\N__17471\&\N__15077\&\N__11840\&\N__17735\&\N__19193\&\N__20111\&\N__10247\;
    \this_vram.mem_mem_1_0_physical_WADDR_wire\ <= \N__13628\&\N__15212\&\N__13961\&\N__14804\&\N__15446\&\N__13355\&\N__14663\&\N__13496\&\N__15698\&\N__13229\&\N__12719\;
    \this_vram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16570\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17577\&'0'&'0'&'0';
    \this_vram.mem_out_bus1_3\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus1_2\ <= \this_vram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_1_1_physical_RADDR_wire\ <= \N__16001\&\N__20420\&\N__12002\&\N__10058\&\N__17465\&\N__15071\&\N__11834\&\N__17729\&\N__19187\&\N__20105\&\N__10241\;
    \this_vram.mem_mem_1_1_physical_WADDR_wire\ <= \N__13622\&\N__15206\&\N__13955\&\N__14798\&\N__15440\&\N__13349\&\N__14657\&\N__13490\&\N__15692\&\N__13223\&\N__12713\;
    \this_vram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18004\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19723\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_1\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_0\ <= \this_vram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_0_physical_RADDR_wire\ <= \N__15995\&\N__20414\&\N__11996\&\N__10052\&\N__17459\&\N__15065\&\N__11828\&\N__17723\&\N__19181\&\N__20099\&\N__10235\;
    \this_vram.mem_mem_2_0_physical_WADDR_wire\ <= \N__13616\&\N__15200\&\N__13949\&\N__14792\&\N__15434\&\N__13343\&\N__14651\&\N__13484\&\N__15686\&\N__13217\&\N__12707\;
    \this_vram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16546\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17565\&'0'&'0'&'0';
    \this_vram.mem_out_bus2_3\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus2_2\ <= \this_vram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_2_1_physical_RADDR_wire\ <= \N__15989\&\N__20408\&\N__11990\&\N__10046\&\N__17453\&\N__15059\&\N__11822\&\N__17717\&\N__19175\&\N__20093\&\N__10229\;
    \this_vram.mem_mem_2_1_physical_WADDR_wire\ <= \N__13610\&\N__15194\&\N__13943\&\N__14786\&\N__15428\&\N__13337\&\N__14645\&\N__13478\&\N__15680\&\N__13211\&\N__12701\;
    \this_vram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17996\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19715\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_1\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_0\ <= \this_vram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_0_physical_RADDR_wire\ <= \N__15983\&\N__20402\&\N__11984\&\N__10040\&\N__17447\&\N__15053\&\N__11816\&\N__17711\&\N__19169\&\N__20087\&\N__10223\;
    \this_vram.mem_mem_3_0_physical_WADDR_wire\ <= \N__13604\&\N__15188\&\N__13937\&\N__14780\&\N__15422\&\N__13331\&\N__14639\&\N__13472\&\N__15674\&\N__13205\&\N__12695\;
    \this_vram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16557\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17581\&'0'&'0'&'0';
    \this_vram.mem_out_bus3_3\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus3_2\ <= \this_vram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_3_1_physical_RADDR_wire\ <= \N__15977\&\N__20396\&\N__11978\&\N__10034\&\N__17441\&\N__15047\&\N__11810\&\N__17705\&\N__19163\&\N__20081\&\N__10217\;
    \this_vram.mem_mem_3_1_physical_WADDR_wire\ <= \N__13598\&\N__15182\&\N__13931\&\N__14774\&\N__15416\&\N__13325\&\N__14633\&\N__13466\&\N__15668\&\N__13199\&\N__12689\;
    \this_vram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17982\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19701\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_1\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_0\ <= \this_vram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_0_physical_RADDR_wire\ <= \N__15971\&\N__20390\&\N__11972\&\N__10028\&\N__17435\&\N__15041\&\N__11804\&\N__17699\&\N__19157\&\N__20075\&\N__10211\;
    \this_vram.mem_mem_4_0_physical_WADDR_wire\ <= \N__13592\&\N__15176\&\N__13925\&\N__14768\&\N__15410\&\N__13319\&\N__14627\&\N__13460\&\N__15662\&\N__13193\&\N__12683\;
    \this_vram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16547\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17573\&'0'&'0'&'0';
    \this_vram.mem_out_bus4_3\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus4_2\ <= \this_vram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_4_1_physical_RADDR_wire\ <= \N__15965\&\N__20384\&\N__11966\&\N__10022\&\N__17429\&\N__15035\&\N__11798\&\N__17693\&\N__19151\&\N__20069\&\N__10205\;
    \this_vram.mem_mem_4_1_physical_WADDR_wire\ <= \N__13586\&\N__15170\&\N__13919\&\N__14762\&\N__15404\&\N__13313\&\N__14621\&\N__13454\&\N__15656\&\N__13187\&\N__12677\;
    \this_vram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17963\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19661\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_1\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_0\ <= \this_vram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_0_physical_RADDR_wire\ <= \N__15959\&\N__20378\&\N__11960\&\N__10016\&\N__17423\&\N__15029\&\N__11792\&\N__17687\&\N__19145\&\N__20063\&\N__10199\;
    \this_vram.mem_mem_5_0_physical_WADDR_wire\ <= \N__13580\&\N__15164\&\N__13913\&\N__14756\&\N__15398\&\N__13307\&\N__14615\&\N__13448\&\N__15650\&\N__13181\&\N__12671\;
    \this_vram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16507\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17519\&'0'&'0'&'0';
    \this_vram.mem_out_bus5_3\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus5_2\ <= \this_vram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_5_1_physical_RADDR_wire\ <= \N__15953\&\N__20372\&\N__11954\&\N__10010\&\N__17417\&\N__15023\&\N__11786\&\N__17681\&\N__19139\&\N__20057\&\N__10193\;
    \this_vram.mem_mem_5_1_physical_WADDR_wire\ <= \N__13574\&\N__15158\&\N__13907\&\N__14750\&\N__15392\&\N__13301\&\N__14609\&\N__13442\&\N__15644\&\N__13175\&\N__12665\;
    \this_vram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17964\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19694\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_1\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_0\ <= \this_vram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_0_physical_RADDR_wire\ <= \N__15947\&\N__20366\&\N__11948\&\N__10004\&\N__17411\&\N__15017\&\N__11780\&\N__17675\&\N__19133\&\N__20051\&\N__10187\;
    \this_vram.mem_mem_6_0_physical_WADDR_wire\ <= \N__13568\&\N__15152\&\N__13901\&\N__14744\&\N__15386\&\N__13295\&\N__14603\&\N__13436\&\N__15638\&\N__13169\&\N__12659\;
    \this_vram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16542\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17555\&'0'&'0'&'0';
    \this_vram.mem_out_bus6_3\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus6_2\ <= \this_vram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_6_1_physical_RADDR_wire\ <= \N__15941\&\N__20360\&\N__11942\&\N__9998\&\N__17405\&\N__15011\&\N__11774\&\N__17669\&\N__19127\&\N__20045\&\N__10181\;
    \this_vram.mem_mem_6_1_physical_WADDR_wire\ <= \N__13562\&\N__15146\&\N__13895\&\N__14738\&\N__15380\&\N__13289\&\N__14597\&\N__13430\&\N__15632\&\N__13163\&\N__12653\;
    \this_vram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__17992\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19711\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_1\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_0\ <= \this_vram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_0_physical_RADDR_wire\ <= \N__15935\&\N__20354\&\N__11936\&\N__9992\&\N__17399\&\N__15005\&\N__11768\&\N__17663\&\N__19121\&\N__20039\&\N__10175\;
    \this_vram.mem_mem_7_0_physical_WADDR_wire\ <= \N__13556\&\N__15140\&\N__13889\&\N__14732\&\N__15374\&\N__13283\&\N__14591\&\N__13424\&\N__15626\&\N__13157\&\N__12647\;
    \this_vram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__16556\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17572\&'0'&'0'&'0';
    \this_vram.mem_out_bus7_3\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_vram.mem_out_bus7_2\ <= \this_vram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_vram.mem_mem_7_1_physical_RADDR_wire\ <= \N__15929\&\N__20348\&\N__11930\&\N__9986\&\N__17393\&\N__14999\&\N__11762\&\N__17657\&\N__19115\&\N__20033\&\N__10169\;
    \this_vram.mem_mem_7_1_physical_WADDR_wire\ <= \N__13550\&\N__15134\&\N__13883\&\N__14726\&\N__15368\&\N__13277\&\N__14585\&\N__13418\&\N__15620\&\N__13151\&\N__12641\;
    \this_vram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18003\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19722\&'0'&'0'&'0';

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18179\,
            RE => \N__14434\,
            WCLKE => \N__18436\,
            WCLK => \N__18180\,
            WE => \N__14418\
        );

    \this_vram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18181\,
            RE => \N__14413\,
            WCLKE => \N__18437\,
            WCLK => \N__18182\,
            WE => \N__14414\
        );

    \this_vram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18183\,
            RE => \N__14412\,
            WCLKE => \N__17375\,
            WCLK => \N__18184\,
            WE => \N__14386\
        );

    \this_vram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18185\,
            RE => \N__14369\,
            WCLKE => \N__17371\,
            WCLK => \N__18186\,
            WE => \N__14385\
        );

    \this_vram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18188\,
            RE => \N__14327\,
            WCLKE => \N__18464\,
            WCLK => \N__18187\,
            WE => \N__14306\
        );

    \this_vram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18190\,
            RE => \N__14311\,
            WCLKE => \N__18460\,
            WCLK => \N__18191\,
            WE => \N__14305\
        );

    \this_vram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18198\,
            RE => \N__14223\,
            WCLKE => \N__17243\,
            WCLK => \N__18199\,
            WE => \N__14172\
        );

    \this_vram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18206\,
            RE => \N__14307\,
            WCLKE => \N__17242\,
            WCLK => \N__18207\,
            WE => \N__14278\
        );

    \this_vram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18210\,
            RE => \N__14368\,
            WCLKE => \N__19789\,
            WCLK => \N__18211\,
            WE => \N__14338\
        );

    \this_vram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18218\,
            RE => \N__14351\,
            WCLKE => \N__19793\,
            WCLK => \N__18219\,
            WE => \N__14339\
        );

    \this_vram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18224\,
            RE => \N__14398\,
            WCLKE => \N__19642\,
            WCLK => \N__18225\,
            WE => \N__14388\
        );

    \this_vram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18228\,
            RE => \N__14399\,
            WCLKE => \N__19643\,
            WCLK => \N__18229\,
            WE => \N__14389\
        );

    \this_vram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18232\,
            RE => \N__14426\,
            WCLKE => \N__19222\,
            WCLK => \N__18233\,
            WE => \N__14271\
        );

    \this_vram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18234\,
            RE => \N__14430\,
            WCLKE => \N__19226\,
            WCLK => \N__18235\,
            WE => \N__14419\
        );

    \this_vram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18236\,
            RE => \N__14440\,
            WCLKE => \N__19621\,
            WCLK => \N__18237\,
            WE => \N__14435\
        );

    \this_vram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18238\,
            RE => \N__14441\,
            WCLKE => \N__19625\,
            WCLK => \N__18239\,
            WE => \N__14436\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__20796\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20798\,
            DIN => \N__20797\,
            DOUT => \N__20796\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20798\,
            PADOUT => \N__20797\,
            PADIN => \N__20796\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20787\,
            DIN => \N__20786\,
            DOUT => \N__20785\,
            PACKAGEPIN => debug_wire
        );

    \debug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20787\,
            PADOUT => \N__20786\,
            PADIN => \N__20785\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__10457\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20778\,
            DIN => \N__20777\,
            DOUT => \N__20776\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20778\,
            PADOUT => \N__20777\,
            PADIN => \N__20776\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7100\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20769\,
            DIN => \N__20768\,
            DOUT => \N__20767\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20769\,
            PADOUT => \N__20768\,
            PADIN => \N__20767\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8726\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20760\,
            DIN => \N__20759\,
            DOUT => \N__20758\,
            PACKAGEPIN => port_address_wire(0)
        );

    \port_address_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20760\,
            PADOUT => \N__20759\,
            PADIN => \N__20758\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20751\,
            DIN => \N__20750\,
            DOUT => \N__20749\,
            PACKAGEPIN => port_address_wire(1)
        );

    \port_address_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20751\,
            PADOUT => \N__20750\,
            PADIN => \N__20749\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20742\,
            DIN => \N__20741\,
            DOUT => \N__20740\,
            PACKAGEPIN => port_address_wire(2)
        );

    \port_address_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20742\,
            PADOUT => \N__20741\,
            PADIN => \N__20740\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20733\,
            DIN => \N__20732\,
            DOUT => \N__20731\,
            PACKAGEPIN => port_address_wire(3)
        );

    \port_address_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20733\,
            PADOUT => \N__20732\,
            PADIN => \N__20731\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20724\,
            DIN => \N__20723\,
            DOUT => \N__20722\,
            PACKAGEPIN => port_address_wire(4)
        );

    \port_address_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20724\,
            PADOUT => \N__20723\,
            PADIN => \N__20722\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20715\,
            DIN => \N__20714\,
            DOUT => \N__20713\,
            PACKAGEPIN => port_address_wire(5)
        );

    \port_address_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20715\,
            PADOUT => \N__20714\,
            PADIN => \N__20713\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20706\,
            DIN => \N__20705\,
            DOUT => \N__20704\,
            PACKAGEPIN => port_address_wire(6)
        );

    \port_address_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20706\,
            PADOUT => \N__20705\,
            PADIN => \N__20704\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20697\,
            DIN => \N__20696\,
            DOUT => \N__20695\,
            PACKAGEPIN => port_address_wire(7)
        );

    \port_address_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20697\,
            PADOUT => \N__20696\,
            PADIN => \N__20695\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20688\,
            DIN => \N__20687\,
            DOUT => \N__20686\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20688\,
            PADOUT => \N__20687\,
            PADIN => \N__20686\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20679\,
            DIN => \N__20678\,
            DOUT => \N__20677\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20679\,
            PADOUT => \N__20678\,
            PADIN => \N__20677\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20670\,
            DIN => \N__20669\,
            DOUT => \N__20668\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20670\,
            PADOUT => \N__20669\,
            PADIN => \N__20668\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20661\,
            DIN => \N__20660\,
            DOUT => \N__20659\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20661\,
            PADOUT => \N__20660\,
            PADIN => \N__20659\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20652\,
            DIN => \N__20651\,
            DOUT => \N__20650\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20652\,
            PADOUT => \N__20651\,
            PADIN => \N__20650\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20643\,
            DIN => \N__20642\,
            DOUT => \N__20641\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20643\,
            PADOUT => \N__20642\,
            PADIN => \N__20641\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20634\,
            DIN => \N__20633\,
            DOUT => \N__20632\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20634\,
            PADOUT => \N__20633\,
            PADIN => \N__20632\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20625\,
            DIN => \N__20624\,
            DOUT => \N__20623\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20625\,
            PADOUT => \N__20624\,
            PADIN => \N__20623\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20616\,
            DIN => \N__20615\,
            DOUT => \N__20614\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20616\,
            PADOUT => \N__20615\,
            PADIN => \N__20614\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7034\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20607\,
            DIN => \N__20606\,
            DOUT => \N__20605\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20607\,
            PADOUT => \N__20606\,
            PADIN => \N__20605\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__14387\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20598\,
            DIN => \N__20597\,
            DOUT => \N__20596\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20598\,
            PADOUT => \N__20597\,
            PADIN => \N__20596\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20589\,
            DIN => \N__20588\,
            DOUT => \N__20587\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20589\,
            PADOUT => \N__20588\,
            PADIN => \N__20587\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7160\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20580\,
            DIN => \N__20579\,
            DOUT => \N__20578\,
            PACKAGEPIN => port_rw_wire
        );

    \port_rw_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20580\,
            PADOUT => \N__20579\,
            PADIN => \N__20578\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20571\,
            DIN => \N__20570\,
            DOUT => \N__20569\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20571\,
            PADOUT => \N__20570\,
            PADIN => \N__20569\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7082\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20562\,
            DIN => \N__20561\,
            DOUT => \N__20560\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20562\,
            PADOUT => \N__20561\,
            PADIN => \N__20560\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7178\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20553\,
            DIN => \N__20552\,
            DOUT => \N__20551\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20553\,
            PADOUT => \N__20552\,
            PADIN => \N__20551\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8828\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20544\,
            DIN => \N__20543\,
            DOUT => \N__20542\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20544\,
            PADOUT => \N__20543\,
            PADIN => \N__20542\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7211\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20535\,
            DIN => \N__20534\,
            DOUT => \N__20533\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20535\,
            PADOUT => \N__20534\,
            PADIN => \N__20533\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__9032\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20526\,
            DIN => \N__20525\,
            DOUT => \N__20524\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20526\,
            PADOUT => \N__20525\,
            PADIN => \N__20524\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7238\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20517\,
            DIN => \N__20516\,
            DOUT => \N__20515\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__20517\,
            PADOUT => \N__20516\,
            PADIN => \N__20515\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20508\,
            DIN => \N__20507\,
            DOUT => \N__20506\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20508\,
            PADOUT => \N__20507\,
            PADIN => \N__20506\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7091\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20499\,
            DIN => \N__20498\,
            DOUT => \N__20497\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__20499\,
            PADOUT => \N__20498\,
            PADIN => \N__20497\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__7343\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__4987\ : InMux
    port map (
            O => \N__20480\,
            I => \N__20477\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__20477\,
            I => \N__20474\
        );

    \I__4985\ : Span12Mux_s10_h
    port map (
            O => \N__20474\,
            I => \N__20470\
        );

    \I__4984\ : InMux
    port map (
            O => \N__20473\,
            I => \N__20467\
        );

    \I__4983\ : Span12Mux_v
    port map (
            O => \N__20470\,
            I => \N__20464\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__20467\,
            I => \this_vga_signals.if_m2_5_0\
        );

    \I__4981\ : Odrv12
    port map (
            O => \N__20464\,
            I => \this_vga_signals.if_m2_5_0\
        );

    \I__4980\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20456\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__20456\,
            I => \N__20453\
        );

    \I__4978\ : Span12Mux_h
    port map (
            O => \N__20453\,
            I => \N__20450\
        );

    \I__4977\ : Span12Mux_v
    port map (
            O => \N__20450\,
            I => \N__20446\
        );

    \I__4976\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20443\
        );

    \I__4975\ : Odrv12
    port map (
            O => \N__20446\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__20443\,
            I => \this_vga_signals.mult1_un68_sum_c3_0\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__4972\ : CascadeBuf
    port map (
            O => \N__20435\,
            I => \N__20432\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__20432\,
            I => \N__20429\
        );

    \I__4970\ : CascadeBuf
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__4969\ : CascadeMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__4968\ : CascadeBuf
    port map (
            O => \N__20423\,
            I => \N__20420\
        );

    \I__4967\ : CascadeMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__4966\ : CascadeBuf
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__4964\ : CascadeBuf
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__4962\ : CascadeBuf
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__4961\ : CascadeMux
    port map (
            O => \N__20402\,
            I => \N__20399\
        );

    \I__4960\ : CascadeBuf
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__4959\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__4958\ : CascadeBuf
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__4956\ : CascadeBuf
    port map (
            O => \N__20387\,
            I => \N__20384\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__4954\ : CascadeBuf
    port map (
            O => \N__20381\,
            I => \N__20378\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__4952\ : CascadeBuf
    port map (
            O => \N__20375\,
            I => \N__20372\
        );

    \I__4951\ : CascadeMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__4950\ : CascadeBuf
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__4949\ : CascadeMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__4948\ : CascadeBuf
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__4946\ : CascadeBuf
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__4944\ : CascadeBuf
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__4942\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20342\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__20342\,
            I => \M_this_vga_signals_address_9\
        );

    \I__4940\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20335\
        );

    \I__4939\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20326\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20320\
        );

    \I__4937\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20317\
        );

    \I__4936\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20314\
        );

    \I__4935\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20311\
        );

    \I__4934\ : InMux
    port map (
            O => \N__20331\,
            I => \N__20305\
        );

    \I__4933\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20302\
        );

    \I__4932\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20299\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__20326\,
            I => \N__20295\
        );

    \I__4930\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20292\
        );

    \I__4929\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20286\
        );

    \I__4928\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20283\
        );

    \I__4927\ : Sp12to4
    port map (
            O => \N__20320\,
            I => \N__20280\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20273\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__20314\,
            I => \N__20273\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__20311\,
            I => \N__20273\
        );

    \I__4923\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20270\
        );

    \I__4922\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20267\
        );

    \I__4921\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20263\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__20305\,
            I => \N__20257\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__20302\,
            I => \N__20257\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20254\
        );

    \I__4917\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20251\
        );

    \I__4916\ : Span4Mux_v
    port map (
            O => \N__20295\,
            I => \N__20246\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20246\
        );

    \I__4914\ : InMux
    port map (
            O => \N__20291\,
            I => \N__20243\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__20290\,
            I => \N__20240\
        );

    \I__4912\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20237\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__20286\,
            I => \N__20232\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__20283\,
            I => \N__20232\
        );

    \I__4909\ : Span12Mux_v
    port map (
            O => \N__20280\,
            I => \N__20225\
        );

    \I__4908\ : Span12Mux_s7_v
    port map (
            O => \N__20273\,
            I => \N__20225\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20225\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__20267\,
            I => \N__20222\
        );

    \I__4905\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20219\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__20263\,
            I => \N__20216\
        );

    \I__4903\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20213\
        );

    \I__4902\ : Span4Mux_h
    port map (
            O => \N__20257\,
            I => \N__20210\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__20254\,
            I => \N__20201\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__20251\,
            I => \N__20201\
        );

    \I__4899\ : Span4Mux_h
    port map (
            O => \N__20246\,
            I => \N__20201\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20201\
        );

    \I__4897\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20198\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20191\
        );

    \I__4895\ : Sp12to4
    port map (
            O => \N__20232\,
            I => \N__20191\
        );

    \I__4894\ : Span12Mux_h
    port map (
            O => \N__20225\,
            I => \N__20191\
        );

    \I__4893\ : Span12Mux_v
    port map (
            O => \N__20222\,
            I => \N__20182\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__20219\,
            I => \N__20182\
        );

    \I__4891\ : Span12Mux_h
    port map (
            O => \N__20216\,
            I => \N__20182\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__20213\,
            I => \N__20182\
        );

    \I__4889\ : Span4Mux_h
    port map (
            O => \N__20210\,
            I => \N__20177\
        );

    \I__4888\ : Span4Mux_h
    port map (
            O => \N__20201\,
            I => \N__20177\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__20198\,
            I => \this_vga_signals.N_9_0\
        );

    \I__4886\ : Odrv12
    port map (
            O => \N__20191\,
            I => \this_vga_signals.N_9_0\
        );

    \I__4885\ : Odrv12
    port map (
            O => \N__20182\,
            I => \this_vga_signals.N_9_0\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__20177\,
            I => \this_vga_signals.N_9_0\
        );

    \I__4883\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20164\
        );

    \I__4882\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20161\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20158\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__20161\,
            I => \N__20155\
        );

    \I__4879\ : Sp12to4
    port map (
            O => \N__20158\,
            I => \N__20150\
        );

    \I__4878\ : Sp12to4
    port map (
            O => \N__20155\,
            I => \N__20150\
        );

    \I__4877\ : Span12Mux_s9_v
    port map (
            O => \N__20150\,
            I => \N__20145\
        );

    \I__4876\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20140\
        );

    \I__4875\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20140\
        );

    \I__4874\ : Odrv12
    port map (
            O => \N__20145\,
            I => \this_vga_signals.mult1_un75_sum_c3_0\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__20140\,
            I => \this_vga_signals.mult1_un75_sum_c3_0\
        );

    \I__4872\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__4870\ : Span12Mux_h
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__4869\ : Odrv12
    port map (
            O => \N__20126\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__20123\,
            I => \N__20120\
        );

    \I__4867\ : CascadeBuf
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__4865\ : CascadeBuf
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__4864\ : CascadeMux
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__4863\ : CascadeBuf
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__4861\ : CascadeBuf
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__4859\ : CascadeBuf
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__4857\ : CascadeBuf
    port map (
            O => \N__20090\,
            I => \N__20087\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__4855\ : CascadeBuf
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__4853\ : CascadeBuf
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__4851\ : CascadeBuf
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__4850\ : CascadeMux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__4849\ : CascadeBuf
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__4847\ : CascadeBuf
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__4846\ : CascadeMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__4845\ : CascadeBuf
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__4843\ : CascadeBuf
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__4842\ : CascadeMux
    port map (
            O => \N__20045\,
            I => \N__20042\
        );

    \I__4841\ : CascadeBuf
    port map (
            O => \N__20042\,
            I => \N__20039\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__20039\,
            I => \N__20036\
        );

    \I__4839\ : CascadeBuf
    port map (
            O => \N__20036\,
            I => \N__20033\
        );

    \I__4838\ : CascadeMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__4837\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__20027\,
            I => \M_this_vga_signals_address_1\
        );

    \I__4835\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__20021\,
            I => port_address_c_5
        );

    \I__4833\ : InMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__4831\ : Span4Mux_v
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__20009\,
            I => port_address_c_6
        );

    \I__4829\ : InMux
    port map (
            O => \N__20006\,
            I => \N__20003\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__4827\ : Span12Mux_s10_h
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__4826\ : Odrv12
    port map (
            O => \N__19997\,
            I => port_address_c_2
        );

    \I__4825\ : InMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__4823\ : Span12Mux_v
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__19985\,
            I => port_address_c_3
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__4820\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__19976\,
            I => port_address_c_4
        );

    \I__4818\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__19967\,
            I => \M_state_q_ns_0_a3_0_0_1_0\
        );

    \I__4815\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19960\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__19963\,
            I => \N__19957\
        );

    \I__4813\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19954\
        );

    \I__4812\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19951\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__19954\,
            I => \N__19946\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__19951\,
            I => \N__19946\
        );

    \I__4809\ : Span12Mux_h
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__4808\ : Span12Mux_h
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__4807\ : Odrv12
    port map (
            O => \N__19940\,
            I => \M_state_q_ns_0_a3_0_0_0\
        );

    \I__4806\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__19934\,
            I => \this_vram.mem_mem_2_0_RNIU0NZ0Z11\
        );

    \I__4804\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__4802\ : Sp12to4
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__4801\ : Span12Mux_v
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__4800\ : Odrv12
    port map (
            O => \N__19919\,
            I => \this_vram.mem_out_bus7_0\
        );

    \I__4799\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__19910\,
            I => \this_vram.mem_out_bus3_0\
        );

    \I__4796\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__19904\,
            I => \this_vram.mem_mem_3_0_RNI05PZ0Z11\
        );

    \I__4794\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__4792\ : Sp12to4
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__4791\ : Span12Mux_v
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__4790\ : Odrv12
    port map (
            O => \N__19889\,
            I => \this_vram.mem_out_bus0_0\
        );

    \I__4789\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__19883\,
            I => \this_vram.mem_out_bus4_0\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__19880\,
            I => \N__19873\
        );

    \I__4786\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19863\
        );

    \I__4785\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19863\
        );

    \I__4784\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19854\
        );

    \I__4783\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19854\
        );

    \I__4782\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19854\
        );

    \I__4781\ : InMux
    port map (
            O => \N__19872\,
            I => \N__19854\
        );

    \I__4780\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19851\
        );

    \I__4779\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19844\
        );

    \I__4778\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19844\
        );

    \I__4777\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19844\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__19863\,
            I => \N__19834\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19834\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19834\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__19844\,
            I => \N__19831\
        );

    \I__4772\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19824\
        );

    \I__4771\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19824\
        );

    \I__4770\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19824\
        );

    \I__4769\ : Span4Mux_v
    port map (
            O => \N__19834\,
            I => \N__19814\
        );

    \I__4768\ : Span4Mux_h
    port map (
            O => \N__19831\,
            I => \N__19814\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__19824\,
            I => \N__19814\
        );

    \I__4766\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19809\
        );

    \I__4765\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19809\
        );

    \I__4764\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19806\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__19814\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__19809\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__19806\,
            I => \this_vram.mem_radregZ0Z_13\
        );

    \I__4760\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__19796\,
            I => \this_vram.mem_mem_0_0_RNIQOIZ0Z11\
        );

    \I__4758\ : CEMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19786\
        );

    \I__4756\ : CEMux
    port map (
            O => \N__19789\,
            I => \N__19783\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__19786\,
            I => \N__19780\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__19783\,
            I => \N__19777\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__19780\,
            I => \this_vram.mem_WE_6\
        );

    \I__4752\ : Odrv4
    port map (
            O => \N__19777\,
            I => \this_vram.mem_WE_6\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__19772\,
            I => \N__19768\
        );

    \I__4750\ : InMux
    port map (
            O => \N__19771\,
            I => \N__19764\
        );

    \I__4749\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19761\
        );

    \I__4748\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19758\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__19764\,
            I => \N__19753\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__19761\,
            I => \N__19753\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__19758\,
            I => \N__19750\
        );

    \I__4744\ : Span4Mux_v
    port map (
            O => \N__19753\,
            I => \N__19747\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__19750\,
            I => \N__19744\
        );

    \I__4742\ : Sp12to4
    port map (
            O => \N__19747\,
            I => \N__19741\
        );

    \I__4741\ : Sp12to4
    port map (
            O => \N__19744\,
            I => \N__19738\
        );

    \I__4740\ : Span12Mux_h
    port map (
            O => \N__19741\,
            I => \N__19735\
        );

    \I__4739\ : Span12Mux_h
    port map (
            O => \N__19738\,
            I => \N__19732\
        );

    \I__4738\ : Odrv12
    port map (
            O => \N__19735\,
            I => port_data_c_2
        );

    \I__4737\ : Odrv12
    port map (
            O => \N__19732\,
            I => port_data_c_2
        );

    \I__4736\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19719\
        );

    \I__4734\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19716\
        );

    \I__4733\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19712\
        );

    \I__4732\ : Span4Mux_h
    port map (
            O => \N__19719\,
            I => \N__19708\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__19716\,
            I => \N__19705\
        );

    \I__4730\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19702\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19698\
        );

    \I__4728\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19695\
        );

    \I__4727\ : Span4Mux_v
    port map (
            O => \N__19708\,
            I => \N__19689\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__19705\,
            I => \N__19689\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__19702\,
            I => \N__19686\
        );

    \I__4724\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19683\
        );

    \I__4723\ : Span4Mux_v
    port map (
            O => \N__19698\,
            I => \N__19678\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__19695\,
            I => \N__19678\
        );

    \I__4721\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19675\
        );

    \I__4720\ : Span4Mux_v
    port map (
            O => \N__19689\,
            I => \N__19670\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__19686\,
            I => \N__19670\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__19683\,
            I => \N__19667\
        );

    \I__4717\ : Span4Mux_v
    port map (
            O => \N__19678\,
            I => \N__19662\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__19675\,
            I => \N__19662\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__19670\,
            I => \N__19656\
        );

    \I__4714\ : Span4Mux_h
    port map (
            O => \N__19667\,
            I => \N__19656\
        );

    \I__4713\ : Span4Mux_v
    port map (
            O => \N__19662\,
            I => \N__19653\
        );

    \I__4712\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19650\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__19656\,
            I => \M_this_vram_write_data_2\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__19653\,
            I => \M_this_vram_write_data_2\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__19650\,
            I => \M_this_vram_write_data_2\
        );

    \I__4708\ : CEMux
    port map (
            O => \N__19643\,
            I => \N__19639\
        );

    \I__4707\ : CEMux
    port map (
            O => \N__19642\,
            I => \N__19636\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__19639\,
            I => \N__19631\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__19636\,
            I => \N__19631\
        );

    \I__4704\ : Span4Mux_v
    port map (
            O => \N__19631\,
            I => \N__19628\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__19628\,
            I => \this_vram.mem_WE_4\
        );

    \I__4702\ : CEMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__19622\,
            I => \N__19618\
        );

    \I__4700\ : CEMux
    port map (
            O => \N__19621\,
            I => \N__19615\
        );

    \I__4699\ : Span4Mux_s2_v
    port map (
            O => \N__19618\,
            I => \N__19610\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__19615\,
            I => \N__19610\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__19604\,
            I => \this_vram.mem_WE_0\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__4693\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19592\
        );

    \I__4692\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19589\
        );

    \I__4691\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19586\
        );

    \I__4690\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19583\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__19592\,
            I => \N__19576\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__19589\,
            I => \N__19571\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__19586\,
            I => \N__19571\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__19583\,
            I => \N__19568\
        );

    \I__4685\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19563\
        );

    \I__4684\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19563\
        );

    \I__4683\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19560\
        );

    \I__4682\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19557\
        );

    \I__4681\ : Span4Mux_v
    port map (
            O => \N__19576\,
            I => \N__19552\
        );

    \I__4680\ : Span4Mux_v
    port map (
            O => \N__19571\,
            I => \N__19552\
        );

    \I__4679\ : Span4Mux_v
    port map (
            O => \N__19568\,
            I => \N__19549\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__19563\,
            I => \N__19546\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__19560\,
            I => \N__19541\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__19557\,
            I => \N__19538\
        );

    \I__4675\ : Span4Mux_h
    port map (
            O => \N__19552\,
            I => \N__19535\
        );

    \I__4674\ : Span4Mux_v
    port map (
            O => \N__19549\,
            I => \N__19530\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__19546\,
            I => \N__19530\
        );

    \I__4672\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19527\
        );

    \I__4671\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19524\
        );

    \I__4670\ : Span12Mux_s10_h
    port map (
            O => \N__19541\,
            I => \N__19519\
        );

    \I__4669\ : Span12Mux_v
    port map (
            O => \N__19538\,
            I => \N__19519\
        );

    \I__4668\ : Span4Mux_h
    port map (
            O => \N__19535\,
            I => \N__19516\
        );

    \I__4667\ : Span4Mux_h
    port map (
            O => \N__19530\,
            I => \N__19513\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__19527\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__19524\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4664\ : Odrv12
    port map (
            O => \N__19519\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__19516\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__19513\,
            I => \M_current_address_qZ0Z_12\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__19502\,
            I => \N__19493\
        );

    \I__4660\ : CascadeMux
    port map (
            O => \N__19501\,
            I => \N__19490\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__19500\,
            I => \N__19487\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__19499\,
            I => \N__19484\
        );

    \I__4657\ : CascadeMux
    port map (
            O => \N__19498\,
            I => \N__19481\
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__19497\,
            I => \N__19477\
        );

    \I__4655\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19472\
        );

    \I__4654\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19472\
        );

    \I__4653\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19469\
        );

    \I__4652\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19466\
        );

    \I__4651\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19463\
        );

    \I__4650\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19459\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19454\
        );

    \I__4648\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19454\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__19472\,
            I => \N__19451\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19448\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__19466\,
            I => \N__19443\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__19463\,
            I => \N__19443\
        );

    \I__4643\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19440\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__19459\,
            I => \N__19433\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__19454\,
            I => \N__19433\
        );

    \I__4640\ : Span4Mux_v
    port map (
            O => \N__19451\,
            I => \N__19433\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__19448\,
            I => \N__19427\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__19443\,
            I => \N__19427\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__19440\,
            I => \N__19424\
        );

    \I__4636\ : Span4Mux_v
    port map (
            O => \N__19433\,
            I => \N__19421\
        );

    \I__4635\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19418\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__19427\,
            I => \N__19415\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__19424\,
            I => \N__19410\
        );

    \I__4632\ : Span4Mux_h
    port map (
            O => \N__19421\,
            I => \N__19410\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__19418\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__19415\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__19410\,
            I => \M_current_address_qZ0Z_13\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19398\
        );

    \I__4627\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19395\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__19401\,
            I => \N__19387\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__19398\,
            I => \N__19383\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__19395\,
            I => \N__19379\
        );

    \I__4623\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19376\
        );

    \I__4622\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19373\
        );

    \I__4621\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19370\
        );

    \I__4620\ : InMux
    port map (
            O => \N__19391\,
            I => \N__19367\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19364\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19359\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19386\,
            I => \N__19359\
        );

    \I__4616\ : Span4Mux_h
    port map (
            O => \N__19383\,
            I => \N__19356\
        );

    \I__4615\ : InMux
    port map (
            O => \N__19382\,
            I => \N__19353\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__19379\,
            I => \N__19350\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19341\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__19373\,
            I => \N__19341\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__19370\,
            I => \N__19341\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__19367\,
            I => \N__19341\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__19364\,
            I => \N__19336\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__19359\,
            I => \N__19336\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__19356\,
            I => \N__19333\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__19353\,
            I => \N__19328\
        );

    \I__4605\ : Span4Mux_h
    port map (
            O => \N__19350\,
            I => \N__19328\
        );

    \I__4604\ : Span12Mux_h
    port map (
            O => \N__19341\,
            I => \N__19325\
        );

    \I__4603\ : Odrv12
    port map (
            O => \N__19336\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__19333\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4601\ : Odrv4
    port map (
            O => \N__19328\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4600\ : Odrv12
    port map (
            O => \N__19325\,
            I => \M_current_address_qZ0Z_11\
        );

    \I__4599\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19306\
        );

    \I__4598\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19301\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19301\
        );

    \I__4596\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19298\
        );

    \I__4595\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19292\
        );

    \I__4594\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19292\
        );

    \I__4593\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19289\
        );

    \I__4592\ : InMux
    port map (
            O => \N__19309\,
            I => \N__19286\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__19306\,
            I => \N__19283\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19278\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__19298\,
            I => \N__19278\
        );

    \I__4588\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19273\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19266\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19266\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19266\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__19283\,
            I => \N__19261\
        );

    \I__4583\ : Span4Mux_v
    port map (
            O => \N__19278\,
            I => \N__19261\
        );

    \I__4582\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19258\
        );

    \I__4581\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19255\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__19273\,
            I => \N__19252\
        );

    \I__4579\ : Span12Mux_h
    port map (
            O => \N__19266\,
            I => \N__19248\
        );

    \I__4578\ : Sp12to4
    port map (
            O => \N__19261\,
            I => \N__19241\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__19258\,
            I => \N__19241\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__19255\,
            I => \N__19241\
        );

    \I__4575\ : Span4Mux_h
    port map (
            O => \N__19252\,
            I => \N__19238\
        );

    \I__4574\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19235\
        );

    \I__4573\ : Odrv12
    port map (
            O => \N__19248\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4572\ : Odrv12
    port map (
            O => \N__19241\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__19238\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__19235\,
            I => \M_this_vram_write_en_0_sqmuxa\
        );

    \I__4569\ : CEMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__19223\,
            I => \N__19219\
        );

    \I__4567\ : CEMux
    port map (
            O => \N__19222\,
            I => \N__19216\
        );

    \I__4566\ : Span4Mux_v
    port map (
            O => \N__19219\,
            I => \N__19211\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__19216\,
            I => \N__19211\
        );

    \I__4564\ : Span4Mux_v
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__4563\ : Odrv4
    port map (
            O => \N__19208\,
            I => \this_vram.mem_WE_2\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__4561\ : CascadeBuf
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__4559\ : CascadeBuf
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__4557\ : CascadeBuf
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__4555\ : CascadeBuf
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__4553\ : CascadeBuf
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__19175\,
            I => \N__19172\
        );

    \I__4551\ : CascadeBuf
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__4550\ : CascadeMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__4549\ : CascadeBuf
    port map (
            O => \N__19166\,
            I => \N__19163\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__4547\ : CascadeBuf
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__4545\ : CascadeBuf
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__4543\ : CascadeBuf
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__4541\ : CascadeBuf
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__4539\ : CascadeBuf
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__4538\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__4537\ : CascadeBuf
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__4535\ : CascadeBuf
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__4533\ : CascadeBuf
    port map (
            O => \N__19118\,
            I => \N__19115\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__4531\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__19106\,
            I => \M_this_vga_signals_address_2\
        );

    \I__4528\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__19097\,
            I => \this_vram.mem_out_bus2_2\
        );

    \I__4525\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__4523\ : Span4Mux_h
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__4522\ : Sp12to4
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__4521\ : Span12Mux_v
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__4520\ : Odrv12
    port map (
            O => \N__19079\,
            I => \this_vram.mem_out_bus6_2\
        );

    \I__4519\ : CascadeMux
    port map (
            O => \N__19076\,
            I => \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__19070\,
            I => \this_vram.mem_mem_0_1_RNISOIZ0Z11\
        );

    \I__4516\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19063\
        );

    \I__4515\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19060\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__19063\,
            I => \N__19055\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__19060\,
            I => \N__19055\
        );

    \I__4512\ : Span4Mux_v
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__19049\,
            I => \this_vram.mem_N_98\
        );

    \I__4509\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__4507\ : Sp12to4
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__4506\ : Span12Mux_v
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__4505\ : Odrv12
    port map (
            O => \N__19034\,
            I => \this_vram.mem_out_bus1_3\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__19028\,
            I => \N__19025\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__4501\ : Span4Mux_v
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__19019\,
            I => \this_vram.mem_out_bus5_3\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__19016\,
            I => \N__19013\
        );

    \I__4498\ : InMux
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__19010\,
            I => \this_vram.mem_out_bus3_3\
        );

    \I__4496\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__4494\ : Span4Mux_v
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__4493\ : Span4Mux_v
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__4492\ : Span4Mux_v
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__4491\ : Span4Mux_v
    port map (
            O => \N__18992\,
            I => \N__18989\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__18989\,
            I => \this_vram.mem_out_bus7_3\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__18986\,
            I => \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_\
        );

    \I__4488\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18980\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__18977\,
            I => \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0\
        );

    \I__4485\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18970\
        );

    \I__4484\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18967\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__18970\,
            I => \N__18962\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__18967\,
            I => \N__18962\
        );

    \I__4481\ : Span4Mux_v
    port map (
            O => \N__18962\,
            I => \N__18959\
        );

    \I__4480\ : Span4Mux_h
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__18956\,
            I => \this_vram.mem_N_102\
        );

    \I__4478\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__4476\ : Odrv4
    port map (
            O => \N__18947\,
            I => \this_vram.mem_mem_1_0_RNISSKZ0Z11\
        );

    \I__4475\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18940\
        );

    \I__4474\ : InMux
    port map (
            O => \N__18943\,
            I => \N__18937\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__18940\,
            I => \N__18931\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__18937\,
            I => \N__18931\
        );

    \I__4471\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18928\
        );

    \I__4470\ : Span4Mux_v
    port map (
            O => \N__18931\,
            I => \N__18925\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__4468\ : Span4Mux_h
    port map (
            O => \N__18925\,
            I => \N__18917\
        );

    \I__4467\ : Span4Mux_v
    port map (
            O => \N__18922\,
            I => \N__18917\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__18914\,
            I => \this_vram_mem_N_109\
        );

    \I__4464\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__18908\,
            I => \this_vram.mem_out_bus3_2\
        );

    \I__4462\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__4460\ : Span4Mux_v
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__4459\ : Sp12to4
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4458\ : Span12Mux_v
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__4457\ : Odrv12
    port map (
            O => \N__18890\,
            I => \this_vram.mem_out_bus7_2\
        );

    \I__4456\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__18884\,
            I => \this_vram.mem_mem_1_1_RNIUSKZ0Z11\
        );

    \I__4454\ : CascadeMux
    port map (
            O => \N__18881\,
            I => \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_\
        );

    \I__4453\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18873\
        );

    \I__4452\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18870\
        );

    \I__4451\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18867\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__18873\,
            I => \N__18858\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__18870\,
            I => \N__18858\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__18867\,
            I => \N__18855\
        );

    \I__4447\ : InMux
    port map (
            O => \N__18866\,
            I => \N__18852\
        );

    \I__4446\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18844\
        );

    \I__4445\ : InMux
    port map (
            O => \N__18864\,
            I => \N__18844\
        );

    \I__4444\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18844\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__18858\,
            I => \N__18837\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__18855\,
            I => \N__18837\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__18852\,
            I => \N__18837\
        );

    \I__4440\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18834\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__18844\,
            I => \N__18827\
        );

    \I__4438\ : Span4Mux_h
    port map (
            O => \N__18837\,
            I => \N__18827\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__18834\,
            I => \N__18827\
        );

    \I__4436\ : Span4Mux_v
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__18824\,
            I => \this_vram.mem_radregZ0Z_12\
        );

    \I__4434\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18815\
        );

    \I__4433\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18815\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__4431\ : Span4Mux_v
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__4430\ : Span4Mux_h
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__4429\ : Odrv4
    port map (
            O => \N__18806\,
            I => \this_vram.mem_N_95\
        );

    \I__4428\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__4426\ : Span4Mux_h
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__4425\ : Sp12to4
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__4424\ : Odrv12
    port map (
            O => \N__18791\,
            I => \this_vram.mem_out_bus6_0\
        );

    \I__4423\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__18779\,
            I => \this_vram.mem_out_bus2_0\
        );

    \I__4419\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__18767\,
            I => \this_vram.mem_out_bus2_1\
        );

    \I__4415\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__4413\ : Span4Mux_v
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__18755\,
            I => \N__18752\
        );

    \I__4411\ : Span4Mux_v
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__18749\,
            I => \this_vram.mem_out_bus6_1\
        );

    \I__4409\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__18743\,
            I => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0_cascade_\
        );

    \I__4406\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18733\
        );

    \I__4405\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18730\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__18733\,
            I => \N__18727\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__18730\,
            I => \N__18724\
        );

    \I__4402\ : Span4Mux_v
    port map (
            O => \N__18727\,
            I => \N__18721\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__18724\,
            I => \N__18718\
        );

    \I__4400\ : Span4Mux_h
    port map (
            O => \N__18721\,
            I => \N__18715\
        );

    \I__4399\ : Span4Mux_h
    port map (
            O => \N__18718\,
            I => \N__18712\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__18715\,
            I => \this_vram.mem_N_91\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__18712\,
            I => \this_vram.mem_N_91\
        );

    \I__4396\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__18704\,
            I => \N__18701\
        );

    \I__4394\ : Sp12to4
    port map (
            O => \N__18701\,
            I => \N__18698\
        );

    \I__4393\ : Odrv12
    port map (
            O => \N__18698\,
            I => \this_vram.mem_out_bus5_1\
        );

    \I__4392\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__4390\ : Sp12to4
    port map (
            O => \N__18689\,
            I => \N__18686\
        );

    \I__4389\ : Span12Mux_v
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__4388\ : Odrv12
    port map (
            O => \N__18683\,
            I => \this_vram.mem_out_bus1_1\
        );

    \I__4387\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__18677\,
            I => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\
        );

    \I__4385\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__18671\,
            I => \this_vram.mem_out_bus3_1\
        );

    \I__4383\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18665\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__18665\,
            I => \N__18662\
        );

    \I__4381\ : Sp12to4
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__4380\ : Span12Mux_v
    port map (
            O => \N__18659\,
            I => \N__18656\
        );

    \I__4379\ : Odrv12
    port map (
            O => \N__18656\,
            I => \this_vram.mem_out_bus7_1\
        );

    \I__4378\ : InMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__18650\,
            I => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\
        );

    \I__4376\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__4374\ : Span4Mux_v
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__4373\ : Odrv4
    port map (
            O => \N__18638\,
            I => \this_vram.mem_out_bus1_0\
        );

    \I__4372\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__4370\ : Span4Mux_v
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__4369\ : Span4Mux_v
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__18623\,
            I => \this_vram.mem_out_bus5_0\
        );

    \I__4367\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__18614\,
            I => \this_vram.mem_out_bus2_3\
        );

    \I__4364\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18608\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__18608\,
            I => \N__18605\
        );

    \I__4362\ : Span4Mux_h
    port map (
            O => \N__18605\,
            I => \N__18602\
        );

    \I__4361\ : Sp12to4
    port map (
            O => \N__18602\,
            I => \N__18599\
        );

    \I__4360\ : Span12Mux_v
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__4359\ : Odrv12
    port map (
            O => \N__18596\,
            I => \this_vram.mem_out_bus6_3\
        );

    \I__4358\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__18590\,
            I => \this_vram.mem_mem_2_1_RNI01N11Z0Z_0\
        );

    \I__4356\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__4354\ : Span4Mux_v
    port map (
            O => \N__18581\,
            I => \N__18578\
        );

    \I__4353\ : Span4Mux_v
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__18575\,
            I => \this_vram.mem_out_bus0_2\
        );

    \I__4351\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__18563\,
            I => \this_vram.mem_out_bus4_2\
        );

    \I__4347\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__18551\,
            I => \this_vram.mem_out_bus1_2\
        );

    \I__4343\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__4341\ : Span4Mux_v
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__18536\,
            I => \this_vram.mem_out_bus5_2\
        );

    \I__4338\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__18521\,
            I => \this_vram.mem_out_bus4_3\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__4332\ : InMux
    port map (
            O => \N__18515\,
            I => \N__18511\
        );

    \I__4331\ : InMux
    port map (
            O => \N__18514\,
            I => \N__18508\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__18511\,
            I => \N__18503\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__18508\,
            I => \N__18503\
        );

    \I__4328\ : Span4Mux_v
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__18497\,
            I => \this_vram.mem_N_88\
        );

    \I__4325\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__18488\,
            I => \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\
        );

    \I__4322\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18481\
        );

    \I__4321\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18478\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__18481\,
            I => \N__18473\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__18478\,
            I => \N__18473\
        );

    \I__4318\ : Span4Mux_v
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__18467\,
            I => \this_vram.mem_N_105\
        );

    \I__4315\ : CEMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__18461\,
            I => \N__18457\
        );

    \I__4313\ : CEMux
    port map (
            O => \N__18460\,
            I => \N__18454\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__18457\,
            I => \N__18451\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__18454\,
            I => \N__18448\
        );

    \I__4310\ : Span4Mux_v
    port map (
            O => \N__18451\,
            I => \N__18445\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__18448\,
            I => \N__18442\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__18445\,
            I => \this_vram.mem_WE_10\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__18442\,
            I => \this_vram.mem_WE_10\
        );

    \I__4306\ : CEMux
    port map (
            O => \N__18437\,
            I => \N__18433\
        );

    \I__4305\ : CEMux
    port map (
            O => \N__18436\,
            I => \N__18430\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__18433\,
            I => \N__18427\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__4301\ : Span12Mux_s2_v
    port map (
            O => \N__18424\,
            I => \N__18418\
        );

    \I__4300\ : Span4Mux_v
    port map (
            O => \N__18421\,
            I => \N__18415\
        );

    \I__4299\ : Span12Mux_v
    port map (
            O => \N__18418\,
            I => \N__18412\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__18415\,
            I => \N__18409\
        );

    \I__4297\ : Odrv12
    port map (
            O => \N__18412\,
            I => \this_vram.mem_WE_14\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__18409\,
            I => \this_vram.mem_WE_14\
        );

    \I__4295\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__4293\ : Span4Mux_v
    port map (
            O => \N__18398\,
            I => \N__18393\
        );

    \I__4292\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18390\
        );

    \I__4291\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18387\
        );

    \I__4290\ : Sp12to4
    port map (
            O => \N__18393\,
            I => \N__18382\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__18390\,
            I => \N__18382\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__18387\,
            I => \N__18379\
        );

    \I__4287\ : Span12Mux_h
    port map (
            O => \N__18382\,
            I => \N__18374\
        );

    \I__4286\ : Span12Mux_v
    port map (
            O => \N__18379\,
            I => \N__18374\
        );

    \I__4285\ : Odrv12
    port map (
            O => \N__18374\,
            I => \this_vram_mem_N_112\
        );

    \I__4284\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18367\
        );

    \I__4283\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18364\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__18367\,
            I => \N__18360\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__18364\,
            I => \N__18355\
        );

    \I__4280\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18352\
        );

    \I__4279\ : Span4Mux_v
    port map (
            O => \N__18360\,
            I => \N__18349\
        );

    \I__4278\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18346\
        );

    \I__4277\ : InMux
    port map (
            O => \N__18358\,
            I => \N__18343\
        );

    \I__4276\ : Span4Mux_v
    port map (
            O => \N__18355\,
            I => \N__18332\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18329\
        );

    \I__4274\ : Sp12to4
    port map (
            O => \N__18349\,
            I => \N__18326\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__18346\,
            I => \N__18323\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__18343\,
            I => \N__18319\
        );

    \I__4271\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18316\
        );

    \I__4270\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18309\
        );

    \I__4269\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18309\
        );

    \I__4268\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18309\
        );

    \I__4267\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18304\
        );

    \I__4266\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18304\
        );

    \I__4265\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18298\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18298\
        );

    \I__4263\ : Sp12to4
    port map (
            O => \N__18332\,
            I => \N__18291\
        );

    \I__4262\ : Span12Mux_v
    port map (
            O => \N__18329\,
            I => \N__18291\
        );

    \I__4261\ : Span12Mux_h
    port map (
            O => \N__18326\,
            I => \N__18288\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__18323\,
            I => \N__18285\
        );

    \I__4259\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18282\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__18319\,
            I => \N__18275\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__18316\,
            I => \N__18275\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__18309\,
            I => \N__18275\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__18304\,
            I => \N__18272\
        );

    \I__4254\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18269\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__18298\,
            I => \N__18266\
        );

    \I__4252\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18263\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18296\,
            I => \N__18260\
        );

    \I__4250\ : Odrv12
    port map (
            O => \N__18291\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4249\ : Odrv12
    port map (
            O => \N__18288\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4248\ : Odrv4
    port map (
            O => \N__18285\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__18282\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__18275\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__18272\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__18269\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__18266\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18263\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18260\,
            I => \this_vga_signals.rgb_1_4\
        );

    \I__4240\ : ClkMux
    port map (
            O => \N__18239\,
            I => \N__18056\
        );

    \I__4239\ : ClkMux
    port map (
            O => \N__18238\,
            I => \N__18056\
        );

    \I__4238\ : ClkMux
    port map (
            O => \N__18237\,
            I => \N__18056\
        );

    \I__4237\ : ClkMux
    port map (
            O => \N__18236\,
            I => \N__18056\
        );

    \I__4236\ : ClkMux
    port map (
            O => \N__18235\,
            I => \N__18056\
        );

    \I__4235\ : ClkMux
    port map (
            O => \N__18234\,
            I => \N__18056\
        );

    \I__4234\ : ClkMux
    port map (
            O => \N__18233\,
            I => \N__18056\
        );

    \I__4233\ : ClkMux
    port map (
            O => \N__18232\,
            I => \N__18056\
        );

    \I__4232\ : ClkMux
    port map (
            O => \N__18231\,
            I => \N__18056\
        );

    \I__4231\ : ClkMux
    port map (
            O => \N__18230\,
            I => \N__18056\
        );

    \I__4230\ : ClkMux
    port map (
            O => \N__18229\,
            I => \N__18056\
        );

    \I__4229\ : ClkMux
    port map (
            O => \N__18228\,
            I => \N__18056\
        );

    \I__4228\ : ClkMux
    port map (
            O => \N__18227\,
            I => \N__18056\
        );

    \I__4227\ : ClkMux
    port map (
            O => \N__18226\,
            I => \N__18056\
        );

    \I__4226\ : ClkMux
    port map (
            O => \N__18225\,
            I => \N__18056\
        );

    \I__4225\ : ClkMux
    port map (
            O => \N__18224\,
            I => \N__18056\
        );

    \I__4224\ : ClkMux
    port map (
            O => \N__18223\,
            I => \N__18056\
        );

    \I__4223\ : ClkMux
    port map (
            O => \N__18222\,
            I => \N__18056\
        );

    \I__4222\ : ClkMux
    port map (
            O => \N__18221\,
            I => \N__18056\
        );

    \I__4221\ : ClkMux
    port map (
            O => \N__18220\,
            I => \N__18056\
        );

    \I__4220\ : ClkMux
    port map (
            O => \N__18219\,
            I => \N__18056\
        );

    \I__4219\ : ClkMux
    port map (
            O => \N__18218\,
            I => \N__18056\
        );

    \I__4218\ : ClkMux
    port map (
            O => \N__18217\,
            I => \N__18056\
        );

    \I__4217\ : ClkMux
    port map (
            O => \N__18216\,
            I => \N__18056\
        );

    \I__4216\ : ClkMux
    port map (
            O => \N__18215\,
            I => \N__18056\
        );

    \I__4215\ : ClkMux
    port map (
            O => \N__18214\,
            I => \N__18056\
        );

    \I__4214\ : ClkMux
    port map (
            O => \N__18213\,
            I => \N__18056\
        );

    \I__4213\ : ClkMux
    port map (
            O => \N__18212\,
            I => \N__18056\
        );

    \I__4212\ : ClkMux
    port map (
            O => \N__18211\,
            I => \N__18056\
        );

    \I__4211\ : ClkMux
    port map (
            O => \N__18210\,
            I => \N__18056\
        );

    \I__4210\ : ClkMux
    port map (
            O => \N__18209\,
            I => \N__18056\
        );

    \I__4209\ : ClkMux
    port map (
            O => \N__18208\,
            I => \N__18056\
        );

    \I__4208\ : ClkMux
    port map (
            O => \N__18207\,
            I => \N__18056\
        );

    \I__4207\ : ClkMux
    port map (
            O => \N__18206\,
            I => \N__18056\
        );

    \I__4206\ : ClkMux
    port map (
            O => \N__18205\,
            I => \N__18056\
        );

    \I__4205\ : ClkMux
    port map (
            O => \N__18204\,
            I => \N__18056\
        );

    \I__4204\ : ClkMux
    port map (
            O => \N__18203\,
            I => \N__18056\
        );

    \I__4203\ : ClkMux
    port map (
            O => \N__18202\,
            I => \N__18056\
        );

    \I__4202\ : ClkMux
    port map (
            O => \N__18201\,
            I => \N__18056\
        );

    \I__4201\ : ClkMux
    port map (
            O => \N__18200\,
            I => \N__18056\
        );

    \I__4200\ : ClkMux
    port map (
            O => \N__18199\,
            I => \N__18056\
        );

    \I__4199\ : ClkMux
    port map (
            O => \N__18198\,
            I => \N__18056\
        );

    \I__4198\ : ClkMux
    port map (
            O => \N__18197\,
            I => \N__18056\
        );

    \I__4197\ : ClkMux
    port map (
            O => \N__18196\,
            I => \N__18056\
        );

    \I__4196\ : ClkMux
    port map (
            O => \N__18195\,
            I => \N__18056\
        );

    \I__4195\ : ClkMux
    port map (
            O => \N__18194\,
            I => \N__18056\
        );

    \I__4194\ : ClkMux
    port map (
            O => \N__18193\,
            I => \N__18056\
        );

    \I__4193\ : ClkMux
    port map (
            O => \N__18192\,
            I => \N__18056\
        );

    \I__4192\ : ClkMux
    port map (
            O => \N__18191\,
            I => \N__18056\
        );

    \I__4191\ : ClkMux
    port map (
            O => \N__18190\,
            I => \N__18056\
        );

    \I__4190\ : ClkMux
    port map (
            O => \N__18189\,
            I => \N__18056\
        );

    \I__4189\ : ClkMux
    port map (
            O => \N__18188\,
            I => \N__18056\
        );

    \I__4188\ : ClkMux
    port map (
            O => \N__18187\,
            I => \N__18056\
        );

    \I__4187\ : ClkMux
    port map (
            O => \N__18186\,
            I => \N__18056\
        );

    \I__4186\ : ClkMux
    port map (
            O => \N__18185\,
            I => \N__18056\
        );

    \I__4185\ : ClkMux
    port map (
            O => \N__18184\,
            I => \N__18056\
        );

    \I__4184\ : ClkMux
    port map (
            O => \N__18183\,
            I => \N__18056\
        );

    \I__4183\ : ClkMux
    port map (
            O => \N__18182\,
            I => \N__18056\
        );

    \I__4182\ : ClkMux
    port map (
            O => \N__18181\,
            I => \N__18056\
        );

    \I__4181\ : ClkMux
    port map (
            O => \N__18180\,
            I => \N__18056\
        );

    \I__4180\ : ClkMux
    port map (
            O => \N__18179\,
            I => \N__18056\
        );

    \I__4179\ : GlobalMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__4178\ : gio2CtrlBuf
    port map (
            O => \N__18053\,
            I => clk_0_c_g
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \N__18046\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18040\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18040\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18045\,
            I => \N__18037\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18040\,
            I => \N__18034\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__18037\,
            I => \N__18031\
        );

    \I__4171\ : Sp12to4
    port map (
            O => \N__18034\,
            I => \N__18028\
        );

    \I__4170\ : Span4Mux_v
    port map (
            O => \N__18031\,
            I => \N__18025\
        );

    \I__4169\ : Span12Mux_v
    port map (
            O => \N__18028\,
            I => \N__18022\
        );

    \I__4168\ : Sp12to4
    port map (
            O => \N__18025\,
            I => \N__18019\
        );

    \I__4167\ : Span12Mux_h
    port map (
            O => \N__18022\,
            I => \N__18016\
        );

    \I__4166\ : Span12Mux_h
    port map (
            O => \N__18019\,
            I => \N__18013\
        );

    \I__4165\ : Odrv12
    port map (
            O => \N__18016\,
            I => port_data_c_3
        );

    \I__4164\ : Odrv12
    port map (
            O => \N__18013\,
            I => port_data_c_3
        );

    \I__4163\ : InMux
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__18005\,
            I => \N__18000\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17997\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17993\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__18000\,
            I => \N__17989\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__17997\,
            I => \N__17986\
        );

    \I__4157\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17983\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__17993\,
            I => \N__17979\
        );

    \I__4155\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17976\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__17989\,
            I => \N__17971\
        );

    \I__4153\ : Span4Mux_h
    port map (
            O => \N__17986\,
            I => \N__17971\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__17983\,
            I => \N__17968\
        );

    \I__4151\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17965\
        );

    \I__4150\ : Span4Mux_h
    port map (
            O => \N__17979\,
            I => \N__17960\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__17976\,
            I => \N__17957\
        );

    \I__4148\ : Span4Mux_v
    port map (
            O => \N__17971\,
            I => \N__17952\
        );

    \I__4147\ : Span4Mux_h
    port map (
            O => \N__17968\,
            I => \N__17952\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__17965\,
            I => \N__17949\
        );

    \I__4145\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17946\
        );

    \I__4144\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17943\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__17960\,
            I => \N__17938\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__17957\,
            I => \N__17938\
        );

    \I__4141\ : Span4Mux_v
    port map (
            O => \N__17952\,
            I => \N__17933\
        );

    \I__4140\ : Span4Mux_h
    port map (
            O => \N__17949\,
            I => \N__17933\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__17946\,
            I => \N__17930\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__17943\,
            I => \N__17927\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__17938\,
            I => \N__17918\
        );

    \I__4136\ : Span4Mux_v
    port map (
            O => \N__17933\,
            I => \N__17918\
        );

    \I__4135\ : Span4Mux_h
    port map (
            O => \N__17930\,
            I => \N__17918\
        );

    \I__4134\ : Span4Mux_h
    port map (
            O => \N__17927\,
            I => \N__17918\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__17918\,
            I => \M_this_vram_write_data_3\
        );

    \I__4132\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__17906\,
            I => \this_vram.mem_out_bus4_1\
        );

    \I__4128\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17900\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__17900\,
            I => \N__17897\
        );

    \I__4126\ : Span4Mux_v
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__4125\ : Span4Mux_v
    port map (
            O => \N__17894\,
            I => \N__17891\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__17891\,
            I => \this_vram.mem_out_bus0_1\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__17888\,
            I => \rgbZ0Z_1_cascade_\
        );

    \I__4122\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17882\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__17882\,
            I => \M_vcounter_q_esr_RNI2RH6LA_9\
        );

    \I__4120\ : InMux
    port map (
            O => \N__17879\,
            I => \N__17875\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__17878\,
            I => \N__17870\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__17875\,
            I => \N__17866\
        );

    \I__4117\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17862\
        );

    \I__4116\ : InMux
    port map (
            O => \N__17873\,
            I => \N__17859\
        );

    \I__4115\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17854\
        );

    \I__4114\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17854\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__17866\,
            I => \N__17850\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__17865\,
            I => \N__17847\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__17862\,
            I => \N__17843\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__17859\,
            I => \N__17840\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__17854\,
            I => \N__17837\
        );

    \I__4108\ : CascadeMux
    port map (
            O => \N__17853\,
            I => \N__17834\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__17850\,
            I => \N__17828\
        );

    \I__4106\ : InMux
    port map (
            O => \N__17847\,
            I => \N__17823\
        );

    \I__4105\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17823\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__17843\,
            I => \N__17816\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__17840\,
            I => \N__17816\
        );

    \I__4102\ : Span4Mux_h
    port map (
            O => \N__17837\,
            I => \N__17816\
        );

    \I__4101\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17809\
        );

    \I__4100\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17809\
        );

    \I__4099\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17809\
        );

    \I__4098\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17806\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__17828\,
            I => \rgbZ0Z_1\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__17823\,
            I => \rgbZ0Z_1\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__17816\,
            I => \rgbZ0Z_1\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__17809\,
            I => \rgbZ0Z_1\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__17806\,
            I => \rgbZ0Z_1\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__4091\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__17789\,
            I => \N__17786\
        );

    \I__4089\ : Odrv12
    port map (
            O => \N__17786\,
            I => \M_vcounter_q_esr_RNIVLNKSA_9\
        );

    \I__4088\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17780\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__17780\,
            I => \N__17776\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__17779\,
            I => \N__17771\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__17776\,
            I => \N__17766\
        );

    \I__4084\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17763\
        );

    \I__4083\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17754\
        );

    \I__4082\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17754\
        );

    \I__4081\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17754\
        );

    \I__4080\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17754\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__17766\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__17763\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__17754\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__17747\,
            I => \N__17744\
        );

    \I__4075\ : CascadeBuf
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__17741\,
            I => \N__17738\
        );

    \I__4073\ : CascadeBuf
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__17735\,
            I => \N__17732\
        );

    \I__4071\ : CascadeBuf
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__4069\ : CascadeBuf
    port map (
            O => \N__17726\,
            I => \N__17723\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__17723\,
            I => \N__17720\
        );

    \I__4067\ : CascadeBuf
    port map (
            O => \N__17720\,
            I => \N__17717\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__4065\ : CascadeBuf
    port map (
            O => \N__17714\,
            I => \N__17711\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__4063\ : CascadeBuf
    port map (
            O => \N__17708\,
            I => \N__17705\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__17705\,
            I => \N__17702\
        );

    \I__4061\ : CascadeBuf
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__4059\ : CascadeBuf
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__17693\,
            I => \N__17690\
        );

    \I__4057\ : CascadeBuf
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__4056\ : CascadeMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__4055\ : CascadeBuf
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__4054\ : CascadeMux
    port map (
            O => \N__17681\,
            I => \N__17678\
        );

    \I__4053\ : CascadeBuf
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__17675\,
            I => \N__17672\
        );

    \I__4051\ : CascadeBuf
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__17669\,
            I => \N__17666\
        );

    \I__4049\ : CascadeBuf
    port map (
            O => \N__17666\,
            I => \N__17663\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__17663\,
            I => \N__17660\
        );

    \I__4047\ : CascadeBuf
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__4045\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17651\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__17651\,
            I => \N__17648\
        );

    \I__4043\ : Span4Mux_h
    port map (
            O => \N__17648\,
            I => \N__17644\
        );

    \I__4042\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17641\
        );

    \I__4041\ : Span4Mux_v
    port map (
            O => \N__17644\,
            I => \N__17638\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__17641\,
            I => \N__17635\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__17638\,
            I => \N__17632\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__17635\,
            I => \M_this_vga_signals_address_3\
        );

    \I__4037\ : Odrv4
    port map (
            O => \N__17632\,
            I => \M_this_vga_signals_address_3\
        );

    \I__4036\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17624\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__17624\,
            I => \N__17619\
        );

    \I__4034\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17616\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__17622\,
            I => \N__17613\
        );

    \I__4032\ : Span4Mux_v
    port map (
            O => \N__17619\,
            I => \N__17610\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__17616\,
            I => \N__17607\
        );

    \I__4030\ : InMux
    port map (
            O => \N__17613\,
            I => \N__17604\
        );

    \I__4029\ : Sp12to4
    port map (
            O => \N__17610\,
            I => \N__17601\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__17607\,
            I => \N__17598\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__17604\,
            I => \N__17595\
        );

    \I__4026\ : Span12Mux_h
    port map (
            O => \N__17601\,
            I => \N__17590\
        );

    \I__4025\ : Sp12to4
    port map (
            O => \N__17598\,
            I => \N__17590\
        );

    \I__4024\ : Span12Mux_v
    port map (
            O => \N__17595\,
            I => \N__17587\
        );

    \I__4023\ : Odrv12
    port map (
            O => \N__17590\,
            I => port_data_c_0
        );

    \I__4022\ : Odrv12
    port map (
            O => \N__17587\,
            I => port_data_c_0
        );

    \I__4021\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17578\
        );

    \I__4020\ : InMux
    port map (
            O => \N__17581\,
            I => \N__17574\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17569\
        );

    \I__4018\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17566\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__17574\,
            I => \N__17562\
        );

    \I__4016\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17559\
        );

    \I__4015\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17556\
        );

    \I__4014\ : Span4Mux_s3_v
    port map (
            O => \N__17569\,
            I => \N__17550\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__17566\,
            I => \N__17550\
        );

    \I__4012\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17547\
        );

    \I__4011\ : Span4Mux_h
    port map (
            O => \N__17562\,
            I => \N__17544\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__17559\,
            I => \N__17541\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__17556\,
            I => \N__17538\
        );

    \I__4008\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17535\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__17550\,
            I => \N__17530\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__17547\,
            I => \N__17530\
        );

    \I__4005\ : Span4Mux_v
    port map (
            O => \N__17544\,
            I => \N__17525\
        );

    \I__4004\ : Span4Mux_h
    port map (
            O => \N__17541\,
            I => \N__17525\
        );

    \I__4003\ : Span4Mux_v
    port map (
            O => \N__17538\,
            I => \N__17520\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__17535\,
            I => \N__17520\
        );

    \I__4001\ : Sp12to4
    port map (
            O => \N__17530\,
            I => \N__17516\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__17525\,
            I => \N__17511\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__17520\,
            I => \N__17511\
        );

    \I__3998\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17508\
        );

    \I__3997\ : Span12Mux_v
    port map (
            O => \N__17516\,
            I => \N__17501\
        );

    \I__3996\ : Sp12to4
    port map (
            O => \N__17511\,
            I => \N__17501\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__17508\,
            I => \N__17501\
        );

    \I__3994\ : Odrv12
    port map (
            O => \N__17501\,
            I => \M_this_vram_write_data_0\
        );

    \I__3993\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17495\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__3991\ : Span4Mux_h
    port map (
            O => \N__17492\,
            I => \N__17489\
        );

    \I__3990\ : Span4Mux_h
    port map (
            O => \N__17489\,
            I => \N__17486\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__17486\,
            I => \this_vga_signals.SUM_3_1\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__17483\,
            I => \N__17480\
        );

    \I__3987\ : CascadeBuf
    port map (
            O => \N__17480\,
            I => \N__17477\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__17477\,
            I => \N__17474\
        );

    \I__3985\ : CascadeBuf
    port map (
            O => \N__17474\,
            I => \N__17471\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__17471\,
            I => \N__17468\
        );

    \I__3983\ : CascadeBuf
    port map (
            O => \N__17468\,
            I => \N__17465\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__17465\,
            I => \N__17462\
        );

    \I__3981\ : CascadeBuf
    port map (
            O => \N__17462\,
            I => \N__17459\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__3979\ : CascadeBuf
    port map (
            O => \N__17456\,
            I => \N__17453\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__3977\ : CascadeBuf
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__17447\,
            I => \N__17444\
        );

    \I__3975\ : CascadeBuf
    port map (
            O => \N__17444\,
            I => \N__17441\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__17441\,
            I => \N__17438\
        );

    \I__3973\ : CascadeBuf
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3971\ : CascadeBuf
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__3969\ : CascadeBuf
    port map (
            O => \N__17426\,
            I => \N__17423\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__17423\,
            I => \N__17420\
        );

    \I__3967\ : CascadeBuf
    port map (
            O => \N__17420\,
            I => \N__17417\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__3965\ : CascadeBuf
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__3963\ : CascadeBuf
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__3961\ : CascadeBuf
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3960\ : CascadeMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3959\ : CascadeBuf
    port map (
            O => \N__17396\,
            I => \N__17393\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__17393\,
            I => \N__17390\
        );

    \I__3957\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__3955\ : Span4Mux_v
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__3954\ : Span4Mux_h
    port map (
            O => \N__17381\,
            I => \N__17378\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__17378\,
            I => \M_this_vga_signals_address_6\
        );

    \I__3952\ : CEMux
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__17372\,
            I => \N__17368\
        );

    \I__3950\ : CEMux
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__17368\,
            I => \N__17360\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__17365\,
            I => \N__17360\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__17360\,
            I => \N__17357\
        );

    \I__3946\ : Span4Mux_v
    port map (
            O => \N__17357\,
            I => \N__17354\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__17354\,
            I => \this_vram.mem_WE_12\
        );

    \I__3944\ : InMux
    port map (
            O => \N__17351\,
            I => \N__17346\
        );

    \I__3943\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17343\
        );

    \I__3942\ : InMux
    port map (
            O => \N__17349\,
            I => \N__17340\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__17346\,
            I => \N__17334\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__17343\,
            I => \N__17334\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17331\
        );

    \I__3938\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17328\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__17334\,
            I => \N__17323\
        );

    \I__3936\ : Span4Mux_h
    port map (
            O => \N__17331\,
            I => \N__17323\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__17328\,
            I => \N__17315\
        );

    \I__3934\ : Span4Mux_h
    port map (
            O => \N__17323\,
            I => \N__17312\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17305\
        );

    \I__3932\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17305\
        );

    \I__3931\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17302\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__17319\,
            I => \N__17295\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__17318\,
            I => \N__17292\
        );

    \I__3928\ : Span12Mux_h
    port map (
            O => \N__17315\,
            I => \N__17289\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__17312\,
            I => \N__17286\
        );

    \I__3926\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17281\
        );

    \I__3925\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17281\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__17305\,
            I => \N__17278\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17302\,
            I => \N__17275\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17301\,
            I => \N__17266\
        );

    \I__3921\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17266\
        );

    \I__3920\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17266\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17266\
        );

    \I__3918\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17263\
        );

    \I__3917\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17260\
        );

    \I__3916\ : Odrv12
    port map (
            O => \N__17289\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__17286\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__17281\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__17278\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__17275\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__17266\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__17263\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__17260\,
            I => \this_vga_signals.rgb_1_2\
        );

    \I__3908\ : CEMux
    port map (
            O => \N__17243\,
            I => \N__17239\
        );

    \I__3907\ : CEMux
    port map (
            O => \N__17242\,
            I => \N__17236\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__17239\,
            I => \N__17233\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__17236\,
            I => \N__17230\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__17233\,
            I => \N__17227\
        );

    \I__3903\ : Span4Mux_h
    port map (
            O => \N__17230\,
            I => \N__17224\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__17227\,
            I => \this_vram.mem_WE_8\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__17224\,
            I => \this_vram.mem_WE_8\
        );

    \I__3900\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__3898\ : Span4Mux_v
    port map (
            O => \N__17213\,
            I => \N__17210\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__17207\,
            I => \N__17204\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__17204\,
            I => \this_vram.mem_out_bus0_3\
        );

    \I__3894\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17194\
        );

    \I__3893\ : InMux
    port map (
            O => \N__17200\,
            I => \N__17191\
        );

    \I__3892\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17188\
        );

    \I__3891\ : InMux
    port map (
            O => \N__17198\,
            I => \N__17182\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17182\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17194\,
            I => \N__17171\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__17191\,
            I => \N__17171\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17188\,
            I => \N__17171\
        );

    \I__3886\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17165\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17182\,
            I => \N__17155\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17181\,
            I => \N__17152\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17145\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17145\
        );

    \I__3881\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17145\
        );

    \I__3880\ : Span4Mux_v
    port map (
            O => \N__17171\,
            I => \N__17142\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17139\
        );

    \I__3878\ : InMux
    port map (
            O => \N__17169\,
            I => \N__17136\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17133\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17129\
        );

    \I__3875\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17126\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17119\
        );

    \I__3873\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17119\
        );

    \I__3872\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17119\
        );

    \I__3871\ : CascadeMux
    port map (
            O => \N__17160\,
            I => \N__17112\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__17159\,
            I => \N__17107\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__17158\,
            I => \N__17104\
        );

    \I__3868\ : Span4Mux_h
    port map (
            O => \N__17155\,
            I => \N__17094\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__17152\,
            I => \N__17094\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17145\,
            I => \N__17094\
        );

    \I__3865\ : Sp12to4
    port map (
            O => \N__17142\,
            I => \N__17087\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__17139\,
            I => \N__17087\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__17136\,
            I => \N__17087\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__17133\,
            I => \N__17084\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17081\
        );

    \I__3860\ : Span4Mux_v
    port map (
            O => \N__17129\,
            I => \N__17074\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17126\,
            I => \N__17074\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__17119\,
            I => \N__17074\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17071\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17064\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17064\
        );

    \I__3854\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17064\
        );

    \I__3853\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17059\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17059\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17050\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17050\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17050\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17103\,
            I => \N__17050\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17045\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17045\
        );

    \I__3845\ : Span4Mux_h
    port map (
            O => \N__17094\,
            I => \N__17042\
        );

    \I__3844\ : Odrv12
    port map (
            O => \N__17087\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__17084\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17081\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__17074\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__17071\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17064\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__17059\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__17050\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__17045\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__17042\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__17015\,
            I => \rgb_1_cry_0_0_c_RNOZ0Z_0\
        );

    \I__3831\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17009\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__17009\,
            I => \M_vcounter_q_esr_RNI1H9RHL_9\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__3828\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16994\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16994\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16987\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16987\
        );

    \I__3824\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16987\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__16994\,
            I => \N__16979\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__16987\,
            I => \N__16979\
        );

    \I__3821\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16972\
        );

    \I__3820\ : InMux
    port map (
            O => \N__16985\,
            I => \N__16972\
        );

    \I__3819\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16972\
        );

    \I__3818\ : Span4Mux_v
    port map (
            O => \N__16979\,
            I => \N__16963\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__16972\,
            I => \N__16960\
        );

    \I__3816\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16951\
        );

    \I__3815\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16951\
        );

    \I__3814\ : InMux
    port map (
            O => \N__16969\,
            I => \N__16951\
        );

    \I__3813\ : InMux
    port map (
            O => \N__16968\,
            I => \N__16951\
        );

    \I__3812\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16948\
        );

    \I__3811\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16945\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__16963\,
            I => rgb_1_3
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__16960\,
            I => rgb_1_3
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__16951\,
            I => rgb_1_3
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__16948\,
            I => rgb_1_3
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__16945\,
            I => rgb_1_3
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__16934\,
            I => \N__16928\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__16933\,
            I => \N__16925\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__16932\,
            I => \N__16921\
        );

    \I__3802\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16916\
        );

    \I__3801\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16916\
        );

    \I__3800\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16909\
        );

    \I__3799\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16909\
        );

    \I__3798\ : InMux
    port map (
            O => \N__16921\,
            I => \N__16909\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__16916\,
            I => \N__16898\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__16909\,
            I => \N__16898\
        );

    \I__3795\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16891\
        );

    \I__3794\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16891\
        );

    \I__3793\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16891\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__16905\,
            I => \N__16888\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__16904\,
            I => \N__16884\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__16903\,
            I => \N__16881\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__16898\,
            I => \N__16876\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__16891\,
            I => \N__16873\
        );

    \I__3787\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16864\
        );

    \I__3786\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16864\
        );

    \I__3785\ : InMux
    port map (
            O => \N__16884\,
            I => \N__16864\
        );

    \I__3784\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16864\
        );

    \I__3783\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16861\
        );

    \I__3782\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16858\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__16876\,
            I => rgb_1_4
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__16873\,
            I => rgb_1_4
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__16864\,
            I => rgb_1_4
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__16861\,
            I => rgb_1_4
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__16858\,
            I => rgb_1_4
        );

    \I__3776\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16837\
        );

    \I__3775\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16837\
        );

    \I__3774\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16830\
        );

    \I__3773\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16830\
        );

    \I__3772\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16830\
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__16842\,
            I => \N__16827\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__16837\,
            I => \N__16818\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__16830\,
            I => \N__16818\
        );

    \I__3768\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16811\
        );

    \I__3767\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16811\
        );

    \I__3766\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16811\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__16824\,
            I => \N__16804\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__16823\,
            I => \N__16801\
        );

    \I__3763\ : Span4Mux_v
    port map (
            O => \N__16818\,
            I => \N__16798\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__16811\,
            I => \N__16795\
        );

    \I__3761\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16786\
        );

    \I__3760\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16786\
        );

    \I__3759\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16786\
        );

    \I__3758\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16786\
        );

    \I__3757\ : InMux
    port map (
            O => \N__16804\,
            I => \N__16783\
        );

    \I__3756\ : InMux
    port map (
            O => \N__16801\,
            I => \N__16780\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__16798\,
            I => rgb_1_5
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__16795\,
            I => rgb_1_5
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__16786\,
            I => rgb_1_5
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__16783\,
            I => rgb_1_5
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__16780\,
            I => rgb_1_5
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__16769\,
            I => \N__16763\
        );

    \I__3749\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16755\
        );

    \I__3748\ : InMux
    port map (
            O => \N__16767\,
            I => \N__16755\
        );

    \I__3747\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16748\
        );

    \I__3746\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16748\
        );

    \I__3745\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16748\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__16761\,
            I => \N__16744\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__16760\,
            I => \N__16741\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__16755\,
            I => \N__16735\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__16748\,
            I => \N__16735\
        );

    \I__3740\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16728\
        );

    \I__3739\ : InMux
    port map (
            O => \N__16744\,
            I => \N__16728\
        );

    \I__3738\ : InMux
    port map (
            O => \N__16741\,
            I => \N__16728\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__16740\,
            I => \N__16724\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__16735\,
            I => \N__16717\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__16728\,
            I => \N__16714\
        );

    \I__3734\ : InMux
    port map (
            O => \N__16727\,
            I => \N__16705\
        );

    \I__3733\ : InMux
    port map (
            O => \N__16724\,
            I => \N__16705\
        );

    \I__3732\ : InMux
    port map (
            O => \N__16723\,
            I => \N__16705\
        );

    \I__3731\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16705\
        );

    \I__3730\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16702\
        );

    \I__3729\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16699\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__16717\,
            I => \rgb_1_6_THRU_CO\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__16714\,
            I => \rgb_1_6_THRU_CO\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__16705\,
            I => \rgb_1_6_THRU_CO\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__16702\,
            I => \rgb_1_6_THRU_CO\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__16699\,
            I => \rgb_1_6_THRU_CO\
        );

    \I__3723\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16682\
        );

    \I__3722\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16682\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__16682\,
            I => m36
        );

    \I__3720\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16675\
        );

    \I__3719\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16672\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__16675\,
            I => \N__16669\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__16672\,
            I => \N__16666\
        );

    \I__3716\ : Span12Mux_h
    port map (
            O => \N__16669\,
            I => \N__16663\
        );

    \I__3715\ : Span12Mux_v
    port map (
            O => \N__16666\,
            I => \N__16660\
        );

    \I__3714\ : Odrv12
    port map (
            O => \N__16663\,
            I => port_address_c_0
        );

    \I__3713\ : Odrv12
    port map (
            O => \N__16660\,
            I => port_address_c_0
        );

    \I__3712\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3710\ : Span12Mux_h
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3709\ : Odrv12
    port map (
            O => \N__16646\,
            I => port_address_c_1
        );

    \I__3708\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__16640\,
            I => \M_state_q_ns_0_a3_0_1_1\
        );

    \I__3706\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16632\
        );

    \I__3705\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16629\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__16635\,
            I => \N__16626\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__16632\,
            I => \N__16623\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__16629\,
            I => \N__16620\
        );

    \I__3701\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16617\
        );

    \I__3700\ : Span4Mux_h
    port map (
            O => \N__16623\,
            I => \N__16614\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__16620\,
            I => \N__16611\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__16617\,
            I => \N__16608\
        );

    \I__3697\ : Span4Mux_v
    port map (
            O => \N__16614\,
            I => \N__16605\
        );

    \I__3696\ : Span4Mux_v
    port map (
            O => \N__16611\,
            I => \N__16602\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__16608\,
            I => \N__16599\
        );

    \I__3694\ : Span4Mux_v
    port map (
            O => \N__16605\,
            I => \N__16596\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__16602\,
            I => \N__16593\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__16599\,
            I => \N__16590\
        );

    \I__3691\ : Span4Mux_h
    port map (
            O => \N__16596\,
            I => \N__16587\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__16593\,
            I => \N__16584\
        );

    \I__3689\ : Span4Mux_v
    port map (
            O => \N__16590\,
            I => \N__16581\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__16587\,
            I => port_data_c_1
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__16584\,
            I => port_data_c_1
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__16581\,
            I => port_data_c_1
        );

    \I__3685\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__16571\,
            I => \N__16567\
        );

    \I__3683\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16564\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__16567\,
            I => \N__16561\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__16564\,
            I => \N__16558\
        );

    \I__3680\ : Span4Mux_v
    port map (
            O => \N__16561\,
            I => \N__16551\
        );

    \I__3679\ : Span4Mux_h
    port map (
            O => \N__16558\,
            I => \N__16551\
        );

    \I__3678\ : InMux
    port map (
            O => \N__16557\,
            I => \N__16548\
        );

    \I__3677\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16543\
        );

    \I__3676\ : Span4Mux_v
    port map (
            O => \N__16551\,
            I => \N__16539\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16536\
        );

    \I__3674\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16533\
        );

    \I__3673\ : InMux
    port map (
            O => \N__16546\,
            I => \N__16530\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__16543\,
            I => \N__16527\
        );

    \I__3671\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16524\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__16539\,
            I => \N__16519\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__16536\,
            I => \N__16519\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__16533\,
            I => \N__16516\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__16530\,
            I => \N__16513\
        );

    \I__3666\ : Span4Mux_v
    port map (
            O => \N__16527\,
            I => \N__16508\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__16524\,
            I => \N__16508\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__16519\,
            I => \N__16502\
        );

    \I__3663\ : Span4Mux_h
    port map (
            O => \N__16516\,
            I => \N__16502\
        );

    \I__3662\ : Span12Mux_h
    port map (
            O => \N__16513\,
            I => \N__16499\
        );

    \I__3661\ : Span4Mux_v
    port map (
            O => \N__16508\,
            I => \N__16496\
        );

    \I__3660\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16493\
        );

    \I__3659\ : Span4Mux_h
    port map (
            O => \N__16502\,
            I => \N__16490\
        );

    \I__3658\ : Span12Mux_v
    port map (
            O => \N__16499\,
            I => \N__16483\
        );

    \I__3657\ : Sp12to4
    port map (
            O => \N__16496\,
            I => \N__16483\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__16493\,
            I => \N__16483\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__16490\,
            I => \M_this_vram_write_data_1\
        );

    \I__3654\ : Odrv12
    port map (
            O => \N__16483\,
            I => \M_this_vram_write_data_1\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__16478\,
            I => \N__16474\
        );

    \I__3652\ : InMux
    port map (
            O => \N__16477\,
            I => \N__16466\
        );

    \I__3651\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16466\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16463\
        );

    \I__3649\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16457\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16454\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__16466\,
            I => \N__16444\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16444\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16439\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16439\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16433\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__16457\,
            I => \N__16430\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__16454\,
            I => \N__16427\
        );

    \I__3640\ : InMux
    port map (
            O => \N__16453\,
            I => \N__16422\
        );

    \I__3639\ : InMux
    port map (
            O => \N__16452\,
            I => \N__16422\
        );

    \I__3638\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16419\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16414\
        );

    \I__3636\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16414\
        );

    \I__3635\ : Span4Mux_v
    port map (
            O => \N__16444\,
            I => \N__16411\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__16439\,
            I => \N__16408\
        );

    \I__3633\ : InMux
    port map (
            O => \N__16438\,
            I => \N__16401\
        );

    \I__3632\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16401\
        );

    \I__3631\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16401\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__16433\,
            I => \N__16396\
        );

    \I__3629\ : Span4Mux_h
    port map (
            O => \N__16430\,
            I => \N__16396\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__16427\,
            I => \N__16391\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__16422\,
            I => \N__16391\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__16419\,
            I => \N_349_0\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__16414\,
            I => \N_349_0\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__16411\,
            I => \N_349_0\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__16408\,
            I => \N_349_0\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__16401\,
            I => \N_349_0\
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__16396\,
            I => \N_349_0\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__16391\,
            I => \N_349_0\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__16376\,
            I => \N__16372\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__16375\,
            I => \N__16369\
        );

    \I__3617\ : InMux
    port map (
            O => \N__16372\,
            I => \N__16366\
        );

    \I__3616\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16363\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__16366\,
            I => \N__16360\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__16363\,
            I => \N__16357\
        );

    \I__3613\ : Span4Mux_v
    port map (
            O => \N__16360\,
            I => \N__16354\
        );

    \I__3612\ : Span4Mux_v
    port map (
            O => \N__16357\,
            I => \N__16351\
        );

    \I__3611\ : Sp12to4
    port map (
            O => \N__16354\,
            I => \N__16348\
        );

    \I__3610\ : Sp12to4
    port map (
            O => \N__16351\,
            I => \N__16345\
        );

    \I__3609\ : Span12Mux_h
    port map (
            O => \N__16348\,
            I => \N__16342\
        );

    \I__3608\ : Span12Mux_h
    port map (
            O => \N__16345\,
            I => \N__16339\
        );

    \I__3607\ : Span12Mux_v
    port map (
            O => \N__16342\,
            I => \N__16336\
        );

    \I__3606\ : Span12Mux_v
    port map (
            O => \N__16339\,
            I => \N__16333\
        );

    \I__3605\ : Odrv12
    port map (
            O => \N__16336\,
            I => port_data_c_6
        );

    \I__3604\ : Odrv12
    port map (
            O => \N__16333\,
            I => port_data_c_6
        );

    \I__3603\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16322\
        );

    \I__3602\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16306\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16303\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__16325\,
            I => \N__16291\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16322\,
            I => \N__16288\
        );

    \I__3598\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16281\
        );

    \I__3597\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16270\
        );

    \I__3596\ : InMux
    port map (
            O => \N__16319\,
            I => \N__16270\
        );

    \I__3595\ : InMux
    port map (
            O => \N__16318\,
            I => \N__16270\
        );

    \I__3594\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16270\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16270\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16315\,
            I => \N__16267\
        );

    \I__3591\ : InMux
    port map (
            O => \N__16314\,
            I => \N__16258\
        );

    \I__3590\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16258\
        );

    \I__3589\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16258\
        );

    \I__3588\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16258\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__16310\,
            I => \N__16255\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16309\,
            I => \N__16252\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__16306\,
            I => \N__16247\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__16303\,
            I => \N__16247\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16242\
        );

    \I__3582\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16242\
        );

    \I__3581\ : InMux
    port map (
            O => \N__16300\,
            I => \N__16235\
        );

    \I__3580\ : InMux
    port map (
            O => \N__16299\,
            I => \N__16235\
        );

    \I__3579\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16224\
        );

    \I__3578\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16224\
        );

    \I__3577\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16224\
        );

    \I__3576\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16224\
        );

    \I__3575\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16224\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16221\
        );

    \I__3573\ : Span4Mux_h
    port map (
            O => \N__16288\,
            I => \N__16218\
        );

    \I__3572\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16215\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16208\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16208\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16208\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__16281\,
            I => \N__16199\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__16270\,
            I => \N__16199\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16267\,
            I => \N__16199\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__16258\,
            I => \N__16199\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16196\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__16252\,
            I => \N__16193\
        );

    \I__3562\ : Span4Mux_v
    port map (
            O => \N__16247\,
            I => \N__16188\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__16242\,
            I => \N__16188\
        );

    \I__3560\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16183\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16183\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16235\,
            I => \M_state_qZ0Z_0\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__16224\,
            I => \M_state_qZ0Z_0\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__16221\,
            I => \M_state_qZ0Z_0\
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__16218\,
            I => \M_state_qZ0Z_0\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__16215\,
            I => \M_state_qZ0Z_0\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__16208\,
            I => \M_state_qZ0Z_0\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__16199\,
            I => \M_state_qZ0Z_0\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16196\,
            I => \M_state_qZ0Z_0\
        );

    \I__3550\ : Odrv4
    port map (
            O => \N__16193\,
            I => \M_state_qZ0Z_0\
        );

    \I__3549\ : Odrv4
    port map (
            O => \N__16188\,
            I => \M_state_qZ0Z_0\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__16183\,
            I => \M_state_qZ0Z_0\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__16160\,
            I => \N__16157\
        );

    \I__3546\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16154\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__16151\,
            I => \N_414\
        );

    \I__3543\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16143\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__16147\,
            I => \N__16137\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__16146\,
            I => \N__16133\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__16143\,
            I => \N__16130\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16142\,
            I => \N__16125\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16141\,
            I => \N__16125\
        );

    \I__3537\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16122\
        );

    \I__3536\ : InMux
    port map (
            O => \N__16137\,
            I => \N__16114\
        );

    \I__3535\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16114\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16114\
        );

    \I__3533\ : Span4Mux_h
    port map (
            O => \N__16130\,
            I => \N__16107\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16125\,
            I => \N__16107\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16107\
        );

    \I__3530\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16104\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__16114\,
            I => \N__16101\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__16107\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__16104\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__16101\,
            I => this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1
        );

    \I__3525\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16090\
        );

    \I__3524\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16079\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__16090\,
            I => \N__16076\
        );

    \I__3522\ : InMux
    port map (
            O => \N__16089\,
            I => \N__16069\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16088\,
            I => \N__16069\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16069\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16086\,
            I => \N__16062\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16062\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16062\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16083\,
            I => \N__16051\
        );

    \I__3515\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16051\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16079\,
            I => \N__16042\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__16076\,
            I => \N__16042\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16069\,
            I => \N__16042\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__16062\,
            I => \N__16042\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16033\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16033\
        );

    \I__3508\ : InMux
    port map (
            O => \N__16059\,
            I => \N__16033\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16058\,
            I => \N__16033\
        );

    \I__3506\ : InMux
    port map (
            O => \N__16057\,
            I => \N__16028\
        );

    \I__3505\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16028\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16051\,
            I => this_vga_signals_un16_address_if_i1_mux_0
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__16042\,
            I => this_vga_signals_un16_address_if_i1_mux_0
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__16033\,
            I => this_vga_signals_un16_address_if_i1_mux_0
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__16028\,
            I => this_vga_signals_un16_address_if_i1_mux_0
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__16019\,
            I => \N__16016\
        );

    \I__3499\ : CascadeBuf
    port map (
            O => \N__16016\,
            I => \N__16013\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__3497\ : CascadeBuf
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__3495\ : CascadeBuf
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__3493\ : CascadeBuf
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__3491\ : CascadeBuf
    port map (
            O => \N__15992\,
            I => \N__15989\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__3489\ : CascadeBuf
    port map (
            O => \N__15986\,
            I => \N__15983\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__3487\ : CascadeBuf
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__15977\,
            I => \N__15974\
        );

    \I__3485\ : CascadeBuf
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__3483\ : CascadeBuf
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__15965\,
            I => \N__15962\
        );

    \I__3481\ : CascadeBuf
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__15959\,
            I => \N__15956\
        );

    \I__3479\ : CascadeBuf
    port map (
            O => \N__15956\,
            I => \N__15953\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__15953\,
            I => \N__15950\
        );

    \I__3477\ : CascadeBuf
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__3475\ : CascadeBuf
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__15941\,
            I => \N__15938\
        );

    \I__3473\ : CascadeBuf
    port map (
            O => \N__15938\,
            I => \N__15935\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__15935\,
            I => \N__15932\
        );

    \I__3471\ : CascadeBuf
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__3469\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__3467\ : Span12Mux_h
    port map (
            O => \N__15920\,
            I => \N__15916\
        );

    \I__3466\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15913\
        );

    \I__3465\ : Span12Mux_v
    port map (
            O => \N__15916\,
            I => \N__15910\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__15913\,
            I => \M_this_vga_signals_address_10\
        );

    \I__3463\ : Odrv12
    port map (
            O => \N__15910\,
            I => \M_this_vga_signals_address_10\
        );

    \I__3462\ : InMux
    port map (
            O => \N__15905\,
            I => \N__15899\
        );

    \I__3461\ : InMux
    port map (
            O => \N__15904\,
            I => \N__15896\
        );

    \I__3460\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15893\
        );

    \I__3459\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15890\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__15899\,
            I => \N__15887\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__15896\,
            I => \N__15882\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__15893\,
            I => \N__15882\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__15890\,
            I => \N__15876\
        );

    \I__3454\ : Span4Mux_v
    port map (
            O => \N__15887\,
            I => \N__15871\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__15882\,
            I => \N__15871\
        );

    \I__3452\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15866\
        );

    \I__3451\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15866\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__15879\,
            I => \N__15863\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__15876\,
            I => \N__15860\
        );

    \I__3448\ : Sp12to4
    port map (
            O => \N__15871\,
            I => \N__15855\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15855\
        );

    \I__3446\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15852\
        );

    \I__3445\ : Sp12to4
    port map (
            O => \N__15860\,
            I => \N__15845\
        );

    \I__3444\ : Span12Mux_h
    port map (
            O => \N__15855\,
            I => \N__15845\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__15852\,
            I => \N__15845\
        );

    \I__3442\ : Odrv12
    port map (
            O => \N__15845\,
            I => \M_this_vram_read_data_2\
        );

    \I__3441\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15833\
        );

    \I__3440\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15830\
        );

    \I__3439\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15825\
        );

    \I__3438\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15825\
        );

    \I__3437\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15820\
        );

    \I__3436\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15820\
        );

    \I__3435\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15817\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__15833\,
            I => \N__15807\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__15830\,
            I => \N__15807\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__15825\,
            I => \N__15807\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__15820\,
            I => \N__15807\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__15817\,
            I => \N__15804\
        );

    \I__3429\ : InMux
    port map (
            O => \N__15816\,
            I => \N__15801\
        );

    \I__3428\ : Span4Mux_v
    port map (
            O => \N__15807\,
            I => \N__15797\
        );

    \I__3427\ : Span4Mux_v
    port map (
            O => \N__15804\,
            I => \N__15794\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__15801\,
            I => \N__15791\
        );

    \I__3425\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15788\
        );

    \I__3424\ : Sp12to4
    port map (
            O => \N__15797\,
            I => \N__15783\
        );

    \I__3423\ : Sp12to4
    port map (
            O => \N__15794\,
            I => \N__15783\
        );

    \I__3422\ : Span4Mux_v
    port map (
            O => \N__15791\,
            I => \N__15778\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__15788\,
            I => \N__15778\
        );

    \I__3420\ : Odrv12
    port map (
            O => \N__15783\,
            I => this_vram_mem_radreg_11
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__15778\,
            I => this_vram_mem_radreg_11
        );

    \I__3418\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__15770\,
            I => \mem_radreg_RNIMTEJ4_11\
        );

    \I__3416\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__15764\,
            I => m14
        );

    \I__3414\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__15758\,
            I => \rgb_1_cry_0_0_c_RNOZ0\
        );

    \I__3412\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__15752\,
            I => \M_vcounter_q_esr_RNIB9J4TN_9\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__3409\ : InMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__15743\,
            I => \N__15740\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__15740\,
            I => \M_vcounter_q_esr_RNICJRF0D_9\
        );

    \I__3406\ : InMux
    port map (
            O => \N__15737\,
            I => rgb_1_cry_0
        );

    \I__3405\ : InMux
    port map (
            O => \N__15734\,
            I => rgb_1_cry_1
        );

    \I__3404\ : InMux
    port map (
            O => \N__15731\,
            I => rgb_1_cry_2
        );

    \I__3403\ : InMux
    port map (
            O => \N__15728\,
            I => rgb_1_6
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__15725\,
            I => \N_403_cascade_\
        );

    \I__3401\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15719\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15716\
        );

    \I__3399\ : Span4Mux_h
    port map (
            O => \N__15716\,
            I => \N__15713\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__15713\,
            I => \M_current_address_q_RNO_1Z0Z_2\
        );

    \I__3397\ : CascadeMux
    port map (
            O => \N__15710\,
            I => \N__15707\
        );

    \I__3396\ : CascadeBuf
    port map (
            O => \N__15707\,
            I => \N__15704\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__15704\,
            I => \N__15701\
        );

    \I__3394\ : CascadeBuf
    port map (
            O => \N__15701\,
            I => \N__15698\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__3392\ : CascadeBuf
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__15692\,
            I => \N__15689\
        );

    \I__3390\ : CascadeBuf
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__3388\ : CascadeBuf
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__3386\ : CascadeBuf
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__3384\ : CascadeBuf
    port map (
            O => \N__15671\,
            I => \N__15668\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__3382\ : CascadeBuf
    port map (
            O => \N__15665\,
            I => \N__15662\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__15662\,
            I => \N__15659\
        );

    \I__3380\ : CascadeBuf
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__3378\ : CascadeBuf
    port map (
            O => \N__15653\,
            I => \N__15650\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__15650\,
            I => \N__15647\
        );

    \I__3376\ : CascadeBuf
    port map (
            O => \N__15647\,
            I => \N__15644\
        );

    \I__3375\ : CascadeMux
    port map (
            O => \N__15644\,
            I => \N__15641\
        );

    \I__3374\ : CascadeBuf
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__3372\ : CascadeBuf
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__3370\ : CascadeBuf
    port map (
            O => \N__15629\,
            I => \N__15626\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__15626\,
            I => \N__15623\
        );

    \I__3368\ : CascadeBuf
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__15620\,
            I => \N__15616\
        );

    \I__3366\ : InMux
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__3365\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15610\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__15613\,
            I => \N__15607\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__15610\,
            I => \N__15603\
        );

    \I__3362\ : Span4Mux_h
    port map (
            O => \N__15607\,
            I => \N__15600\
        );

    \I__3361\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15597\
        );

    \I__3360\ : Span12Mux_h
    port map (
            O => \N__15603\,
            I => \N__15594\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__15600\,
            I => \M_current_address_qZ0Z_2\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__15597\,
            I => \M_current_address_qZ0Z_2\
        );

    \I__3357\ : Odrv12
    port map (
            O => \N__15594\,
            I => \M_current_address_qZ0Z_2\
        );

    \I__3356\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15584\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__15584\,
            I => \N__15581\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__15581\,
            I => \M_current_address_q_RNO_1Z0Z_13\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__15578\,
            I => \N__15570\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__15577\,
            I => \N__15566\
        );

    \I__3351\ : InMux
    port map (
            O => \N__15576\,
            I => \N__15559\
        );

    \I__3350\ : InMux
    port map (
            O => \N__15575\,
            I => \N__15548\
        );

    \I__3349\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15548\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15548\
        );

    \I__3347\ : InMux
    port map (
            O => \N__15570\,
            I => \N__15541\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15569\,
            I => \N__15541\
        );

    \I__3345\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15541\
        );

    \I__3344\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15538\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15564\,
            I => \N__15531\
        );

    \I__3342\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15531\
        );

    \I__3341\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15531\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__15559\,
            I => \N__15526\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15523\
        );

    \I__3338\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15517\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15556\,
            I => \N__15517\
        );

    \I__3336\ : InMux
    port map (
            O => \N__15555\,
            I => \N__15514\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__15548\,
            I => \N__15511\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15504\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__15538\,
            I => \N__15504\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__15531\,
            I => \N__15504\
        );

    \I__3331\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15501\
        );

    \I__3330\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15498\
        );

    \I__3329\ : Span4Mux_v
    port map (
            O => \N__15526\,
            I => \N__15493\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__15523\,
            I => \N__15493\
        );

    \I__3327\ : InMux
    port map (
            O => \N__15522\,
            I => \N__15490\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__15517\,
            I => \M_state_qZ0Z_1\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__15514\,
            I => \M_state_qZ0Z_1\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__15511\,
            I => \M_state_qZ0Z_1\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__15504\,
            I => \M_state_qZ0Z_1\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__15501\,
            I => \M_state_qZ0Z_1\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__15498\,
            I => \M_state_qZ0Z_1\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__15493\,
            I => \M_state_qZ0Z_1\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__15490\,
            I => \M_state_qZ0Z_1\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__15473\,
            I => \N_407_cascade_\
        );

    \I__3317\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__15467\,
            I => \N__15464\
        );

    \I__3315\ : Span4Mux_h
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__15461\,
            I => \M_current_address_q_RNO_1Z0Z_6\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__3312\ : CascadeBuf
    port map (
            O => \N__15455\,
            I => \N__15452\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__3310\ : CascadeBuf
    port map (
            O => \N__15449\,
            I => \N__15446\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__3308\ : CascadeBuf
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__3306\ : CascadeBuf
    port map (
            O => \N__15437\,
            I => \N__15434\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__3304\ : CascadeBuf
    port map (
            O => \N__15431\,
            I => \N__15428\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__3302\ : CascadeBuf
    port map (
            O => \N__15425\,
            I => \N__15422\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__15422\,
            I => \N__15419\
        );

    \I__3300\ : CascadeBuf
    port map (
            O => \N__15419\,
            I => \N__15416\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__3298\ : CascadeBuf
    port map (
            O => \N__15413\,
            I => \N__15410\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__15410\,
            I => \N__15407\
        );

    \I__3296\ : CascadeBuf
    port map (
            O => \N__15407\,
            I => \N__15404\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__15404\,
            I => \N__15401\
        );

    \I__3294\ : CascadeBuf
    port map (
            O => \N__15401\,
            I => \N__15398\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__15398\,
            I => \N__15395\
        );

    \I__3292\ : CascadeBuf
    port map (
            O => \N__15395\,
            I => \N__15392\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__15392\,
            I => \N__15389\
        );

    \I__3290\ : CascadeBuf
    port map (
            O => \N__15389\,
            I => \N__15386\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__15386\,
            I => \N__15383\
        );

    \I__3288\ : CascadeBuf
    port map (
            O => \N__15383\,
            I => \N__15380\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__3286\ : CascadeBuf
    port map (
            O => \N__15377\,
            I => \N__15374\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \N__15371\
        );

    \I__3284\ : CascadeBuf
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__3282\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15362\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__3280\ : Span4Mux_s2_v
    port map (
            O => \N__15359\,
            I => \N__15355\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15352\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__15355\,
            I => \N__15349\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__15352\,
            I => \N__15346\
        );

    \I__3276\ : Span4Mux_v
    port map (
            O => \N__15349\,
            I => \N__15342\
        );

    \I__3275\ : Span4Mux_h
    port map (
            O => \N__15346\,
            I => \N__15339\
        );

    \I__3274\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15336\
        );

    \I__3273\ : Span4Mux_v
    port map (
            O => \N__15342\,
            I => \N__15333\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__15339\,
            I => \M_current_address_qZ0Z_6\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__15336\,
            I => \M_current_address_qZ0Z_6\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__15333\,
            I => \M_current_address_qZ0Z_6\
        );

    \I__3269\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15316\
        );

    \I__3268\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15316\
        );

    \I__3267\ : SRMux
    port map (
            O => \N__15324\,
            I => \N__15313\
        );

    \I__3266\ : SRMux
    port map (
            O => \N__15323\,
            I => \N__15309\
        );

    \I__3265\ : SRMux
    port map (
            O => \N__15322\,
            I => \N__15303\
        );

    \I__3264\ : SRMux
    port map (
            O => \N__15321\,
            I => \N__15300\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__15316\,
            I => \N__15295\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__15313\,
            I => \N__15295\
        );

    \I__3261\ : SRMux
    port map (
            O => \N__15312\,
            I => \N__15292\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15309\,
            I => \N__15289\
        );

    \I__3259\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15286\
        );

    \I__3258\ : SRMux
    port map (
            O => \N__15307\,
            I => \N__15283\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15280\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15277\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15300\,
            I => \N__15274\
        );

    \I__3254\ : Span4Mux_v
    port map (
            O => \N__15295\,
            I => \N__15271\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__15292\,
            I => \N__15264\
        );

    \I__3252\ : Span4Mux_v
    port map (
            O => \N__15289\,
            I => \N__15264\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__15286\,
            I => \N__15264\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15283\,
            I => \N__15261\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__15280\,
            I => \N__15258\
        );

    \I__3248\ : Span4Mux_h
    port map (
            O => \N__15277\,
            I => \N__15249\
        );

    \I__3247\ : Span4Mux_v
    port map (
            O => \N__15274\,
            I => \N__15249\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__15271\,
            I => \N__15249\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__15264\,
            I => \N__15244\
        );

    \I__3244\ : Span4Mux_h
    port map (
            O => \N__15261\,
            I => \N__15244\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__15258\,
            I => \N__15241\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15257\,
            I => \N__15236\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15236\
        );

    \I__3240\ : Sp12to4
    port map (
            O => \N__15249\,
            I => \N__15227\
        );

    \I__3239\ : Sp12to4
    port map (
            O => \N__15244\,
            I => \N__15227\
        );

    \I__3238\ : Sp12to4
    port map (
            O => \N__15241\,
            I => \N__15227\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15227\
        );

    \I__3236\ : Odrv12
    port map (
            O => \N__15227\,
            I => \M_this_reset_cond_out_0\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__3234\ : CascadeBuf
    port map (
            O => \N__15221\,
            I => \N__15218\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__15218\,
            I => \N__15215\
        );

    \I__3232\ : CascadeBuf
    port map (
            O => \N__15215\,
            I => \N__15212\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__15212\,
            I => \N__15209\
        );

    \I__3230\ : CascadeBuf
    port map (
            O => \N__15209\,
            I => \N__15206\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__3228\ : CascadeBuf
    port map (
            O => \N__15203\,
            I => \N__15200\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__15200\,
            I => \N__15197\
        );

    \I__3226\ : CascadeBuf
    port map (
            O => \N__15197\,
            I => \N__15194\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__15194\,
            I => \N__15191\
        );

    \I__3224\ : CascadeBuf
    port map (
            O => \N__15191\,
            I => \N__15188\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__15188\,
            I => \N__15185\
        );

    \I__3222\ : CascadeBuf
    port map (
            O => \N__15185\,
            I => \N__15182\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__15182\,
            I => \N__15179\
        );

    \I__3220\ : CascadeBuf
    port map (
            O => \N__15179\,
            I => \N__15176\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__3218\ : CascadeBuf
    port map (
            O => \N__15173\,
            I => \N__15170\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__3216\ : CascadeBuf
    port map (
            O => \N__15167\,
            I => \N__15164\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__15164\,
            I => \N__15161\
        );

    \I__3214\ : CascadeBuf
    port map (
            O => \N__15161\,
            I => \N__15158\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__15158\,
            I => \N__15155\
        );

    \I__3212\ : CascadeBuf
    port map (
            O => \N__15155\,
            I => \N__15152\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__15152\,
            I => \N__15149\
        );

    \I__3210\ : CascadeBuf
    port map (
            O => \N__15149\,
            I => \N__15146\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__15146\,
            I => \N__15143\
        );

    \I__3208\ : CascadeBuf
    port map (
            O => \N__15143\,
            I => \N__15140\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__15140\,
            I => \N__15137\
        );

    \I__3206\ : CascadeBuf
    port map (
            O => \N__15137\,
            I => \N__15134\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__15134\,
            I => \N__15131\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15131\,
            I => \N__15128\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__15128\,
            I => \N__15123\
        );

    \I__3202\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15120\
        );

    \I__3201\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15117\
        );

    \I__3200\ : Span12Mux_s9_v
    port map (
            O => \N__15123\,
            I => \N__15114\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__15120\,
            I => \M_current_address_qZ0Z_9\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__15117\,
            I => \M_current_address_qZ0Z_9\
        );

    \I__3197\ : Odrv12
    port map (
            O => \N__15114\,
            I => \M_current_address_qZ0Z_9\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__15107\,
            I => \N__15104\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15101\,
            I => \N_410\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15095\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__15095\,
            I => \N__15092\
        );

    \I__3191\ : Odrv12
    port map (
            O => \N__15092\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__15089\,
            I => \N__15086\
        );

    \I__3189\ : CascadeBuf
    port map (
            O => \N__15086\,
            I => \N__15083\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__15083\,
            I => \N__15080\
        );

    \I__3187\ : CascadeBuf
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__3185\ : CascadeBuf
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__15071\,
            I => \N__15068\
        );

    \I__3183\ : CascadeBuf
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__15065\,
            I => \N__15062\
        );

    \I__3181\ : CascadeBuf
    port map (
            O => \N__15062\,
            I => \N__15059\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__15059\,
            I => \N__15056\
        );

    \I__3179\ : CascadeBuf
    port map (
            O => \N__15056\,
            I => \N__15053\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__15053\,
            I => \N__15050\
        );

    \I__3177\ : CascadeBuf
    port map (
            O => \N__15050\,
            I => \N__15047\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__3175\ : CascadeBuf
    port map (
            O => \N__15044\,
            I => \N__15041\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__15041\,
            I => \N__15038\
        );

    \I__3173\ : CascadeBuf
    port map (
            O => \N__15038\,
            I => \N__15035\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__15035\,
            I => \N__15032\
        );

    \I__3171\ : CascadeBuf
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__15029\,
            I => \N__15026\
        );

    \I__3169\ : CascadeBuf
    port map (
            O => \N__15026\,
            I => \N__15023\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__3167\ : CascadeBuf
    port map (
            O => \N__15020\,
            I => \N__15017\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__3165\ : CascadeBuf
    port map (
            O => \N__15014\,
            I => \N__15011\
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__15011\,
            I => \N__15008\
        );

    \I__3163\ : CascadeBuf
    port map (
            O => \N__15008\,
            I => \N__15005\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__15005\,
            I => \N__15002\
        );

    \I__3161\ : CascadeBuf
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__14999\,
            I => \N__14996\
        );

    \I__3159\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__14993\,
            I => \N__14990\
        );

    \I__3157\ : Span4Mux_h
    port map (
            O => \N__14990\,
            I => \N__14987\
        );

    \I__3156\ : Sp12to4
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__3155\ : Span12Mux_s9_v
    port map (
            O => \N__14984\,
            I => \N__14981\
        );

    \I__3154\ : Odrv12
    port map (
            O => \N__14981\,
            I => \M_this_vga_signals_address_5\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__3152\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14972\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__3150\ : Span4Mux_h
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__14966\,
            I => \mem_radreg_RNIETEJ4_11\
        );

    \I__3148\ : InMux
    port map (
            O => \N__14963\,
            I => \N__14959\
        );

    \I__3147\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14956\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__14959\,
            I => m19
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__14956\,
            I => m19
        );

    \I__3144\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14944\
        );

    \I__3143\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14939\
        );

    \I__3142\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14939\
        );

    \I__3141\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14931\
        );

    \I__3140\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14931\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__14944\,
            I => \N__14926\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__14939\,
            I => \N__14926\
        );

    \I__3137\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14923\
        );

    \I__3136\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14920\
        );

    \I__3135\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14917\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__14931\,
            I => rgb_1_axb_0
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__14926\,
            I => rgb_1_axb_0
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__14923\,
            I => rgb_1_axb_0
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__14920\,
            I => rgb_1_axb_0
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__14917\,
            I => rgb_1_axb_0
        );

    \I__3129\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14901\
        );

    \I__3128\ : InMux
    port map (
            O => \N__14905\,
            I => \N__14898\
        );

    \I__3127\ : InMux
    port map (
            O => \N__14904\,
            I => \N__14895\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__14901\,
            I => \N__14892\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__14898\,
            I => \N__14884\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__14895\,
            I => \N__14884\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__14892\,
            I => \N__14881\
        );

    \I__3122\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14878\
        );

    \I__3121\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14875\
        );

    \I__3120\ : InMux
    port map (
            O => \N__14889\,
            I => \N__14872\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__14884\,
            I => a0_b_0
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__14881\,
            I => a0_b_0
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__14878\,
            I => a0_b_0
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__14875\,
            I => a0_b_0
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__14872\,
            I => a0_b_0
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__14861\,
            I => \m46_am_cascade_\
        );

    \I__3113\ : InMux
    port map (
            O => \N__14858\,
            I => \N__14855\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__14852\,
            I => m46_bm
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__14849\,
            I => \N__14846\
        );

    \I__3109\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__14843\,
            I => \N__14840\
        );

    \I__3107\ : Span12Mux_h
    port map (
            O => \N__14840\,
            I => \N__14837\
        );

    \I__3106\ : Odrv12
    port map (
            O => \N__14837\,
            I => rgb_2_5
        );

    \I__3105\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14831\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N_352\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__14828\,
            I => \N_408_cascade_\
        );

    \I__3102\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__14819\,
            I => \M_current_address_q_RNO_1Z0Z_7\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__3098\ : CascadeBuf
    port map (
            O => \N__14813\,
            I => \N__14810\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__3096\ : CascadeBuf
    port map (
            O => \N__14807\,
            I => \N__14804\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__3094\ : CascadeBuf
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__14798\,
            I => \N__14795\
        );

    \I__3092\ : CascadeBuf
    port map (
            O => \N__14795\,
            I => \N__14792\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__14792\,
            I => \N__14789\
        );

    \I__3090\ : CascadeBuf
    port map (
            O => \N__14789\,
            I => \N__14786\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__3088\ : CascadeBuf
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__14780\,
            I => \N__14777\
        );

    \I__3086\ : CascadeBuf
    port map (
            O => \N__14777\,
            I => \N__14774\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__3084\ : CascadeBuf
    port map (
            O => \N__14771\,
            I => \N__14768\
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__14768\,
            I => \N__14765\
        );

    \I__3082\ : CascadeBuf
    port map (
            O => \N__14765\,
            I => \N__14762\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__3080\ : CascadeBuf
    port map (
            O => \N__14759\,
            I => \N__14756\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__3078\ : CascadeBuf
    port map (
            O => \N__14753\,
            I => \N__14750\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__3076\ : CascadeBuf
    port map (
            O => \N__14747\,
            I => \N__14744\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__3074\ : CascadeBuf
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__14738\,
            I => \N__14735\
        );

    \I__3072\ : CascadeBuf
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__14732\,
            I => \N__14729\
        );

    \I__3070\ : CascadeBuf
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \N__14723\
        );

    \I__3068\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14720\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__14717\,
            I => \N__14713\
        );

    \I__3065\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14709\
        );

    \I__3064\ : Sp12to4
    port map (
            O => \N__14713\,
            I => \N__14706\
        );

    \I__3063\ : InMux
    port map (
            O => \N__14712\,
            I => \N__14703\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N__14698\
        );

    \I__3061\ : Span12Mux_s11_v
    port map (
            O => \N__14706\,
            I => \N__14698\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__14703\,
            I => \M_current_address_qZ0Z_7\
        );

    \I__3059\ : Odrv12
    port map (
            O => \N__14698\,
            I => \M_current_address_qZ0Z_7\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__3057\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14687\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__14687\,
            I => \N_405\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__3053\ : Odrv4
    port map (
            O => \N__14678\,
            I => \M_current_address_q_RNO_1Z0Z_4\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__3051\ : CascadeBuf
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__3049\ : CascadeBuf
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__3047\ : CascadeBuf
    port map (
            O => \N__14660\,
            I => \N__14657\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__3045\ : CascadeBuf
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__3043\ : CascadeBuf
    port map (
            O => \N__14648\,
            I => \N__14645\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__3041\ : CascadeBuf
    port map (
            O => \N__14642\,
            I => \N__14639\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__14639\,
            I => \N__14636\
        );

    \I__3039\ : CascadeBuf
    port map (
            O => \N__14636\,
            I => \N__14633\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__14633\,
            I => \N__14630\
        );

    \I__3037\ : CascadeBuf
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__3035\ : CascadeBuf
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__3033\ : CascadeBuf
    port map (
            O => \N__14618\,
            I => \N__14615\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__3031\ : CascadeBuf
    port map (
            O => \N__14612\,
            I => \N__14609\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__14609\,
            I => \N__14606\
        );

    \I__3029\ : CascadeBuf
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__3027\ : CascadeBuf
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__3025\ : CascadeBuf
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__14591\,
            I => \N__14588\
        );

    \I__3023\ : CascadeBuf
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__14585\,
            I => \N__14582\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14579\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__14579\,
            I => \N__14576\
        );

    \I__3019\ : Span4Mux_s1_v
    port map (
            O => \N__14576\,
            I => \N__14572\
        );

    \I__3018\ : InMux
    port map (
            O => \N__14575\,
            I => \N__14569\
        );

    \I__3017\ : Sp12to4
    port map (
            O => \N__14572\,
            I => \N__14565\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__14569\,
            I => \N__14562\
        );

    \I__3015\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14559\
        );

    \I__3014\ : Span12Mux_h
    port map (
            O => \N__14565\,
            I => \N__14556\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__14562\,
            I => \M_current_address_qZ0Z_4\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__14559\,
            I => \M_current_address_qZ0Z_4\
        );

    \I__3011\ : Odrv12
    port map (
            O => \N__14556\,
            I => \M_current_address_qZ0Z_4\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__3009\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14542\
        );

    \I__3008\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14539\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__14542\,
            I => \N__14536\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__14536\,
            I => \N__14530\
        );

    \I__3004\ : Span4Mux_h
    port map (
            O => \N__14533\,
            I => \N__14527\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__14530\,
            I => \M_state_q_ns_0_a3_0_2_0\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__14527\,
            I => \M_state_q_ns_0_a3_0_2_0\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__14522\,
            I => \N__14519\
        );

    \I__3000\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N_351\
        );

    \I__2998\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14509\
        );

    \I__2997\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14506\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__14509\,
            I => m24
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__14506\,
            I => m24
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__14501\,
            I => \m40_cascade_\
        );

    \I__2993\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__14495\,
            I => m41
        );

    \I__2991\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14486\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14486\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__14486\,
            I => m10
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__14483\,
            I => \rgb_1_axb_0_cascade_\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14480\,
            I => \N__14474\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14474\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__14474\,
            I => \N__14471\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__14471\,
            I => \N__14468\
        );

    \I__2983\ : Odrv4
    port map (
            O => \N__14468\,
            I => m15
        );

    \I__2982\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14458\
        );

    \I__2980\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14455\
        );

    \I__2979\ : Span4Mux_v
    port map (
            O => \N__14458\,
            I => \N__14450\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__14455\,
            I => \N__14450\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__14450\,
            I => rgb_1_0
        );

    \I__2976\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14444\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__14444\,
            I => m37
        );

    \I__2974\ : SRMux
    port map (
            O => \N__14441\,
            I => \N__14437\
        );

    \I__2973\ : SRMux
    port map (
            O => \N__14440\,
            I => \N__14431\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14427\
        );

    \I__2971\ : SRMux
    port map (
            O => \N__14436\,
            I => \N__14423\
        );

    \I__2970\ : SRMux
    port map (
            O => \N__14435\,
            I => \N__14420\
        );

    \I__2969\ : SRMux
    port map (
            O => \N__14434\,
            I => \N__14415\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__14431\,
            I => \N__14409\
        );

    \I__2967\ : SRMux
    port map (
            O => \N__14430\,
            I => \N__14406\
        );

    \I__2966\ : Span4Mux_s3_v
    port map (
            O => \N__14427\,
            I => \N__14403\
        );

    \I__2965\ : SRMux
    port map (
            O => \N__14426\,
            I => \N__14400\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__14423\,
            I => \N__14393\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14420\,
            I => \N__14393\
        );

    \I__2962\ : SRMux
    port map (
            O => \N__14419\,
            I => \N__14390\
        );

    \I__2961\ : SRMux
    port map (
            O => \N__14418\,
            I => \N__14382\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__14415\,
            I => \N__14379\
        );

    \I__2959\ : SRMux
    port map (
            O => \N__14414\,
            I => \N__14376\
        );

    \I__2958\ : SRMux
    port map (
            O => \N__14413\,
            I => \N__14373\
        );

    \I__2957\ : SRMux
    port map (
            O => \N__14412\,
            I => \N__14370\
        );

    \I__2956\ : Span4Mux_h
    port map (
            O => \N__14409\,
            I => \N__14363\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__14406\,
            I => \N__14363\
        );

    \I__2954\ : Span4Mux_v
    port map (
            O => \N__14403\,
            I => \N__14358\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__14400\,
            I => \N__14358\
        );

    \I__2952\ : SRMux
    port map (
            O => \N__14399\,
            I => \N__14355\
        );

    \I__2951\ : SRMux
    port map (
            O => \N__14398\,
            I => \N__14352\
        );

    \I__2950\ : Span4Mux_s3_v
    port map (
            O => \N__14393\,
            I => \N__14346\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__14390\,
            I => \N__14346\
        );

    \I__2948\ : SRMux
    port map (
            O => \N__14389\,
            I => \N__14343\
        );

    \I__2947\ : SRMux
    port map (
            O => \N__14388\,
            I => \N__14340\
        );

    \I__2946\ : IoInMux
    port map (
            O => \N__14387\,
            I => \N__14334\
        );

    \I__2945\ : SRMux
    port map (
            O => \N__14386\,
            I => \N__14331\
        );

    \I__2944\ : SRMux
    port map (
            O => \N__14385\,
            I => \N__14328\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__14382\,
            I => \N__14320\
        );

    \I__2942\ : Span4Mux_h
    port map (
            O => \N__14379\,
            I => \N__14320\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__14376\,
            I => \N__14320\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__14373\,
            I => \N__14315\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__14370\,
            I => \N__14315\
        );

    \I__2938\ : SRMux
    port map (
            O => \N__14369\,
            I => \N__14312\
        );

    \I__2937\ : SRMux
    port map (
            O => \N__14368\,
            I => \N__14308\
        );

    \I__2936\ : Span4Mux_v
    port map (
            O => \N__14363\,
            I => \N__14298\
        );

    \I__2935\ : Span4Mux_h
    port map (
            O => \N__14358\,
            I => \N__14298\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__14355\,
            I => \N__14298\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__14352\,
            I => \N__14295\
        );

    \I__2932\ : SRMux
    port map (
            O => \N__14351\,
            I => \N__14292\
        );

    \I__2931\ : Span4Mux_v
    port map (
            O => \N__14346\,
            I => \N__14285\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14343\,
            I => \N__14285\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14340\,
            I => \N__14285\
        );

    \I__2928\ : SRMux
    port map (
            O => \N__14339\,
            I => \N__14282\
        );

    \I__2927\ : SRMux
    port map (
            O => \N__14338\,
            I => \N__14279\
        );

    \I__2926\ : InMux
    port map (
            O => \N__14337\,
            I => \N__14275\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__14334\,
            I => \N__14272\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14331\,
            I => \N__14266\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14328\,
            I => \N__14266\
        );

    \I__2922\ : SRMux
    port map (
            O => \N__14327\,
            I => \N__14263\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__14320\,
            I => \N__14256\
        );

    \I__2920\ : Span4Mux_v
    port map (
            O => \N__14315\,
            I => \N__14256\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__14312\,
            I => \N__14256\
        );

    \I__2918\ : SRMux
    port map (
            O => \N__14311\,
            I => \N__14253\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__14308\,
            I => \N__14250\
        );

    \I__2916\ : SRMux
    port map (
            O => \N__14307\,
            I => \N__14247\
        );

    \I__2915\ : SRMux
    port map (
            O => \N__14306\,
            I => \N__14244\
        );

    \I__2914\ : SRMux
    port map (
            O => \N__14305\,
            I => \N__14241\
        );

    \I__2913\ : Span4Mux_v
    port map (
            O => \N__14298\,
            I => \N__14234\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__14295\,
            I => \N__14234\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__14292\,
            I => \N__14234\
        );

    \I__2910\ : Span4Mux_v
    port map (
            O => \N__14285\,
            I => \N__14227\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__14282\,
            I => \N__14227\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__14279\,
            I => \N__14227\
        );

    \I__2907\ : SRMux
    port map (
            O => \N__14278\,
            I => \N__14224\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__14275\,
            I => \N__14220\
        );

    \I__2905\ : Span4Mux_s2_h
    port map (
            O => \N__14272\,
            I => \N__14217\
        );

    \I__2904\ : SRMux
    port map (
            O => \N__14271\,
            I => \N__14214\
        );

    \I__2903\ : Span4Mux_v
    port map (
            O => \N__14266\,
            I => \N__14209\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14209\
        );

    \I__2901\ : Span4Mux_v
    port map (
            O => \N__14256\,
            I => \N__14204\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__14253\,
            I => \N__14204\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__14250\,
            I => \N__14199\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__14247\,
            I => \N__14199\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__14244\,
            I => \N__14194\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14194\
        );

    \I__2895\ : Span4Mux_v
    port map (
            O => \N__14234\,
            I => \N__14187\
        );

    \I__2894\ : Span4Mux_v
    port map (
            O => \N__14227\,
            I => \N__14187\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14187\
        );

    \I__2892\ : SRMux
    port map (
            O => \N__14223\,
            I => \N__14184\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__14220\,
            I => \N__14179\
        );

    \I__2890\ : Sp12to4
    port map (
            O => \N__14217\,
            I => \N__14176\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__14214\,
            I => \N__14173\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__14209\,
            I => \N__14169\
        );

    \I__2887\ : Span4Mux_v
    port map (
            O => \N__14204\,
            I => \N__14164\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__14199\,
            I => \N__14164\
        );

    \I__2885\ : Span4Mux_v
    port map (
            O => \N__14194\,
            I => \N__14157\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__14187\,
            I => \N__14157\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14184\,
            I => \N__14157\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__14183\,
            I => \N__14154\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__14182\,
            I => \N__14151\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__14179\,
            I => \N__14147\
        );

    \I__2879\ : Span12Mux_v
    port map (
            O => \N__14176\,
            I => \N__14144\
        );

    \I__2878\ : Span12Mux_h
    port map (
            O => \N__14173\,
            I => \N__14141\
        );

    \I__2877\ : SRMux
    port map (
            O => \N__14172\,
            I => \N__14138\
        );

    \I__2876\ : Span4Mux_v
    port map (
            O => \N__14169\,
            I => \N__14131\
        );

    \I__2875\ : Span4Mux_h
    port map (
            O => \N__14164\,
            I => \N__14131\
        );

    \I__2874\ : Span4Mux_h
    port map (
            O => \N__14157\,
            I => \N__14131\
        );

    \I__2873\ : InMux
    port map (
            O => \N__14154\,
            I => \N__14128\
        );

    \I__2872\ : InMux
    port map (
            O => \N__14151\,
            I => \N__14123\
        );

    \I__2871\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14123\
        );

    \I__2870\ : Span4Mux_v
    port map (
            O => \N__14147\,
            I => \N__14120\
        );

    \I__2869\ : Span12Mux_h
    port map (
            O => \N__14144\,
            I => \N__14113\
        );

    \I__2868\ : Span12Mux_v
    port map (
            O => \N__14141\,
            I => \N__14113\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__14138\,
            I => \N__14113\
        );

    \I__2866\ : Span4Mux_h
    port map (
            O => \N__14131\,
            I => \N__14110\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__14128\,
            I => \N__14105\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__14123\,
            I => \N__14105\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__14120\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2862\ : Odrv12
    port map (
            O => \N__14113\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__14110\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__14105\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14096\,
            I => rgb291
        );

    \I__2858\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14085\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14085\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14081\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14078\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__14085\,
            I => \N__14074\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14071\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14081\,
            I => \N__14068\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14078\,
            I => \N__14065\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14062\
        );

    \I__2849\ : Span4Mux_h
    port map (
            O => \N__14074\,
            I => \N__14057\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__14071\,
            I => \N__14057\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__14068\,
            I => \N__14054\
        );

    \I__2846\ : Span4Mux_v
    port map (
            O => \N__14065\,
            I => \N__14049\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__14062\,
            I => \N__14049\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__14057\,
            I => \N__14046\
        );

    \I__2843\ : Sp12to4
    port map (
            O => \N__14054\,
            I => \N__14043\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__14049\,
            I => \N__14040\
        );

    \I__2841\ : Sp12to4
    port map (
            O => \N__14046\,
            I => \N__14037\
        );

    \I__2840\ : Span12Mux_h
    port map (
            O => \N__14043\,
            I => \N__14034\
        );

    \I__2839\ : Span4Mux_h
    port map (
            O => \N__14040\,
            I => \N__14031\
        );

    \I__2838\ : Odrv12
    port map (
            O => \N__14037\,
            I => \this_vga_signals.rgb_1_sqmuxa\
        );

    \I__2837\ : Odrv12
    port map (
            O => \N__14034\,
            I => \this_vga_signals.rgb_1_sqmuxa\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__14031\,
            I => \this_vga_signals.rgb_1_sqmuxa\
        );

    \I__2835\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__14021\,
            I => \mem_radreg_RNIMTEJ4_0_11\
        );

    \I__2833\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__14015\,
            I => \mem_radreg_RNIETEJ4_0_11\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__14012\,
            I => \m44_cascade_\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__14009\,
            I => \m22_am_cascade_\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__14003\,
            I => \N__14000\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__14000\,
            I => m22_ns
        );

    \I__2826\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__13994\,
            I => m22_bm
        );

    \I__2824\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13988\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__13988\,
            I => \M_current_address_q_RNO_1Z0Z_8\
        );

    \I__2822\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2820\ : Span4Mux_h
    port map (
            O => \N__13979\,
            I => \N__13976\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__13976\,
            I => \N_409\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__2817\ : CascadeBuf
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__13967\,
            I => \N__13964\
        );

    \I__2815\ : CascadeBuf
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__2813\ : CascadeBuf
    port map (
            O => \N__13958\,
            I => \N__13955\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__2811\ : CascadeBuf
    port map (
            O => \N__13952\,
            I => \N__13949\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__13949\,
            I => \N__13946\
        );

    \I__2809\ : CascadeBuf
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__2807\ : CascadeBuf
    port map (
            O => \N__13940\,
            I => \N__13937\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__2805\ : CascadeBuf
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__2803\ : CascadeBuf
    port map (
            O => \N__13928\,
            I => \N__13925\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__13925\,
            I => \N__13922\
        );

    \I__2801\ : CascadeBuf
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__2799\ : CascadeBuf
    port map (
            O => \N__13916\,
            I => \N__13913\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__13913\,
            I => \N__13910\
        );

    \I__2797\ : CascadeBuf
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__13907\,
            I => \N__13904\
        );

    \I__2795\ : CascadeBuf
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__2793\ : CascadeBuf
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2791\ : CascadeBuf
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__13889\,
            I => \N__13886\
        );

    \I__2789\ : CascadeBuf
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__2787\ : InMux
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__2785\ : Span4Mux_s3_v
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__2784\ : Span4Mux_h
    port map (
            O => \N__13871\,
            I => \N__13867\
        );

    \I__2783\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13863\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__13867\,
            I => \N__13860\
        );

    \I__2781\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13857\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__13863\,
            I => \N__13854\
        );

    \I__2779\ : Span4Mux_v
    port map (
            O => \N__13860\,
            I => \N__13851\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__13857\,
            I => \M_current_address_qZ0Z_8\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__13854\,
            I => \M_current_address_qZ0Z_8\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__13851\,
            I => \M_current_address_qZ0Z_8\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13844\,
            I => \N__13841\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__2773\ : Odrv12
    port map (
            O => \N__13838\,
            I => \N_412\
        );

    \I__2772\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13832\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__13832\,
            I => \M_current_address_q_RNO_1Z0Z_11\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__13829\,
            I => \N__13825\
        );

    \I__2769\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__2768\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13819\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__13822\,
            I => \N__13814\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__13819\,
            I => \N__13814\
        );

    \I__2765\ : Span4Mux_v
    port map (
            O => \N__13814\,
            I => \N__13811\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__13811\,
            I => \N__13808\
        );

    \I__2763\ : Sp12to4
    port map (
            O => \N__13808\,
            I => \N__13805\
        );

    \I__2762\ : Span12Mux_h
    port map (
            O => \N__13805\,
            I => \N__13802\
        );

    \I__2761\ : Odrv12
    port map (
            O => \N__13802\,
            I => port_data_c_4
        );

    \I__2760\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13796\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__13796\,
            I => \M_current_address_q_RNO_1Z0Z_9\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__13793\,
            I => \N__13789\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__13792\,
            I => \N__13784\
        );

    \I__2756\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13779\
        );

    \I__2755\ : InMux
    port map (
            O => \N__13788\,
            I => \N__13779\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__13787\,
            I => \N__13776\
        );

    \I__2753\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13771\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__13779\,
            I => \N__13766\
        );

    \I__2751\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13761\
        );

    \I__2750\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13761\
        );

    \I__2749\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13758\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__13771\,
            I => \N__13755\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__13770\,
            I => \N__13752\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__13769\,
            I => \N__13747\
        );

    \I__2745\ : Span4Mux_v
    port map (
            O => \N__13766\,
            I => \N__13742\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__13761\,
            I => \N__13742\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__13758\,
            I => \N__13739\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__13755\,
            I => \N__13736\
        );

    \I__2741\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13731\
        );

    \I__2740\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13731\
        );

    \I__2739\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13726\
        );

    \I__2738\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13726\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__13742\,
            I => \N__13721\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__13739\,
            I => \N__13721\
        );

    \I__2735\ : Span4Mux_h
    port map (
            O => \N__13736\,
            I => \N__13714\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__13731\,
            I => \N__13714\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__13726\,
            I => \N__13714\
        );

    \I__2732\ : Span4Mux_h
    port map (
            O => \N__13721\,
            I => \N__13711\
        );

    \I__2731\ : Span4Mux_v
    port map (
            O => \N__13714\,
            I => \N__13708\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__13711\,
            I => \N__13705\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__13708\,
            I => \N__13702\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__13705\,
            I => \M_this_vram_read_data_1\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__13702\,
            I => \M_this_vram_read_data_1\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__13697\,
            I => \N__13693\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__13696\,
            I => \N__13690\
        );

    \I__2724\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13687\
        );

    \I__2723\ : InMux
    port map (
            O => \N__13690\,
            I => \N__13684\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__13687\,
            I => \N__13681\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__13684\,
            I => \N__13678\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__13681\,
            I => \N__13673\
        );

    \I__2719\ : Span4Mux_v
    port map (
            O => \N__13678\,
            I => \N__13673\
        );

    \I__2718\ : Sp12to4
    port map (
            O => \N__13673\,
            I => \N__13670\
        );

    \I__2717\ : Span12Mux_h
    port map (
            O => \N__13670\,
            I => \N__13667\
        );

    \I__2716\ : Odrv12
    port map (
            O => \N__13667\,
            I => port_data_c_5
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__13664\,
            I => \N_413_cascade_\
        );

    \I__2714\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13658\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__13658\,
            I => \M_current_address_q_RNO_1Z0Z_12\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__13655\,
            I => \N__13652\
        );

    \I__2711\ : InMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__13649\,
            I => \N_411\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13646\,
            I => \N__13643\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__13643\,
            I => \M_current_address_q_RNO_1Z0Z_10\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__2706\ : CascadeBuf
    port map (
            O => \N__13637\,
            I => \N__13634\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__13634\,
            I => \N__13631\
        );

    \I__2704\ : CascadeBuf
    port map (
            O => \N__13631\,
            I => \N__13628\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__13628\,
            I => \N__13625\
        );

    \I__2702\ : CascadeBuf
    port map (
            O => \N__13625\,
            I => \N__13622\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__13622\,
            I => \N__13619\
        );

    \I__2700\ : CascadeBuf
    port map (
            O => \N__13619\,
            I => \N__13616\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__2698\ : CascadeBuf
    port map (
            O => \N__13613\,
            I => \N__13610\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__13610\,
            I => \N__13607\
        );

    \I__2696\ : CascadeBuf
    port map (
            O => \N__13607\,
            I => \N__13604\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__13604\,
            I => \N__13601\
        );

    \I__2694\ : CascadeBuf
    port map (
            O => \N__13601\,
            I => \N__13598\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__13598\,
            I => \N__13595\
        );

    \I__2692\ : CascadeBuf
    port map (
            O => \N__13595\,
            I => \N__13592\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__13592\,
            I => \N__13589\
        );

    \I__2690\ : CascadeBuf
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__13586\,
            I => \N__13583\
        );

    \I__2688\ : CascadeBuf
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__13580\,
            I => \N__13577\
        );

    \I__2686\ : CascadeBuf
    port map (
            O => \N__13577\,
            I => \N__13574\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__13574\,
            I => \N__13571\
        );

    \I__2684\ : CascadeBuf
    port map (
            O => \N__13571\,
            I => \N__13568\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__13568\,
            I => \N__13565\
        );

    \I__2682\ : CascadeBuf
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2680\ : CascadeBuf
    port map (
            O => \N__13559\,
            I => \N__13556\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__13556\,
            I => \N__13553\
        );

    \I__2678\ : CascadeBuf
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__13550\,
            I => \N__13547\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13544\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__13544\,
            I => \N__13539\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13536\
        );

    \I__2673\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13533\
        );

    \I__2672\ : Span12Mux_h
    port map (
            O => \N__13539\,
            I => \N__13530\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__13536\,
            I => \M_current_address_qZ0Z_10\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__13533\,
            I => \M_current_address_qZ0Z_10\
        );

    \I__2669\ : Odrv12
    port map (
            O => \N__13530\,
            I => \M_current_address_qZ0Z_10\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__13523\,
            I => \N__13520\
        );

    \I__2667\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13517\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__13517\,
            I => \N_404\
        );

    \I__2665\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13511\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__13511\,
            I => \M_current_address_q_RNO_1Z0Z_3\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__2662\ : CascadeBuf
    port map (
            O => \N__13505\,
            I => \N__13502\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__13502\,
            I => \N__13499\
        );

    \I__2660\ : CascadeBuf
    port map (
            O => \N__13499\,
            I => \N__13496\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__13496\,
            I => \N__13493\
        );

    \I__2658\ : CascadeBuf
    port map (
            O => \N__13493\,
            I => \N__13490\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__2656\ : CascadeBuf
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__13484\,
            I => \N__13481\
        );

    \I__2654\ : CascadeBuf
    port map (
            O => \N__13481\,
            I => \N__13478\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2652\ : CascadeBuf
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__2650\ : CascadeBuf
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__2648\ : CascadeBuf
    port map (
            O => \N__13463\,
            I => \N__13460\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__13460\,
            I => \N__13457\
        );

    \I__2646\ : CascadeBuf
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__2644\ : CascadeBuf
    port map (
            O => \N__13451\,
            I => \N__13448\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__2642\ : CascadeBuf
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__13442\,
            I => \N__13439\
        );

    \I__2640\ : CascadeBuf
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2638\ : CascadeBuf
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2636\ : CascadeBuf
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__13424\,
            I => \N__13421\
        );

    \I__2634\ : CascadeBuf
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__13418\,
            I => \N__13415\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13412\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__13412\,
            I => \N__13409\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__13409\,
            I => \N__13404\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__13408\,
            I => \N__13401\
        );

    \I__2628\ : InMux
    port map (
            O => \N__13407\,
            I => \N__13398\
        );

    \I__2627\ : Sp12to4
    port map (
            O => \N__13404\,
            I => \N__13395\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13392\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__13398\,
            I => \N__13387\
        );

    \I__2624\ : Span12Mux_s11_v
    port map (
            O => \N__13395\,
            I => \N__13387\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__13392\,
            I => \M_current_address_qZ0Z_3\
        );

    \I__2622\ : Odrv12
    port map (
            O => \N__13387\,
            I => \M_current_address_qZ0Z_3\
        );

    \I__2621\ : InMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__13379\,
            I => \M_current_address_q_RNO_1Z0Z_5\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__2618\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13370\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__13370\,
            I => \N_406\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__13367\,
            I => \N__13364\
        );

    \I__2615\ : CascadeBuf
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__13361\,
            I => \N__13358\
        );

    \I__2613\ : CascadeBuf
    port map (
            O => \N__13358\,
            I => \N__13355\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__13355\,
            I => \N__13352\
        );

    \I__2611\ : CascadeBuf
    port map (
            O => \N__13352\,
            I => \N__13349\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__13349\,
            I => \N__13346\
        );

    \I__2609\ : CascadeBuf
    port map (
            O => \N__13346\,
            I => \N__13343\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__13343\,
            I => \N__13340\
        );

    \I__2607\ : CascadeBuf
    port map (
            O => \N__13340\,
            I => \N__13337\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__13337\,
            I => \N__13334\
        );

    \I__2605\ : CascadeBuf
    port map (
            O => \N__13334\,
            I => \N__13331\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__2603\ : CascadeBuf
    port map (
            O => \N__13328\,
            I => \N__13325\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__13325\,
            I => \N__13322\
        );

    \I__2601\ : CascadeBuf
    port map (
            O => \N__13322\,
            I => \N__13319\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__13319\,
            I => \N__13316\
        );

    \I__2599\ : CascadeBuf
    port map (
            O => \N__13316\,
            I => \N__13313\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__13313\,
            I => \N__13310\
        );

    \I__2597\ : CascadeBuf
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__13307\,
            I => \N__13304\
        );

    \I__2595\ : CascadeBuf
    port map (
            O => \N__13304\,
            I => \N__13301\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__13301\,
            I => \N__13298\
        );

    \I__2593\ : CascadeBuf
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__13295\,
            I => \N__13292\
        );

    \I__2591\ : CascadeBuf
    port map (
            O => \N__13292\,
            I => \N__13289\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__2589\ : CascadeBuf
    port map (
            O => \N__13286\,
            I => \N__13283\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__13283\,
            I => \N__13280\
        );

    \I__2587\ : CascadeBuf
    port map (
            O => \N__13280\,
            I => \N__13277\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__2585\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13271\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__13271\,
            I => \N__13266\
        );

    \I__2583\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13263\
        );

    \I__2582\ : InMux
    port map (
            O => \N__13269\,
            I => \N__13260\
        );

    \I__2581\ : Span12Mux_s11_v
    port map (
            O => \N__13266\,
            I => \N__13257\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__13263\,
            I => \M_current_address_qZ0Z_5\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13260\,
            I => \M_current_address_qZ0Z_5\
        );

    \I__2578\ : Odrv12
    port map (
            O => \N__13257\,
            I => \M_current_address_qZ0Z_5\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__13250\,
            I => \N_402_cascade_\
        );

    \I__2576\ : InMux
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__13244\,
            I => \M_current_address_q_RNO_1Z0Z_1\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__13241\,
            I => \N__13238\
        );

    \I__2573\ : CascadeBuf
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__2571\ : CascadeBuf
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2569\ : CascadeBuf
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__2567\ : CascadeBuf
    port map (
            O => \N__13220\,
            I => \N__13217\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__13217\,
            I => \N__13214\
        );

    \I__2565\ : CascadeBuf
    port map (
            O => \N__13214\,
            I => \N__13211\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__13211\,
            I => \N__13208\
        );

    \I__2563\ : CascadeBuf
    port map (
            O => \N__13208\,
            I => \N__13205\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__13205\,
            I => \N__13202\
        );

    \I__2561\ : CascadeBuf
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__13199\,
            I => \N__13196\
        );

    \I__2559\ : CascadeBuf
    port map (
            O => \N__13196\,
            I => \N__13193\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__2557\ : CascadeBuf
    port map (
            O => \N__13190\,
            I => \N__13187\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \N__13184\
        );

    \I__2555\ : CascadeBuf
    port map (
            O => \N__13184\,
            I => \N__13181\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__13181\,
            I => \N__13178\
        );

    \I__2553\ : CascadeBuf
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__13175\,
            I => \N__13172\
        );

    \I__2551\ : CascadeBuf
    port map (
            O => \N__13172\,
            I => \N__13169\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__13169\,
            I => \N__13166\
        );

    \I__2549\ : CascadeBuf
    port map (
            O => \N__13166\,
            I => \N__13163\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__13163\,
            I => \N__13160\
        );

    \I__2547\ : CascadeBuf
    port map (
            O => \N__13160\,
            I => \N__13157\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__13157\,
            I => \N__13154\
        );

    \I__2545\ : CascadeBuf
    port map (
            O => \N__13154\,
            I => \N__13151\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__13151\,
            I => \N__13148\
        );

    \I__2543\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__13145\,
            I => \N__13142\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__13142\,
            I => \N__13139\
        );

    \I__2540\ : Span4Mux_h
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__2539\ : Span4Mux_h
    port map (
            O => \N__13136\,
            I => \N__13131\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13135\,
            I => \N__13128\
        );

    \I__2537\ : InMux
    port map (
            O => \N__13134\,
            I => \N__13125\
        );

    \I__2536\ : Span4Mux_v
    port map (
            O => \N__13131\,
            I => \N__13122\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__13128\,
            I => \M_current_address_qZ0Z_1\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__13125\,
            I => \M_current_address_qZ0Z_1\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__13122\,
            I => \M_current_address_qZ0Z_1\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__13115\,
            I => \m32_am_cascade_\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13109\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__13109\,
            I => m7_bm
        );

    \I__2529\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13103\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13103\,
            I => m32_bm
        );

    \I__2527\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13096\
        );

    \I__2526\ : InMux
    port map (
            O => \N__13099\,
            I => \N__13093\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__13096\,
            I => \N__13090\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__13093\,
            I => \N__13087\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__13090\,
            I => m32_ns
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__13087\,
            I => m32_ns
        );

    \I__2521\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13079\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13079\,
            I => \N__13076\
        );

    \I__2519\ : Span4Mux_h
    port map (
            O => \N__13076\,
            I => \N__13073\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__13073\,
            I => rgb_2_4
        );

    \I__2517\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13067\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13067\,
            I => \N__13063\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13060\
        );

    \I__2514\ : Odrv12
    port map (
            O => \N__13063\,
            I => m29
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__13060\,
            I => m29
        );

    \I__2512\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13052\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13049\
        );

    \I__2510\ : Span12Mux_h
    port map (
            O => \N__13049\,
            I => \N__13046\
        );

    \I__2509\ : Odrv12
    port map (
            O => \N__13046\,
            I => \this_vga_signals.rgb_bmZ0Z_3\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13043\,
            I => \un1_M_current_address_q_cry_12\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13033\
        );

    \I__2506\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13033\
        );

    \I__2505\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13029\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13033\,
            I => \N__13026\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13032\,
            I => \N__13023\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__13029\,
            I => \N__13020\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__13026\,
            I => \N__13017\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13023\,
            I => \this_pixel_clock.M_counter_qZ0Z_0\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__13020\,
            I => \this_pixel_clock.M_counter_qZ0Z_0\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__13017\,
            I => \this_pixel_clock.M_counter_qZ0Z_0\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__13010\,
            I => \N__13003\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13009\,
            I => \N__12998\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13008\,
            I => \N__12998\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13007\,
            I => \N__12995\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13006\,
            I => \N__12992\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13003\,
            I => \N__12989\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__12998\,
            I => \N__12981\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__12995\,
            I => \N__12981\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12992\,
            I => \N__12976\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__12989\,
            I => \N__12976\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__12988\,
            I => \N__12973\
        );

    \I__2486\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12968\
        );

    \I__2485\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12968\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__12981\,
            I => \N__12963\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__12976\,
            I => \N__12963\
        );

    \I__2482\ : InMux
    port map (
            O => \N__12973\,
            I => \N__12960\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__12968\,
            I => \N__12955\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__12963\,
            I => \N__12952\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__12960\,
            I => \N__12949\
        );

    \I__2478\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12946\
        );

    \I__2477\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12943\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__12955\,
            I => \N__12940\
        );

    \I__2475\ : Sp12to4
    port map (
            O => \N__12952\,
            I => \N__12931\
        );

    \I__2474\ : Span12Mux_s8_h
    port map (
            O => \N__12949\,
            I => \N__12931\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__12946\,
            I => \N__12931\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__12943\,
            I => \N__12931\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__12940\,
            I => \M_this_vram_read_data_3\
        );

    \I__2470\ : Odrv12
    port map (
            O => \N__12931\,
            I => \M_this_vram_read_data_3\
        );

    \I__2469\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12923\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__12923\,
            I => \N__12920\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__12920\,
            I => \N__12917\
        );

    \I__2466\ : Span4Mux_h
    port map (
            O => \N__12917\,
            I => \N__12914\
        );

    \I__2465\ : Span4Mux_h
    port map (
            O => \N__12914\,
            I => \N__12911\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__12911\,
            I => \this_vga_signals.rgb_bmZ0Z_0\
        );

    \I__2463\ : InMux
    port map (
            O => \N__12908\,
            I => \N__12905\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__12905\,
            I => \N__12902\
        );

    \I__2461\ : Odrv12
    port map (
            O => \N__12902\,
            I => \this_vga_signals.rgb_bmZ0Z_2\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__12899\,
            I => \m7_am_cascade_\
        );

    \I__2459\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12893\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__12893\,
            I => m7_ns
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__12890\,
            I => \m28_cascade_\
        );

    \I__2456\ : InMux
    port map (
            O => \N__12887\,
            I => \un1_M_current_address_q_cry_3\
        );

    \I__2455\ : InMux
    port map (
            O => \N__12884\,
            I => \un1_M_current_address_q_cry_4\
        );

    \I__2454\ : InMux
    port map (
            O => \N__12881\,
            I => \un1_M_current_address_q_cry_5\
        );

    \I__2453\ : InMux
    port map (
            O => \N__12878\,
            I => \un1_M_current_address_q_cry_6\
        );

    \I__2452\ : InMux
    port map (
            O => \N__12875\,
            I => \bfn_15_22_0_\
        );

    \I__2451\ : InMux
    port map (
            O => \N__12872\,
            I => \un1_M_current_address_q_cry_8\
        );

    \I__2450\ : InMux
    port map (
            O => \N__12869\,
            I => \un1_M_current_address_q_cry_9\
        );

    \I__2449\ : InMux
    port map (
            O => \N__12866\,
            I => \un1_M_current_address_q_cry_10\
        );

    \I__2448\ : InMux
    port map (
            O => \N__12863\,
            I => \un1_M_current_address_q_cry_11\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__12860\,
            I => \N_349_0_cascade_\
        );

    \I__2446\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12852\
        );

    \I__2445\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12847\
        );

    \I__2444\ : InMux
    port map (
            O => \N__12855\,
            I => \N__12847\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__12852\,
            I => \N__12842\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__12847\,
            I => \N__12842\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__12842\,
            I => \N__12838\
        );

    \I__2440\ : InMux
    port map (
            O => \N__12841\,
            I => \N__12835\
        );

    \I__2439\ : Sp12to4
    port map (
            O => \N__12838\,
            I => \N__12830\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__12835\,
            I => \N__12830\
        );

    \I__2437\ : Span12Mux_h
    port map (
            O => \N__12830\,
            I => \N__12827\
        );

    \I__2436\ : Odrv12
    port map (
            O => \N__12827\,
            I => port_enb_c
        );

    \I__2435\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12818\
        );

    \I__2434\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12811\
        );

    \I__2433\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12811\
        );

    \I__2432\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12811\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__12818\,
            I => \N__12808\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__12811\,
            I => \N__12805\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__12808\,
            I => \this_delay_clk.M_this_delay_clk_out_0\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__12805\,
            I => \this_delay_clk.M_this_delay_clk_out_0\
        );

    \I__2427\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12797\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__12797\,
            I => debug_0
        );

    \I__2425\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12791\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__12791\,
            I => \N__12788\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__12788\,
            I => \N__12785\
        );

    \I__2422\ : Sp12to4
    port map (
            O => \N__12785\,
            I => \N__12782\
        );

    \I__2421\ : Span12Mux_h
    port map (
            O => \N__12782\,
            I => \N__12778\
        );

    \I__2420\ : InMux
    port map (
            O => \N__12781\,
            I => \N__12775\
        );

    \I__2419\ : Odrv12
    port map (
            O => \N__12778\,
            I => port_rw_c
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__12775\,
            I => port_rw_c
        );

    \I__2417\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__12767\,
            I => \N__12764\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__12764\,
            I => \N__12761\
        );

    \I__2414\ : Sp12to4
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__2413\ : Span12Mux_h
    port map (
            O => \N__12758\,
            I => \N__12755\
        );

    \I__2412\ : Span12Mux_v
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__12752\,
            I => port_address_c_7
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__12749\,
            I => \debug_0_cascade_\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__12746\,
            I => \N__12741\
        );

    \I__2408\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12734\
        );

    \I__2407\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12734\
        );

    \I__2406\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12734\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__12734\,
            I => \this_start_data_delay_M_last_q\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__2403\ : CascadeBuf
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__12725\,
            I => \N__12722\
        );

    \I__2401\ : CascadeBuf
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__12719\,
            I => \N__12716\
        );

    \I__2399\ : CascadeBuf
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__12713\,
            I => \N__12710\
        );

    \I__2397\ : CascadeBuf
    port map (
            O => \N__12710\,
            I => \N__12707\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__12707\,
            I => \N__12704\
        );

    \I__2395\ : CascadeBuf
    port map (
            O => \N__12704\,
            I => \N__12701\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__12701\,
            I => \N__12698\
        );

    \I__2393\ : CascadeBuf
    port map (
            O => \N__12698\,
            I => \N__12695\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__12695\,
            I => \N__12692\
        );

    \I__2391\ : CascadeBuf
    port map (
            O => \N__12692\,
            I => \N__12689\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__12689\,
            I => \N__12686\
        );

    \I__2389\ : CascadeBuf
    port map (
            O => \N__12686\,
            I => \N__12683\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__12683\,
            I => \N__12680\
        );

    \I__2387\ : CascadeBuf
    port map (
            O => \N__12680\,
            I => \N__12677\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__2385\ : CascadeBuf
    port map (
            O => \N__12674\,
            I => \N__12671\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__2383\ : CascadeBuf
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__2381\ : CascadeBuf
    port map (
            O => \N__12662\,
            I => \N__12659\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__2379\ : CascadeBuf
    port map (
            O => \N__12656\,
            I => \N__12653\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__12653\,
            I => \N__12650\
        );

    \I__2377\ : CascadeBuf
    port map (
            O => \N__12650\,
            I => \N__12647\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__12647\,
            I => \N__12644\
        );

    \I__2375\ : CascadeBuf
    port map (
            O => \N__12644\,
            I => \N__12641\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__12641\,
            I => \N__12638\
        );

    \I__2373\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12635\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__12635\,
            I => \N__12632\
        );

    \I__2371\ : Sp12to4
    port map (
            O => \N__12632\,
            I => \N__12629\
        );

    \I__2370\ : Span12Mux_s4_v
    port map (
            O => \N__12629\,
            I => \N__12624\
        );

    \I__2369\ : InMux
    port map (
            O => \N__12628\,
            I => \N__12621\
        );

    \I__2368\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12618\
        );

    \I__2367\ : Span12Mux_h
    port map (
            O => \N__12624\,
            I => \N__12615\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__12621\,
            I => \M_current_address_qZ0Z_0\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__12618\,
            I => \M_current_address_qZ0Z_0\
        );

    \I__2364\ : Odrv12
    port map (
            O => \N__12615\,
            I => \M_current_address_qZ0Z_0\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__12608\,
            I => \N__12604\
        );

    \I__2362\ : InMux
    port map (
            O => \N__12607\,
            I => \N__12601\
        );

    \I__2361\ : InMux
    port map (
            O => \N__12604\,
            I => \N__12598\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12601\,
            I => \N_312_0\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__12598\,
            I => \N_312_0\
        );

    \I__2358\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12590\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__12590\,
            I => \M_current_address_q_RNO_1Z0Z_0\
        );

    \I__2356\ : InMux
    port map (
            O => \N__12587\,
            I => \un1_M_current_address_q_cry_0\
        );

    \I__2355\ : InMux
    port map (
            O => \N__12584\,
            I => \un1_M_current_address_q_cry_1\
        );

    \I__2354\ : InMux
    port map (
            O => \N__12581\,
            I => \un1_M_current_address_q_cry_2\
        );

    \I__2353\ : InMux
    port map (
            O => \N__12578\,
            I => \N__12575\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__12575\,
            I => \this_vga_signals.if_N_16_i_0\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__12569\,
            I => \N__12566\
        );

    \I__2349\ : Odrv12
    port map (
            O => \N__12566\,
            I => \this_vga_signals.g0_1_N_5L8\
        );

    \I__2348\ : InMux
    port map (
            O => \N__12563\,
            I => \N__12559\
        );

    \I__2347\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12556\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__12559\,
            I => \N__12553\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__12556\,
            I => \N__12549\
        );

    \I__2344\ : Span12Mux_h
    port map (
            O => \N__12553\,
            I => \N__12545\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12552\,
            I => \N__12542\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__12549\,
            I => \N__12539\
        );

    \I__2341\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12536\
        );

    \I__2340\ : Odrv12
    port map (
            O => \N__12545\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__12542\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__12539\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__12536\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\
        );

    \I__2336\ : InMux
    port map (
            O => \N__12527\,
            I => \N__12524\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__12524\,
            I => \N__12520\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__12523\,
            I => \N__12517\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__12520\,
            I => \N__12513\
        );

    \I__2332\ : InMux
    port map (
            O => \N__12517\,
            I => \N__12510\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12516\,
            I => \N__12505\
        );

    \I__2330\ : Sp12to4
    port map (
            O => \N__12513\,
            I => \N__12500\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__12510\,
            I => \N__12500\
        );

    \I__2328\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12497\
        );

    \I__2327\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12494\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__12505\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2325\ : Odrv12
    port map (
            O => \N__12500\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__12497\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12494\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_d\
        );

    \I__2322\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12482\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__12482\,
            I => \N__12479\
        );

    \I__2320\ : Odrv12
    port map (
            O => \N__12479\,
            I => \this_vga_signals.g0_1_N_3L3\
        );

    \I__2319\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12470\
        );

    \I__2318\ : InMux
    port map (
            O => \N__12475\,
            I => \N__12467\
        );

    \I__2317\ : InMux
    port map (
            O => \N__12474\,
            I => \N__12464\
        );

    \I__2316\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12461\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__12470\,
            I => \N__12456\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__12467\,
            I => \N__12453\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__12464\,
            I => \N__12448\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__12461\,
            I => \N__12448\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12460\,
            I => \N__12445\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12442\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__12456\,
            I => \N__12437\
        );

    \I__2308\ : Span4Mux_v
    port map (
            O => \N__12453\,
            I => \N__12434\
        );

    \I__2307\ : Span4Mux_v
    port map (
            O => \N__12448\,
            I => \N__12429\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__12445\,
            I => \N__12429\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12426\
        );

    \I__2304\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12423\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12420\
        );

    \I__2302\ : Span4Mux_v
    port map (
            O => \N__12437\,
            I => \N__12415\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__12434\,
            I => \N__12415\
        );

    \I__2300\ : Span4Mux_h
    port map (
            O => \N__12429\,
            I => \N__12410\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__12426\,
            I => \N__12410\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__12423\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__12420\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__12415\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__12410\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__12401\,
            I => \this_vga_signals.g0_1_N_6L11_cascade_\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__12398\,
            I => \N__12395\
        );

    \I__2292\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12391\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12394\,
            I => \N__12387\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__12391\,
            I => \N__12384\
        );

    \I__2289\ : InMux
    port map (
            O => \N__12390\,
            I => \N__12381\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__12387\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__12384\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__12381\,
            I => \this_vga_signals.mult1_un61_sum_c2_0\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12374\,
            I => \N__12371\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__12371\,
            I => \this_vga_signals.g0_1_N_7L13\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__12368\,
            I => \this_vga_signals.g0_1_N_8L15_cascade_\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__12365\,
            I => \N__12360\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__12364\,
            I => \N__12357\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__12363\,
            I => \N__12344\
        );

    \I__2279\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12337\
        );

    \I__2278\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12337\
        );

    \I__2277\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12337\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__12355\,
            I => \N__12327\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__12354\,
            I => \N__12324\
        );

    \I__2274\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12321\
        );

    \I__2273\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12316\
        );

    \I__2272\ : InMux
    port map (
            O => \N__12351\,
            I => \N__12316\
        );

    \I__2271\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12313\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12306\
        );

    \I__2269\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12306\
        );

    \I__2268\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12306\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12344\,
            I => \N__12301\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12337\,
            I => \N__12298\
        );

    \I__2265\ : InMux
    port map (
            O => \N__12336\,
            I => \N__12294\
        );

    \I__2264\ : InMux
    port map (
            O => \N__12335\,
            I => \N__12291\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12334\,
            I => \N__12286\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12333\,
            I => \N__12286\
        );

    \I__2261\ : InMux
    port map (
            O => \N__12332\,
            I => \N__12281\
        );

    \I__2260\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12281\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12278\
        );

    \I__2258\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12273\
        );

    \I__2257\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12273\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__12321\,
            I => \N__12264\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12316\,
            I => \N__12264\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__12313\,
            I => \N__12264\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__12306\,
            I => \N__12264\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12305\,
            I => \N__12259\
        );

    \I__2251\ : InMux
    port map (
            O => \N__12304\,
            I => \N__12259\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__12301\,
            I => \N__12254\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__12298\,
            I => \N__12251\
        );

    \I__2248\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12248\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12294\,
            I => \N__12242\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12291\,
            I => \N__12242\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12286\,
            I => \N__12237\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__12281\,
            I => \N__12237\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12234\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__12273\,
            I => \N__12227\
        );

    \I__2241\ : Span4Mux_v
    port map (
            O => \N__12264\,
            I => \N__12227\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__12259\,
            I => \N__12227\
        );

    \I__2239\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12224\
        );

    \I__2238\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12221\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__12254\,
            I => \N__12218\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__12251\,
            I => \N__12215\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__12248\,
            I => \N__12212\
        );

    \I__2234\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12209\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__12242\,
            I => \N__12204\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__12237\,
            I => \N__12204\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__12234\,
            I => \N__12199\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__12227\,
            I => \N__12199\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__12224\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12221\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__12218\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__12215\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__12212\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__12209\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__12204\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__12199\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__12182\,
            I => \N__12175\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12165\
        );

    \I__2219\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12162\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12157\
        );

    \I__2217\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12157\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12152\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12152\
        );

    \I__2214\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12149\
        );

    \I__2213\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12144\
        );

    \I__2212\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12144\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__12170\,
            I => \N__12141\
        );

    \I__2210\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12135\
        );

    \I__2209\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12132\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12165\,
            I => \N__12127\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__12162\,
            I => \N__12127\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__12157\,
            I => \N__12124\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__12152\,
            I => \N__12117\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__12149\,
            I => \N__12117\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12144\,
            I => \N__12117\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12114\
        );

    \I__2201\ : InMux
    port map (
            O => \N__12140\,
            I => \N__12109\
        );

    \I__2200\ : InMux
    port map (
            O => \N__12139\,
            I => \N__12109\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__12138\,
            I => \N__12105\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__12135\,
            I => \N__12102\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__12132\,
            I => \N__12095\
        );

    \I__2196\ : Span4Mux_h
    port map (
            O => \N__12127\,
            I => \N__12095\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__12124\,
            I => \N__12095\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__12117\,
            I => \N__12092\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__12114\,
            I => \N__12087\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12109\,
            I => \N__12087\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12084\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12081\
        );

    \I__2189\ : Span4Mux_h
    port map (
            O => \N__12102\,
            I => \N__12076\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__12095\,
            I => \N__12076\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__12092\,
            I => \N__12073\
        );

    \I__2186\ : Span4Mux_v
    port map (
            O => \N__12087\,
            I => \N__12070\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__12084\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__12081\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__12076\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__12073\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__12070\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12052\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12049\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12046\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12041\
        );

    \I__2176\ : InMux
    port map (
            O => \N__12055\,
            I => \N__12041\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12052\,
            I => \this_vga_signals.mult1_un68_sum_axb2_0\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12049\,
            I => \this_vga_signals.mult1_un68_sum_axb2_0\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__12046\,
            I => \this_vga_signals.mult1_un68_sum_axb2_0\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12041\,
            I => \this_vga_signals.mult1_un68_sum_axb2_0\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__12032\,
            I => \this_vga_signals.mult1_un68_sum_c2_0_0_cascade_\
        );

    \I__2170\ : InMux
    port map (
            O => \N__12029\,
            I => \N__12026\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__12026\,
            I => \this_vga_signals.if_N_6_3_0\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__12023\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0_cascade_\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__12020\,
            I => \N__12017\
        );

    \I__2166\ : CascadeBuf
    port map (
            O => \N__12017\,
            I => \N__12014\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__12014\,
            I => \N__12011\
        );

    \I__2164\ : CascadeBuf
    port map (
            O => \N__12011\,
            I => \N__12008\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__12008\,
            I => \N__12005\
        );

    \I__2162\ : CascadeBuf
    port map (
            O => \N__12005\,
            I => \N__12002\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__12002\,
            I => \N__11999\
        );

    \I__2160\ : CascadeBuf
    port map (
            O => \N__11999\,
            I => \N__11996\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__11996\,
            I => \N__11993\
        );

    \I__2158\ : CascadeBuf
    port map (
            O => \N__11993\,
            I => \N__11990\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__11990\,
            I => \N__11987\
        );

    \I__2156\ : CascadeBuf
    port map (
            O => \N__11987\,
            I => \N__11984\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__11984\,
            I => \N__11981\
        );

    \I__2154\ : CascadeBuf
    port map (
            O => \N__11981\,
            I => \N__11978\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__11978\,
            I => \N__11975\
        );

    \I__2152\ : CascadeBuf
    port map (
            O => \N__11975\,
            I => \N__11972\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__11972\,
            I => \N__11969\
        );

    \I__2150\ : CascadeBuf
    port map (
            O => \N__11969\,
            I => \N__11966\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__11966\,
            I => \N__11963\
        );

    \I__2148\ : CascadeBuf
    port map (
            O => \N__11963\,
            I => \N__11960\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__2146\ : CascadeBuf
    port map (
            O => \N__11957\,
            I => \N__11954\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__11954\,
            I => \N__11951\
        );

    \I__2144\ : CascadeBuf
    port map (
            O => \N__11951\,
            I => \N__11948\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__11948\,
            I => \N__11945\
        );

    \I__2142\ : CascadeBuf
    port map (
            O => \N__11945\,
            I => \N__11942\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__11942\,
            I => \N__11939\
        );

    \I__2140\ : CascadeBuf
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__11936\,
            I => \N__11933\
        );

    \I__2138\ : CascadeBuf
    port map (
            O => \N__11933\,
            I => \N__11930\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__11930\,
            I => \N__11927\
        );

    \I__2136\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11924\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__11924\,
            I => \N__11921\
        );

    \I__2134\ : Sp12to4
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__2133\ : Span12Mux_v
    port map (
            O => \N__11918\,
            I => \N__11915\
        );

    \I__2132\ : Odrv12
    port map (
            O => \N__11915\,
            I => \M_this_vga_signals_address_8\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__11912\,
            I => \N__11909\
        );

    \I__2130\ : InMux
    port map (
            O => \N__11909\,
            I => \N__11906\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__11906\,
            I => \N_401\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__11903\,
            I => \N__11898\
        );

    \I__2127\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11893\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11888\
        );

    \I__2125\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11888\
        );

    \I__2124\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11885\
        );

    \I__2123\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11882\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__11893\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__11888\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__11885\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__11882\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\
        );

    \I__2118\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11867\
        );

    \I__2117\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11864\
        );

    \I__2116\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11859\
        );

    \I__2115\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11859\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__11867\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__11864\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__11859\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__11852\,
            I => \N__11849\
        );

    \I__2110\ : CascadeBuf
    port map (
            O => \N__11849\,
            I => \N__11846\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__11846\,
            I => \N__11843\
        );

    \I__2108\ : CascadeBuf
    port map (
            O => \N__11843\,
            I => \N__11840\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__11840\,
            I => \N__11837\
        );

    \I__2106\ : CascadeBuf
    port map (
            O => \N__11837\,
            I => \N__11834\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__11834\,
            I => \N__11831\
        );

    \I__2104\ : CascadeBuf
    port map (
            O => \N__11831\,
            I => \N__11828\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__2102\ : CascadeBuf
    port map (
            O => \N__11825\,
            I => \N__11822\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__11822\,
            I => \N__11819\
        );

    \I__2100\ : CascadeBuf
    port map (
            O => \N__11819\,
            I => \N__11816\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__11816\,
            I => \N__11813\
        );

    \I__2098\ : CascadeBuf
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__11810\,
            I => \N__11807\
        );

    \I__2096\ : CascadeBuf
    port map (
            O => \N__11807\,
            I => \N__11804\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__11804\,
            I => \N__11801\
        );

    \I__2094\ : CascadeBuf
    port map (
            O => \N__11801\,
            I => \N__11798\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__11798\,
            I => \N__11795\
        );

    \I__2092\ : CascadeBuf
    port map (
            O => \N__11795\,
            I => \N__11792\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__11792\,
            I => \N__11789\
        );

    \I__2090\ : CascadeBuf
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__2088\ : CascadeBuf
    port map (
            O => \N__11783\,
            I => \N__11780\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__2086\ : CascadeBuf
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__11774\,
            I => \N__11771\
        );

    \I__2084\ : CascadeBuf
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__2082\ : CascadeBuf
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__11762\,
            I => \N__11759\
        );

    \I__2080\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__2078\ : Span12Mux_h
    port map (
            O => \N__11753\,
            I => \N__11750\
        );

    \I__2077\ : Odrv12
    port map (
            O => \N__11750\,
            I => \M_this_vga_signals_address_4\
        );

    \I__2076\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11742\
        );

    \I__2075\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11737\
        );

    \I__2074\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11737\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__11742\,
            I => \N__11732\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__11737\,
            I => \N__11729\
        );

    \I__2071\ : InMux
    port map (
            O => \N__11736\,
            I => \N__11726\
        );

    \I__2070\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11723\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__11732\,
            I => \N__11720\
        );

    \I__2068\ : Span4Mux_h
    port map (
            O => \N__11729\,
            I => \N__11715\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__11726\,
            I => \N__11715\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__11723\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__11720\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__11715\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__2063\ : InMux
    port map (
            O => \N__11708\,
            I => \N__11694\
        );

    \I__2062\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11694\
        );

    \I__2061\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11690\
        );

    \I__2060\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11677\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11677\
        );

    \I__2058\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11677\
        );

    \I__2057\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11677\
        );

    \I__2056\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11670\
        );

    \I__2055\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11670\
        );

    \I__2054\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11670\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__11694\,
            I => \N__11667\
        );

    \I__2052\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11664\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__11690\,
            I => \N__11661\
        );

    \I__2050\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11655\
        );

    \I__2049\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11655\
        );

    \I__2048\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11650\
        );

    \I__2047\ : InMux
    port map (
            O => \N__11686\,
            I => \N__11650\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__11677\,
            I => \N__11647\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__11670\,
            I => \N__11644\
        );

    \I__2044\ : Span4Mux_h
    port map (
            O => \N__11667\,
            I => \N__11639\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__11664\,
            I => \N__11639\
        );

    \I__2042\ : Span12Mux_v
    port map (
            O => \N__11661\,
            I => \N__11636\
        );

    \I__2041\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11633\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__11655\,
            I => \M_counter_q_RNIJR071_1\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__11650\,
            I => \M_counter_q_RNIJR071_1\
        );

    \I__2038\ : Odrv12
    port map (
            O => \N__11647\,
            I => \M_counter_q_RNIJR071_1\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__11644\,
            I => \M_counter_q_RNIJR071_1\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__11639\,
            I => \M_counter_q_RNIJR071_1\
        );

    \I__2035\ : Odrv12
    port map (
            O => \N__11636\,
            I => \M_counter_q_RNIJR071_1\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__11633\,
            I => \M_counter_q_RNIJR071_1\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11611\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__11614\,
            I => \N__11607\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__11611\,
            I => \N__11603\
        );

    \I__2029\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11600\
        );

    \I__2028\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11595\
        );

    \I__2027\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11595\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__11603\,
            I => \N__11592\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__11600\,
            I => \N__11589\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__11595\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__11592\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__11589\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__2021\ : SRMux
    port map (
            O => \N__11582\,
            I => \N__11579\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__11579\,
            I => \N__11574\
        );

    \I__2019\ : SRMux
    port map (
            O => \N__11578\,
            I => \N__11571\
        );

    \I__2018\ : SRMux
    port map (
            O => \N__11577\,
            I => \N__11568\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__11574\,
            I => \N__11562\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__11571\,
            I => \N__11562\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__11568\,
            I => \N__11559\
        );

    \I__2014\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11556\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__11562\,
            I => \N__11553\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__11559\,
            I => \N__11550\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__11556\,
            I => \N__11547\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__11553\,
            I => \M_counter_q_RNIQR4I2_1\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__11550\,
            I => \M_counter_q_RNIQR4I2_1\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__11547\,
            I => \M_counter_q_RNIQR4I2_1\
        );

    \I__2007\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__11537\,
            I => \N__11534\
        );

    \I__2005\ : Odrv12
    port map (
            O => \N__11534\,
            I => \this_vga_signals.rgb_bmZ0Z_1\
        );

    \I__2004\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11528\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__11528\,
            I => \N__11525\
        );

    \I__2002\ : Span4Mux_h
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__2001\ : Span4Mux_h
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__11519\,
            I => \N__11516\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__11516\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__1998\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11509\
        );

    \I__1997\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11506\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__11509\,
            I => \N__11500\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__11506\,
            I => \N__11497\
        );

    \I__1994\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11493\
        );

    \I__1993\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11488\
        );

    \I__1992\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11488\
        );

    \I__1991\ : Span4Mux_h
    port map (
            O => \N__11500\,
            I => \N__11485\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__11497\,
            I => \N__11482\
        );

    \I__1989\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11479\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__11493\,
            I => \N__11474\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__11488\,
            I => \N__11474\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__11485\,
            I => \this_vga_signals.mult1_un54_sum_axb1_5\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__11482\,
            I => \this_vga_signals.mult1_un54_sum_axb1_5\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__11479\,
            I => \this_vga_signals.mult1_un54_sum_axb1_5\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__11474\,
            I => \this_vga_signals.mult1_un54_sum_axb1_5\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__11465\,
            I => \N__11452\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__11464\,
            I => \N__11447\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__11463\,
            I => \N__11444\
        );

    \I__1979\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11439\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__11461\,
            I => \N__11432\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__11460\,
            I => \N__11429\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__11459\,
            I => \N__11423\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__11458\,
            I => \N__11419\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__11457\,
            I => \N__11414\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__11456\,
            I => \N__11410\
        );

    \I__1972\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11403\
        );

    \I__1971\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11396\
        );

    \I__1970\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11396\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11396\
        );

    \I__1968\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11391\
        );

    \I__1967\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11388\
        );

    \I__1966\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11383\
        );

    \I__1965\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11383\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__11439\,
            I => \N__11380\
        );

    \I__1963\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11377\
        );

    \I__1962\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11368\
        );

    \I__1961\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11368\
        );

    \I__1960\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11368\
        );

    \I__1959\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11368\
        );

    \I__1958\ : InMux
    port map (
            O => \N__11429\,
            I => \N__11363\
        );

    \I__1957\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11363\
        );

    \I__1956\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11360\
        );

    \I__1955\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11357\
        );

    \I__1954\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11354\
        );

    \I__1953\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11349\
        );

    \I__1952\ : InMux
    port map (
            O => \N__11419\,
            I => \N__11349\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__11418\,
            I => \N__11345\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11417\,
            I => \N__11342\
        );

    \I__1949\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11337\
        );

    \I__1948\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11337\
        );

    \I__1947\ : InMux
    port map (
            O => \N__11410\,
            I => \N__11332\
        );

    \I__1946\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11332\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__11408\,
            I => \N__11328\
        );

    \I__1944\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11323\
        );

    \I__1943\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11323\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__11403\,
            I => \N__11318\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11396\,
            I => \N__11318\
        );

    \I__1940\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11313\
        );

    \I__1939\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11313\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__11391\,
            I => \N__11310\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__11388\,
            I => \N__11307\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__11383\,
            I => \N__11298\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__11380\,
            I => \N__11298\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__11377\,
            I => \N__11298\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__11368\,
            I => \N__11298\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__11363\,
            I => \N__11295\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__11360\,
            I => \N__11290\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__11357\,
            I => \N__11290\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11354\,
            I => \N__11284\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11349\,
            I => \N__11284\
        );

    \I__1927\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11281\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11278\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11271\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__11337\,
            I => \N__11271\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__11332\,
            I => \N__11271\
        );

    \I__1922\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11265\
        );

    \I__1921\ : InMux
    port map (
            O => \N__11328\,
            I => \N__11265\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__11323\,
            I => \N__11262\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__11318\,
            I => \N__11259\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__11313\,
            I => \N__11254\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__11310\,
            I => \N__11254\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__11307\,
            I => \N__11245\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__11298\,
            I => \N__11245\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__11295\,
            I => \N__11245\
        );

    \I__1913\ : Span4Mux_h
    port map (
            O => \N__11290\,
            I => \N__11245\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11289\,
            I => \N__11242\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__11284\,
            I => \N__11235\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11235\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11235\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__11271\,
            I => \N__11232\
        );

    \I__1907\ : InMux
    port map (
            O => \N__11270\,
            I => \N__11229\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__11265\,
            I => \N__11226\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__11262\,
            I => \N__11219\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__11259\,
            I => \N__11219\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__11254\,
            I => \N__11219\
        );

    \I__1902\ : Span4Mux_v
    port map (
            O => \N__11245\,
            I => \N__11216\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__11242\,
            I => \N__11209\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__11235\,
            I => \N__11209\
        );

    \I__1899\ : Span4Mux_h
    port map (
            O => \N__11232\,
            I => \N__11209\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__11229\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__11226\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__11219\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__11216\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__11209\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__11198\,
            I => \this_vga_signals.if_N_13_i_i_0_cascade_\
        );

    \I__1892\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11187\
        );

    \I__1891\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11184\
        );

    \I__1890\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11180\
        );

    \I__1889\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11175\
        );

    \I__1888\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11175\
        );

    \I__1887\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11170\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__11187\,
            I => \N__11166\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11184\,
            I => \N__11163\
        );

    \I__1884\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11160\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__11180\,
            I => \N__11155\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__11175\,
            I => \N__11155\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11150\
        );

    \I__1880\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11150\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__11170\,
            I => \N__11140\
        );

    \I__1878\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11137\
        );

    \I__1877\ : Span4Mux_h
    port map (
            O => \N__11166\,
            I => \N__11126\
        );

    \I__1876\ : Span4Mux_h
    port map (
            O => \N__11163\,
            I => \N__11126\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11160\,
            I => \N__11126\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__11155\,
            I => \N__11126\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__11150\,
            I => \N__11126\
        );

    \I__1872\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11119\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11119\
        );

    \I__1870\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11119\
        );

    \I__1869\ : InMux
    port map (
            O => \N__11146\,
            I => \N__11114\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11114\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11109\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11109\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__11140\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__11137\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__11126\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11119\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11114\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__11109\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_0\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__11096\,
            I => \this_vga_signals.g0_1_0_0_cascade_\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__11087\,
            I => \this_vga_signals.g4_0\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__11084\,
            I => \this_vga_signals.mult1_un68_sum_ac0_3_d_0_cascade_\
        );

    \I__1854\ : InMux
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__11078\,
            I => \N__11073\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11077\,
            I => \N__11070\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11067\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__11073\,
            I => \this_vga_signals.mult1_un68_sum_ac0_4\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__11070\,
            I => \this_vga_signals.mult1_un68_sum_ac0_4\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__11067\,
            I => \this_vga_signals.mult1_un68_sum_ac0_4\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__11060\,
            I => \this_vga_signals.g0_i_o2_0_0_x2_0_cascade_\
        );

    \I__1846\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11054\,
            I => \this_vga_signals.N_16\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__11051\,
            I => \N__11048\
        );

    \I__1843\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__11045\,
            I => \N__11040\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11037\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11034\
        );

    \I__1839\ : Span4Mux_v
    port map (
            O => \N__11040\,
            I => \N__11029\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__11037\,
            I => \N__11029\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__11024\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__11029\,
            I => \N__11021\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11018\
        );

    \I__1834\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11015\
        );

    \I__1833\ : Odrv12
    port map (
            O => \N__11024\,
            I => \this_vga_signals.mult1_un54_sum_i_1\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__11021\,
            I => \this_vga_signals.mult1_un54_sum_i_1\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__11018\,
            I => \this_vga_signals.mult1_un54_sum_i_1\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11015\,
            I => \this_vga_signals.mult1_un54_sum_i_1\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11006\,
            I => \N__11002\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__11005\,
            I => \N__10999\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__11002\,
            I => \N__10996\
        );

    \I__1826\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10993\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__10996\,
            I => \this_vga_signals.if_N_1_i_0\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__10993\,
            I => \this_vga_signals.if_N_1_i_0\
        );

    \I__1823\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10982\
        );

    \I__1822\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10982\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10977\
        );

    \I__1820\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10972\
        );

    \I__1819\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10972\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__10977\,
            I => \N__10959\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__10972\,
            I => \N__10959\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__10971\,
            I => \N__10956\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__10970\,
            I => \N__10953\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__10969\,
            I => \N__10950\
        );

    \I__1813\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10944\
        );

    \I__1812\ : InMux
    port map (
            O => \N__10967\,
            I => \N__10944\
        );

    \I__1811\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10937\
        );

    \I__1810\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10937\
        );

    \I__1809\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10937\
        );

    \I__1808\ : Span4Mux_h
    port map (
            O => \N__10959\,
            I => \N__10934\
        );

    \I__1807\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10925\
        );

    \I__1806\ : InMux
    port map (
            O => \N__10953\,
            I => \N__10925\
        );

    \I__1805\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10925\
        );

    \I__1804\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10925\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__10944\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__10937\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__10934\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__10925\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1799\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10907\
        );

    \I__1798\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10907\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__10914\,
            I => \N__10903\
        );

    \I__1796\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10894\
        );

    \I__1795\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10894\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__10907\,
            I => \N__10891\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10884\
        );

    \I__1792\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10884\
        );

    \I__1791\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10884\
        );

    \I__1790\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10877\
        );

    \I__1789\ : InMux
    port map (
            O => \N__10900\,
            I => \N__10874\
        );

    \I__1788\ : InMux
    port map (
            O => \N__10899\,
            I => \N__10871\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__10894\,
            I => \N__10868\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__10891\,
            I => \N__10865\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__10884\,
            I => \N__10862\
        );

    \I__1784\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10853\
        );

    \I__1783\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10853\
        );

    \I__1782\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10853\
        );

    \I__1781\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10853\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__10877\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__10874\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__10871\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__10868\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__10865\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__10862\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__10853\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__1773\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10835\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__10835\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0\
        );

    \I__1771\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__1769\ : Span4Mux_h
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__10823\,
            I => \this_vga_signals.mult1_un61_sum_axb1\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__10820\,
            I => \this_vga_signals.if_m3_5_cascade_\
        );

    \I__1766\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__10814\,
            I => \this_vga_signals.if_N_3_i\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__10811\,
            I => \this_vga_signals.if_m5_4_cascade_\
        );

    \I__1763\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__10805\,
            I => \this_vga_signals.g1_1_4\
        );

    \I__1761\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10799\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__10799\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_1\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__10796\,
            I => \this_vga_signals.mult1_un68_sum_axb2_0_1_cascade_\
        );

    \I__1758\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__10790\,
            I => \this_vga_signals.g1_1_1\
        );

    \I__1756\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__10784\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_0\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__10781\,
            I => \this_vga_signals.SUM_3_cascade_\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1752\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10766\
        );

    \I__1751\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10763\
        );

    \I__1750\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10758\
        );

    \I__1749\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10758\
        );

    \I__1748\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10751\
        );

    \I__1747\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10751\
        );

    \I__1746\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10751\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__10766\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__10763\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__10758\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10751\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__10742\,
            I => \N__10734\
        );

    \I__1740\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10730\
        );

    \I__1739\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10727\
        );

    \I__1738\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10722\
        );

    \I__1737\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10722\
        );

    \I__1736\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10715\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10715\
        );

    \I__1734\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10715\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__10730\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__10727\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__10722\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__10715\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1729\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10696\
        );

    \I__1728\ : InMux
    port map (
            O => \N__10705\,
            I => \N__10696\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__10704\,
            I => \N__10693\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__10703\,
            I => \N__10690\
        );

    \I__1725\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10686\
        );

    \I__1724\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10683\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__10696\,
            I => \N__10680\
        );

    \I__1722\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10673\
        );

    \I__1721\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10673\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10673\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__10686\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__10683\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__10680\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__10673\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1715\ : InMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__10661\,
            I => \this_vga_signals.N_34\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__10658\,
            I => \this_vga_signals.N_34_cascade_\
        );

    \I__1712\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10650\
        );

    \I__1711\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10645\
        );

    \I__1710\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10645\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__10650\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__10645\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__10640\,
            I => \N__10633\
        );

    \I__1706\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10627\
        );

    \I__1705\ : InMux
    port map (
            O => \N__10638\,
            I => \N__10624\
        );

    \I__1704\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10621\
        );

    \I__1703\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10616\
        );

    \I__1702\ : InMux
    port map (
            O => \N__10633\,
            I => \N__10616\
        );

    \I__1701\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10609\
        );

    \I__1700\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10609\
        );

    \I__1699\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10609\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__10627\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__10624\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__10621\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10616\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__10609\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__10598\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0_cascade_\
        );

    \I__1692\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10584\
        );

    \I__1691\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10581\
        );

    \I__1690\ : InMux
    port map (
            O => \N__10593\,
            I => \N__10578\
        );

    \I__1689\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10575\
        );

    \I__1688\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10564\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10564\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10564\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10564\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10564\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__10584\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__10581\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__10578\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__10575\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__10564\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1678\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10545\
        );

    \I__1677\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10536\
        );

    \I__1676\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10536\
        );

    \I__1675\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10536\
        );

    \I__1674\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10536\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10531\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__10545\,
            I => \N__10526\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__10536\,
            I => \N__10526\
        );

    \I__1670\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10523\
        );

    \I__1669\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10520\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__10531\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__10526\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__10523\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__10520\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1664\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10502\
        );

    \I__1663\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10499\
        );

    \I__1662\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10494\
        );

    \I__1661\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10494\
        );

    \I__1660\ : InMux
    port map (
            O => \N__10507\,
            I => \N__10487\
        );

    \I__1659\ : InMux
    port map (
            O => \N__10506\,
            I => \N__10487\
        );

    \I__1658\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10487\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__10502\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__10499\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__10494\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__10487\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__10478\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10469\
        );

    \I__1651\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10469\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10469\,
            I => \this_vga_signals.mult1_un68_sum_c2_0\
        );

    \I__1649\ : CEMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__10463\,
            I => \N__10460\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__10460\,
            I => \this_vga_signals.N_469_1\
        );

    \I__1646\ : IoInMux
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__1644\ : IoSpan4Mux
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__1643\ : Span4Mux_s3_v
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__1642\ : Sp12to4
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1641\ : Span12Mux_v
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__1640\ : Odrv12
    port map (
            O => \N__10439\,
            I => debug_0_i
        );

    \I__1639\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__1637\ : Span4Mux_h
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__1636\ : Span4Mux_h
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__10424\,
            I => \this_vga_signals.rgb_cnst_i_a5_0_0Z0Z_3\
        );

    \I__1634\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10417\
        );

    \I__1633\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10414\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__10417\,
            I => \N__10405\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10405\
        );

    \I__1630\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10402\
        );

    \I__1629\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10399\
        );

    \I__1628\ : InMux
    port map (
            O => \N__10411\,
            I => \N__10396\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__10410\,
            I => \N__10393\
        );

    \I__1626\ : Span4Mux_v
    port map (
            O => \N__10405\,
            I => \N__10387\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__10402\,
            I => \N__10387\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__10399\,
            I => \N__10382\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__10396\,
            I => \N__10382\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10377\
        );

    \I__1621\ : InMux
    port map (
            O => \N__10392\,
            I => \N__10377\
        );

    \I__1620\ : Span4Mux_h
    port map (
            O => \N__10387\,
            I => \N__10373\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__10382\,
            I => \N__10370\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10377\,
            I => \N__10367\
        );

    \I__1617\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10364\
        );

    \I__1616\ : Span4Mux_h
    port map (
            O => \N__10373\,
            I => \N__10361\
        );

    \I__1615\ : Span4Mux_h
    port map (
            O => \N__10370\,
            I => \N__10354\
        );

    \I__1614\ : Span4Mux_v
    port map (
            O => \N__10367\,
            I => \N__10354\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10354\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__10361\,
            I => \M_this_vram_read_data_0\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__10354\,
            I => \M_this_vram_read_data_0\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__10349\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__10346\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__10343\,
            I => \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\
        );

    \I__1607\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__10337\,
            I => \this_vga_signals.mult1_un61_sum_axbxc1\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \N__10327\
        );

    \I__1604\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10318\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10318\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10318\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10313\
        );

    \I__1600\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10313\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__10326\,
            I => \N__10310\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10305\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10300\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10300\
        );

    \I__1595\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10293\
        );

    \I__1594\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10293\
        );

    \I__1593\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10293\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__10305\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__10300\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__10293\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__10286\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_0_0_cascade_\
        );

    \I__1588\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__10280\,
            I => \this_vga_signals.if_N_9_0_0\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10269\
        );

    \I__1585\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10269\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10264\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10264\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__10269\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__10264\,
            I => \this_vga_signals.mult1_un68_sum_axb1\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__1579\ : CascadeBuf
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1577\ : CascadeBuf
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__1575\ : CascadeBuf
    port map (
            O => \N__10244\,
            I => \N__10241\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__10241\,
            I => \N__10238\
        );

    \I__1573\ : CascadeBuf
    port map (
            O => \N__10238\,
            I => \N__10235\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__10235\,
            I => \N__10232\
        );

    \I__1571\ : CascadeBuf
    port map (
            O => \N__10232\,
            I => \N__10229\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__10229\,
            I => \N__10226\
        );

    \I__1569\ : CascadeBuf
    port map (
            O => \N__10226\,
            I => \N__10223\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__10223\,
            I => \N__10220\
        );

    \I__1567\ : CascadeBuf
    port map (
            O => \N__10220\,
            I => \N__10217\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__1565\ : CascadeBuf
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__1563\ : CascadeBuf
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__10205\,
            I => \N__10202\
        );

    \I__1561\ : CascadeBuf
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__10199\,
            I => \N__10196\
        );

    \I__1559\ : CascadeBuf
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__1557\ : CascadeBuf
    port map (
            O => \N__10190\,
            I => \N__10187\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__10187\,
            I => \N__10184\
        );

    \I__1555\ : CascadeBuf
    port map (
            O => \N__10184\,
            I => \N__10181\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__10181\,
            I => \N__10178\
        );

    \I__1553\ : CascadeBuf
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__1551\ : CascadeBuf
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10163\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__10163\,
            I => \N__10160\
        );

    \I__1547\ : Span12Mux_s2_v
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1546\ : Span12Mux_h
    port map (
            O => \N__10157\,
            I => \N__10154\
        );

    \I__1545\ : Odrv12
    port map (
            O => \N__10154\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__10151\,
            I => \this_vga_signals.if_N_8_i_cascade_\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__10145\,
            I => \this_vga_signals.mult1_un82_sum_axb1\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__10139\,
            I => \this_vga_signals.mult1_un89_sum_c3\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__10136\,
            I => \this_vga_signals.mult1_un82_sum_c3_cascade_\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__10133\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_\
        );

    \I__1537\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10127\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_2\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10121\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__10121\,
            I => \this_vga_signals.mult1_un82_sum_c2_0\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10118\,
            I => \N__10115\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__10115\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_0\
        );

    \I__1531\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__10109\,
            I => \this_vga_signals.g0_i_x2_5\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__10106\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10100\,
            I => \this_vga_signals.N_9_1_0\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__10088\,
            I => \this_vga_signals.g1_5\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10082\,
            I => \this_vga_signals.N_6\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__10079\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_0_0_1_cascade_\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__1518\ : CascadeBuf
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__1516\ : CascadeBuf
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__1514\ : CascadeBuf
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__1512\ : CascadeBuf
    port map (
            O => \N__10055\,
            I => \N__10052\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__1510\ : CascadeBuf
    port map (
            O => \N__10049\,
            I => \N__10046\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__1508\ : CascadeBuf
    port map (
            O => \N__10043\,
            I => \N__10040\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10040\,
            I => \N__10037\
        );

    \I__1506\ : CascadeBuf
    port map (
            O => \N__10037\,
            I => \N__10034\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__10034\,
            I => \N__10031\
        );

    \I__1504\ : CascadeBuf
    port map (
            O => \N__10031\,
            I => \N__10028\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__10028\,
            I => \N__10025\
        );

    \I__1502\ : CascadeBuf
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__10022\,
            I => \N__10019\
        );

    \I__1500\ : CascadeBuf
    port map (
            O => \N__10019\,
            I => \N__10016\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__10016\,
            I => \N__10013\
        );

    \I__1498\ : CascadeBuf
    port map (
            O => \N__10013\,
            I => \N__10010\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__10010\,
            I => \N__10007\
        );

    \I__1496\ : CascadeBuf
    port map (
            O => \N__10007\,
            I => \N__10004\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__10004\,
            I => \N__10001\
        );

    \I__1494\ : CascadeBuf
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__1492\ : CascadeBuf
    port map (
            O => \N__9995\,
            I => \N__9992\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__1490\ : CascadeBuf
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__1488\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9980\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__1485\ : Span4Mux_v
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__1483\ : Span4Mux_h
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__9962\,
            I => \M_this_vga_signals_address_7\
        );

    \I__1480\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__9956\,
            I => \this_vga_signals.g2_0_1_0\
        );

    \I__1478\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__9950\,
            I => \this_vga_signals.g0_i_x2_2\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__9947\,
            I => \this_vga_signals.g0_i_0_N_4L5_cascade_\
        );

    \I__1475\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__9941\,
            I => \this_vga_signals.g0_i_0_N_5L7\
        );

    \I__1473\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9935\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__9935\,
            I => \this_vga_signals.if_i4_mux_0_0_0_1\
        );

    \I__1471\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9929\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__9929\,
            I => \this_vga_signals.N_6_i\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__1468\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1466\ : Span4Mux_v
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__9914\,
            I => \this_vga_signals.g1_1_2\
        );

    \I__1464\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__9908\,
            I => \this_vga_signals.g1_4_1\
        );

    \I__1462\ : InMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__9902\,
            I => \N__9898\
        );

    \I__1460\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9894\
        );

    \I__1459\ : Span4Mux_h
    port map (
            O => \N__9898\,
            I => \N__9891\
        );

    \I__1458\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9888\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__9894\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__9891\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__9888\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__1454\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9878\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__9878\,
            I => \this_vga_signals.g0_i_0_N_2L1\
        );

    \I__1452\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9868\
        );

    \I__1451\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9868\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__9873\,
            I => \N__9864\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__9868\,
            I => \N__9856\
        );

    \I__1448\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9853\
        );

    \I__1447\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9849\
        );

    \I__1446\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9844\
        );

    \I__1445\ : InMux
    port map (
            O => \N__9862\,
            I => \N__9844\
        );

    \I__1444\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9841\
        );

    \I__1443\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9836\
        );

    \I__1442\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9836\
        );

    \I__1441\ : Span4Mux_v
    port map (
            O => \N__9856\,
            I => \N__9825\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__9853\,
            I => \N__9825\
        );

    \I__1439\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9822\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9814\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__9844\,
            I => \N__9814\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__9841\,
            I => \N__9814\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9811\
        );

    \I__1434\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9808\
        );

    \I__1433\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9801\
        );

    \I__1432\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9801\
        );

    \I__1431\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9801\
        );

    \I__1430\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9796\
        );

    \I__1429\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9796\
        );

    \I__1428\ : Span4Mux_h
    port map (
            O => \N__9825\,
            I => \N__9785\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__9822\,
            I => \N__9785\
        );

    \I__1426\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9782\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__9814\,
            I => \N__9775\
        );

    \I__1424\ : Span4Mux_v
    port map (
            O => \N__9811\,
            I => \N__9775\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__9808\,
            I => \N__9775\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__9801\,
            I => \N__9770\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__9796\,
            I => \N__9770\
        );

    \I__1420\ : InMux
    port map (
            O => \N__9795\,
            I => \N__9763\
        );

    \I__1419\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9763\
        );

    \I__1418\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9763\
        );

    \I__1417\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9756\
        );

    \I__1416\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9756\
        );

    \I__1415\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9756\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__9785\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__9782\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__9775\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__9770\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__9763\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__9756\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__1408\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9736\
        );

    \I__1407\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9733\
        );

    \I__1406\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9729\
        );

    \I__1405\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9722\
        );

    \I__1404\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9722\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__9736\,
            I => \N__9718\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__9733\,
            I => \N__9715\
        );

    \I__1401\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9712\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__9729\,
            I => \N__9706\
        );

    \I__1399\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9701\
        );

    \I__1398\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9701\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__9722\,
            I => \N__9698\
        );

    \I__1396\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9694\
        );

    \I__1395\ : Span4Mux_h
    port map (
            O => \N__9718\,
            I => \N__9691\
        );

    \I__1394\ : Span4Mux_h
    port map (
            O => \N__9715\,
            I => \N__9688\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9712\,
            I => \N__9685\
        );

    \I__1392\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9680\
        );

    \I__1391\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9680\
        );

    \I__1390\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9677\
        );

    \I__1389\ : Span4Mux_h
    port map (
            O => \N__9706\,
            I => \N__9670\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__9701\,
            I => \N__9670\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__9698\,
            I => \N__9670\
        );

    \I__1386\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9667\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__9694\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__9691\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__9688\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__9685\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__9680\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__9677\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__9670\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__9667\,
            I => \this_vga_signals.M_vcounter_qZ0Z_7\
        );

    \I__1377\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__9647\,
            I => \N__9644\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__9641\,
            I => \this_vga_signals.M_vcounter_d_1_sqmuxa_i_a3_1\
        );

    \I__1373\ : InMux
    port map (
            O => \N__9638\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1372\ : InMux
    port map (
            O => \N__9635\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1371\ : InMux
    port map (
            O => \N__9632\,
            I => \bfn_12_25_0_\
        );

    \I__1370\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9626\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__9623\,
            I => \this_vga_signals.N_22\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__9620\,
            I => \this_vga_signals.g1_0_0_2_cascade_\
        );

    \I__1366\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9614\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__9614\,
            I => \this_vga_signals.N_21\
        );

    \I__1364\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9608\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__1362\ : Odrv12
    port map (
            O => \N__9605\,
            I => \this_vga_signals.g0_i_x2_1\
        );

    \I__1361\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9599\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__9599\,
            I => \this_vga_signals.g4_1\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__9596\,
            I => \this_vga_signals.g0_1_0_cascade_\
        );

    \I__1358\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__9590\,
            I => \N__9586\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9583\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__9586\,
            I => \this_vga_signals.CO0_i_i\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__9583\,
            I => \this_vga_signals.CO0_i_i\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__9578\,
            I => \this_vga_signals.N_45_cascade_\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__9575\,
            I => \N__9571\
        );

    \I__1351\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9567\
        );

    \I__1350\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9564\
        );

    \I__1349\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9561\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__9567\,
            I => \N_23_0\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__9564\,
            I => \N_23_0\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__9561\,
            I => \N_23_0\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__9554\,
            I => \N_23_0_cascade_\
        );

    \I__1344\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9546\
        );

    \I__1343\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9541\
        );

    \I__1342\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9541\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__9546\,
            I => \this_pixel_clock.M_counter_q_i_1\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__9541\,
            I => \this_pixel_clock.M_counter_q_i_1\
        );

    \I__1339\ : InMux
    port map (
            O => \N__9536\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1338\ : InMux
    port map (
            O => \N__9533\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1337\ : InMux
    port map (
            O => \N__9530\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1336\ : InMux
    port map (
            O => \N__9527\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1335\ : InMux
    port map (
            O => \N__9524\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__9521\,
            I => \this_vga_signals.N_28_0_cascade_\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__9518\,
            I => \this_vga_signals.N_42_cascade_\
        );

    \I__1332\ : IoInMux
    port map (
            O => \N__9515\,
            I => \N__9512\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__9512\,
            I => \N__9509\
        );

    \I__1330\ : Span4Mux_s2_v
    port map (
            O => \N__9509\,
            I => \N__9506\
        );

    \I__1329\ : Span4Mux_v
    port map (
            O => \N__9506\,
            I => \N__9503\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__9500\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIVV6F6Z0Z_9\
        );

    \I__1326\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9492\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9496\,
            I => \N__9489\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9486\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__9492\,
            I => \N__9481\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__9489\,
            I => \N__9476\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__9486\,
            I => \N__9476\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__9485\,
            I => \N__9466\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__9484\,
            I => \N__9462\
        );

    \I__1318\ : Span4Mux_v
    port map (
            O => \N__9481\,
            I => \N__9459\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__9476\,
            I => \N__9456\
        );

    \I__1316\ : InMux
    port map (
            O => \N__9475\,
            I => \N__9453\
        );

    \I__1315\ : InMux
    port map (
            O => \N__9474\,
            I => \N__9448\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9448\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9445\
        );

    \I__1312\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9440\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9440\
        );

    \I__1310\ : InMux
    port map (
            O => \N__9469\,
            I => \N__9435\
        );

    \I__1309\ : InMux
    port map (
            O => \N__9466\,
            I => \N__9435\
        );

    \I__1308\ : InMux
    port map (
            O => \N__9465\,
            I => \N__9430\
        );

    \I__1307\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9430\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__9459\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__9456\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__9453\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__9448\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__9445\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__9440\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__9435\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__9430\,
            I => \this_vga_signals.M_vcounter_qZ0Z_8\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__9413\,
            I => \this_vga_signals.rgb297_i_a3_0_cascade_\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__1296\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9399\
        );

    \I__1295\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9396\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9405\,
            I => \N__9393\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9385\
        );

    \I__1292\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9385\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__9402\,
            I => \N__9382\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__9399\,
            I => \N__9375\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__9396\,
            I => \N__9372\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__9393\,
            I => \N__9369\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__9392\,
            I => \N__9366\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__9391\,
            I => \N__9361\
        );

    \I__1285\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9354\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9351\
        );

    \I__1283\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9344\
        );

    \I__1282\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9344\
        );

    \I__1281\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9344\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9339\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9339\
        );

    \I__1278\ : Span4Mux_v
    port map (
            O => \N__9375\,
            I => \N__9336\
        );

    \I__1277\ : Span4Mux_h
    port map (
            O => \N__9372\,
            I => \N__9331\
        );

    \I__1276\ : Span4Mux_h
    port map (
            O => \N__9369\,
            I => \N__9331\
        );

    \I__1275\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9324\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9324\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9324\
        );

    \I__1272\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9321\
        );

    \I__1271\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9312\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9312\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9312\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9312\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__9354\,
            I => \N__9309\
        );

    \I__1266\ : Span4Mux_h
    port map (
            O => \N__9351\,
            I => \N__9302\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__9344\,
            I => \N__9302\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9339\,
            I => \N__9302\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__9336\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__9331\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__9324\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9321\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__9312\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__9309\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__9302\,
            I => \this_vga_signals.M_vcounter_qZ0Z_6\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__9284\,
            I => \this_vga_signals.SUM_2_i_a4_0_a0_2_3\
        );

    \I__1254\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__1250\ : Span4Mux_h
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__9266\,
            I => \this_vga_signals.N_33_0\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9254\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9251\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9247\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9244\
        );

    \I__1244\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9241\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9236\
        );

    \I__1242\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9236\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__9254\,
            I => \N__9233\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9230\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__9250\,
            I => \N__9224\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9247\,
            I => \N__9220\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9244\,
            I => \N__9217\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__9241\,
            I => \N__9212\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__9236\,
            I => \N__9212\
        );

    \I__1234\ : Span4Mux_h
    port map (
            O => \N__9233\,
            I => \N__9208\
        );

    \I__1233\ : Span4Mux_h
    port map (
            O => \N__9230\,
            I => \N__9205\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9200\
        );

    \I__1231\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9200\
        );

    \I__1230\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9197\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9192\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9192\
        );

    \I__1227\ : Span4Mux_v
    port map (
            O => \N__9220\,
            I => \N__9185\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__9217\,
            I => \N__9185\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__9212\,
            I => \N__9185\
        );

    \I__1224\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9182\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__9208\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__9205\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__9200\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__9197\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__9192\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__9185\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__9182\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__1216\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9164\,
            I => \N__9160\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__1213\ : Odrv12
    port map (
            O => \N__9160\,
            I => \this_vga_signals.N_49\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__9157\,
            I => \this_vga_signals.N_49\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__9152\,
            I => \this_vga_signals.N_33_0_cascade_\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__9146\,
            I => \this_vga_signals.N_11_i\
        );

    \I__1208\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9139\
        );

    \I__1207\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9132\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__9139\,
            I => \N__9129\
        );

    \I__1205\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9122\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9122\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9122\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9119\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__9132\,
            I => \this_vga_signals.mult1_un40_sum_axb1\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__9129\,
            I => \this_vga_signals.mult1_un40_sum_axb1\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9122\,
            I => \this_vga_signals.mult1_un40_sum_axb1\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__9119\,
            I => \this_vga_signals.mult1_un40_sum_axb1\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9104\,
            I => \this_vga_signals.g0_5_0_0\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__9098\,
            I => \this_vga_signals.mult1_un54_sum_axb1_5_4\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__9095\,
            I => \this_vga_signals.g0_25_1_cascade_\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9086\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9083\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9078\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9078\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9086\,
            I => \N__9075\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9083\,
            I => \N__9072\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__9078\,
            I => \N__9069\
        );

    \I__1184\ : Span4Mux_v
    port map (
            O => \N__9075\,
            I => \N__9066\
        );

    \I__1183\ : Span4Mux_h
    port map (
            O => \N__9072\,
            I => \N__9063\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__9069\,
            I => \N__9060\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__9066\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__9063\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__9060\,
            I => \this_vga_signals.mult1_un47_sum_ac0_3_c\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__9053\,
            I => \this_vga_signals.if_N_13_i_i_1_0_0_cascade_\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9047\,
            I => \this_vga_signals.g2_0_0_0\
        );

    \I__1175\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__9035\,
            I => \this_vga_signals.N_371_0\
        );

    \I__1171\ : IoInMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__1169\ : Span12Mux_s11_h
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__1168\ : Odrv12
    port map (
            O => \N__9023\,
            I => rgb_c_4
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \N__9007\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9019\,
            I => \N__9004\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__9018\,
            I => \N__9001\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__9017\,
            I => \N__8997\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__9016\,
            I => \N__8994\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__9015\,
            I => \N__8991\
        );

    \I__1161\ : InMux
    port map (
            O => \N__9014\,
            I => \N__8987\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9013\,
            I => \N__8983\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8980\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8975\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9010\,
            I => \N__8975\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8972\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9004\,
            I => \N__8969\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8962\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8962\
        );

    \I__1152\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8962\
        );

    \I__1151\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8957\
        );

    \I__1150\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8957\
        );

    \I__1149\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8954\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8951\
        );

    \I__1147\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8948\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__8983\,
            I => \N__8945\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__8980\,
            I => \N__8936\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__8975\,
            I => \N__8936\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__8972\,
            I => \N__8936\
        );

    \I__1142\ : Span4Mux_h
    port map (
            O => \N__8969\,
            I => \N__8929\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__8962\,
            I => \N__8929\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__8957\,
            I => \N__8929\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__8954\,
            I => \N__8926\
        );

    \I__1138\ : Span4Mux_h
    port map (
            O => \N__8951\,
            I => \N__8919\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8919\
        );

    \I__1136\ : Span4Mux_v
    port map (
            O => \N__8945\,
            I => \N__8919\
        );

    \I__1135\ : InMux
    port map (
            O => \N__8944\,
            I => \N__8914\
        );

    \I__1134\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8914\
        );

    \I__1133\ : Span4Mux_h
    port map (
            O => \N__8936\,
            I => \N__8911\
        );

    \I__1132\ : Span4Mux_v
    port map (
            O => \N__8929\,
            I => \N__8908\
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__8926\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__8919\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__8914\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__8911\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__8908\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__8897\,
            I => \this_vga_signals.un11_address_0_7_cascade_\
        );

    \I__1125\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8888\
        );

    \I__1124\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8885\
        );

    \I__1123\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8880\
        );

    \I__1122\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8880\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__8888\,
            I => \N__8877\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__8885\,
            I => \this_vga_signals.SUM_2\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__8880\,
            I => \this_vga_signals.SUM_2\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__8877\,
            I => \this_vga_signals.SUM_2\
        );

    \I__1117\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__8867\,
            I => \N__8864\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__8864\,
            I => \this_vga_signals.g0_3_0\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__8861\,
            I => \this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_cascade_\
        );

    \I__1113\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__8855\,
            I => \this_vga_signals.g0_i_x2_1_1\
        );

    \I__1111\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__8849\,
            I => \this_vga_signals.g0_i_x1\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__8846\,
            I => \this_vga_signals.g0_i_x0_cascade_\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__8843\,
            I => \this_vga_signals_un16_address_if_i1_mux_0_cascade_\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__8840\,
            I => \this_vga_signals.N_6_i_cascade_\
        );

    \I__1106\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__8834\,
            I => \this_vga_signals.g1_1_0\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__8831\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIO6OD01Z0Z_9_cascade_\
        );

    \I__1103\ : IoInMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__8825\,
            I => \N__8822\
        );

    \I__1101\ : Span12Mux_s5_h
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__8819\,
            I => rgb_c_2
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__1098\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__8807\,
            I => \this_vga_signals.g0_i_x2_1_0\
        );

    \I__1095\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8801\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__8801\,
            I => \this_vga_signals.N_10_i\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__8798\,
            I => \this_vga_signals.N_10_i_cascade_\
        );

    \I__1092\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__8792\,
            I => \this_vga_signals.g0_i_x2_5_1\
        );

    \I__1090\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__8783\,
            I => \this_vga_signals.if_N_13_i_i_1\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__8780\,
            I => \this_vga_signals.g4_0_0_cascade_\
        );

    \I__1086\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__8774\,
            I => \N__8771\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__8771\,
            I => \this_vga_signals.g0_i_0_N_3L3\
        );

    \I__1083\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__8765\,
            I => \N__8762\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__8762\,
            I => \this_vga_signals.N_3_1_0_1\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__8759\,
            I => \this_vga_signals.g0_i_x2_1_1_cascade_\
        );

    \I__1079\ : InMux
    port map (
            O => \N__8756\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__1078\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8749\
        );

    \I__1077\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8746\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__8749\,
            I => \N__8740\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__8746\,
            I => \N__8740\
        );

    \I__1074\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8737\
        );

    \I__1073\ : Span4Mux_h
    port map (
            O => \N__8740\,
            I => \N__8734\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__8737\,
            I => \N__8731\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__8734\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__8731\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__1069\ : IoInMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1067\ : Span4Mux_s2_v
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__1066\ : Sp12to4
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__1065\ : Span12Mux_s10_h
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__1064\ : Odrv12
    port map (
            O => \N__8711\,
            I => \N_18\
        );

    \I__1063\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__8705\,
            I => \this_vga_signals.hsync_1_i_0_1\
        );

    \I__1061\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8697\
        );

    \I__1060\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8692\
        );

    \I__1059\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8692\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8697\,
            I => \N__8689\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__8692\,
            I => \N__8686\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__8689\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1055\ : Odrv12
    port map (
            O => \N__8686\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__1054\ : CEMux
    port map (
            O => \N__8681\,
            I => \N__8657\
        );

    \I__1053\ : CEMux
    port map (
            O => \N__8680\,
            I => \N__8657\
        );

    \I__1052\ : CEMux
    port map (
            O => \N__8679\,
            I => \N__8657\
        );

    \I__1051\ : CEMux
    port map (
            O => \N__8678\,
            I => \N__8657\
        );

    \I__1050\ : CEMux
    port map (
            O => \N__8677\,
            I => \N__8657\
        );

    \I__1049\ : CEMux
    port map (
            O => \N__8676\,
            I => \N__8657\
        );

    \I__1048\ : CEMux
    port map (
            O => \N__8675\,
            I => \N__8657\
        );

    \I__1047\ : CEMux
    port map (
            O => \N__8674\,
            I => \N__8657\
        );

    \I__1046\ : GlobalMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1045\ : gio2CtrlBuf
    port map (
            O => \N__8654\,
            I => \this_vga_signals.N_469_0_g\
        );

    \I__1044\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8636\
        );

    \I__1042\ : SRMux
    port map (
            O => \N__8647\,
            I => \N__8615\
        );

    \I__1041\ : SRMux
    port map (
            O => \N__8646\,
            I => \N__8615\
        );

    \I__1040\ : SRMux
    port map (
            O => \N__8645\,
            I => \N__8615\
        );

    \I__1039\ : SRMux
    port map (
            O => \N__8644\,
            I => \N__8615\
        );

    \I__1038\ : SRMux
    port map (
            O => \N__8643\,
            I => \N__8615\
        );

    \I__1037\ : SRMux
    port map (
            O => \N__8642\,
            I => \N__8615\
        );

    \I__1036\ : SRMux
    port map (
            O => \N__8641\,
            I => \N__8615\
        );

    \I__1035\ : SRMux
    port map (
            O => \N__8640\,
            I => \N__8615\
        );

    \I__1034\ : SRMux
    port map (
            O => \N__8639\,
            I => \N__8615\
        );

    \I__1033\ : Glb2LocalMux
    port map (
            O => \N__8636\,
            I => \N__8615\
        );

    \I__1032\ : GlobalMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1031\ : gio2CtrlBuf
    port map (
            O => \N__8612\,
            I => \this_vga_signals.N_608_g\
        );

    \I__1030\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__8606\,
            I => \this_vga_signals.N_381_0\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__8603\,
            I => \this_vga_signals.N_390_cascade_\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__8600\,
            I => \this_vga_signals.rgb_cnst_i_0_2_cascade_\
        );

    \I__1026\ : InMux
    port map (
            O => \N__8597\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__1025\ : InMux
    port map (
            O => \N__8594\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__1024\ : InMux
    port map (
            O => \N__8591\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8588\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8578\
        );

    \I__1020\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8575\
        );

    \I__1019\ : Span4Mux_h
    port map (
            O => \N__8578\,
            I => \N__8569\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8575\,
            I => \N__8569\
        );

    \I__1017\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8566\
        );

    \I__1016\ : Odrv4
    port map (
            O => \N__8569\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__8566\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__1014\ : InMux
    port map (
            O => \N__8561\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__1013\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__1011\ : Span12Mux_v
    port map (
            O => \N__8552\,
            I => \N__8547\
        );

    \I__1010\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8542\
        );

    \I__1009\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8542\
        );

    \I__1008\ : Odrv12
    port map (
            O => \N__8547\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__8542\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__1006\ : InMux
    port map (
            O => \N__8537\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8531\,
            I => \N__8526\
        );

    \I__1003\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8521\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8529\,
            I => \N__8521\
        );

    \I__1001\ : Odrv4
    port map (
            O => \N__8526\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__8521\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__999\ : InMux
    port map (
            O => \N__8516\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__998\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8509\
        );

    \I__997\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8506\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8502\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8499\
        );

    \I__994\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8496\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__8502\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__8499\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__8496\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__990\ : InMux
    port map (
            O => \N__8489\,
            I => \bfn_11_24_0_\
        );

    \I__989\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__8483\,
            I => \this_vga_signals.un11_address_c4_i\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__8480\,
            I => \this_vga_signals.SUM_2_i_a4_1_0_3_cascade_\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__8477\,
            I => \this_vga_signals.un11_address_c5_a0_0_cascade_\
        );

    \I__985\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8470\
        );

    \I__984\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8467\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__8470\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8467\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1\
        );

    \I__981\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8455\
        );

    \I__980\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8455\
        );

    \I__979\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8449\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__8455\,
            I => \N__8443\
        );

    \I__977\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8440\
        );

    \I__976\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8435\
        );

    \I__975\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8435\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__8449\,
            I => \N__8432\
        );

    \I__973\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8425\
        );

    \I__972\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8425\
        );

    \I__971\ : InMux
    port map (
            O => \N__8446\,
            I => \N__8425\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__8443\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8440\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__8435\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__8432\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__8425\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__8414\,
            I => \N__8406\
        );

    \I__964\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8401\
        );

    \I__963\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8401\
        );

    \I__962\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8396\
        );

    \I__961\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8396\
        );

    \I__960\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8391\
        );

    \I__959\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8391\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__8401\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__8396\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__8391\,
            I => \this_vga_signals.M_vcounter_q_9_repZ0Z1\
        );

    \I__955\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__8381\,
            I => \N__8375\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__8380\,
            I => \N__8372\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__8379\,
            I => \N__8368\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__8378\,
            I => \N__8364\
        );

    \I__950\ : Span4Mux_h
    port map (
            O => \N__8375\,
            I => \N__8359\
        );

    \I__949\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8356\
        );

    \I__948\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8353\
        );

    \I__947\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8346\
        );

    \I__946\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8346\
        );

    \I__945\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8346\
        );

    \I__944\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8343\
        );

    \I__943\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8340\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__8359\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__8356\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__8353\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8346\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8343\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__8340\,
            I => \this_vga_signals.M_vcounter_q_8_repZ0Z1\
        );

    \I__936\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8315\
        );

    \I__935\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8315\
        );

    \I__934\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8312\
        );

    \I__933\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8305\
        );

    \I__932\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8305\
        );

    \I__931\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8305\
        );

    \I__930\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8300\
        );

    \I__929\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8300\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__8315\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__8312\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__8305\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__8300\,
            I => \this_vga_signals.M_vcounter_q_7_repZ0Z1\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__8291\,
            I => \N__8285\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__8290\,
            I => \N__8277\
        );

    \I__922\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8274\
        );

    \I__921\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8271\
        );

    \I__920\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8268\
        );

    \I__919\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8263\
        );

    \I__918\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8263\
        );

    \I__917\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8258\
        );

    \I__916\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8258\
        );

    \I__915\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8253\
        );

    \I__914\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8253\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__8274\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__8271\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8268\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__8263\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__8258\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__8253\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__907\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8230\
        );

    \I__906\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8230\
        );

    \I__905\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8230\
        );

    \I__904\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8225\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8230\,
            I => \N__8215\
        );

    \I__902\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8210\
        );

    \I__901\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8210\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8225\,
            I => \N__8207\
        );

    \I__899\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8198\
        );

    \I__898\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8198\
        );

    \I__897\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8198\
        );

    \I__896\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8198\
        );

    \I__895\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8193\
        );

    \I__894\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8193\
        );

    \I__893\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8190\
        );

    \I__892\ : Span4Mux_v
    port map (
            O => \N__8215\,
            I => \N__8185\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__8210\,
            I => \N__8185\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__8207\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__8198\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8193\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__8190\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__8185\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__8174\,
            I => \this_vga_signals.SUM_2_i_a4_0_a0_2_3_cascade_\
        );

    \I__884\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__8168\,
            I => \this_vga_signals.SUM_2_i_a4_a0_2_3\
        );

    \I__882\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8162\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8162\,
            I => \this_vga_signals.SUM_2_i_1_0_3\
        );

    \I__880\ : InMux
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__8156\,
            I => \this_vga_signals.SUM_2_i_0_1_3\
        );

    \I__878\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8150\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__8150\,
            I => \this_vga_signals.SUM_2_i_0_3\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__8147\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\
        );

    \I__875\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__8141\,
            I => \N__8138\
        );

    \I__873\ : Span4Mux_h
    port map (
            O => \N__8138\,
            I => \N__8135\
        );

    \I__872\ : Odrv4
    port map (
            O => \N__8135\,
            I => \this_vga_signals.g0_1\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__8132\,
            I => \this_vga_signals.un11_address_c4_i_cascade_\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__8129\,
            I => \this_vga_signals.mult1_un54_sum_axb1_5_4_1_cascade_\
        );

    \I__869\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8120\
        );

    \I__868\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8120\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8120\,
            I => \N__8116\
        );

    \I__866\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8113\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__8116\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__8113\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__8108\,
            I => \this_vga_signals.mult1_un54_sum_axb1_5_4_cascade_\
        );

    \I__862\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8095\
        );

    \I__861\ : InMux
    port map (
            O => \N__8104\,
            I => \N__8095\
        );

    \I__860\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8095\
        );

    \I__859\ : InMux
    port map (
            O => \N__8102\,
            I => \N__8092\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8095\,
            I => \N__8087\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__8092\,
            I => \N__8084\
        );

    \I__856\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8081\
        );

    \I__855\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8078\
        );

    \I__854\ : Span4Mux_h
    port map (
            O => \N__8087\,
            I => \N__8075\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__8084\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8081\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8078\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__8075\,
            I => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0\
        );

    \I__849\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8058\
        );

    \I__848\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8058\
        );

    \I__847\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8053\
        );

    \I__846\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8053\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8058\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__8053\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__8048\,
            I => \N__8043\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__8047\,
            I => \N__8040\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__8046\,
            I => \N__8037\
        );

    \I__840\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8034\
        );

    \I__839\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8029\
        );

    \I__838\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8029\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8034\,
            I => \N__8026\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8029\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__8026\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__834\ : InMux
    port map (
            O => \N__8021\,
            I => \N__8016\
        );

    \I__833\ : InMux
    port map (
            O => \N__8020\,
            I => \N__8011\
        );

    \I__832\ : InMux
    port map (
            O => \N__8019\,
            I => \N__8011\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8016\,
            I => \N__8008\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8011\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__8008\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__828\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7998\
        );

    \I__827\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7995\
        );

    \I__826\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7992\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__7998\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__7995\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__7992\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__7985\,
            I => \N__7981\
        );

    \I__821\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7976\
        );

    \I__820\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7976\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__818\ : Span4Mux_h
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__7970\,
            I => \this_vga_signals.if_N_3_0_i\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__7967\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_c_cascade_\
        );

    \I__815\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7958\
        );

    \I__814\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7953\
        );

    \I__813\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7953\
        );

    \I__812\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7950\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__7958\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__7953\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__7950\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1\
        );

    \I__808\ : InMux
    port map (
            O => \N__7943\,
            I => \N__7937\
        );

    \I__807\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7937\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__7937\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_c\
        );

    \I__805\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__7925\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1_0\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__800\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__798\ : Span4Mux_h
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__797\ : Odrv4
    port map (
            O => \N__7910\,
            I => \this_vga_signals.if_N_3_0_i_0\
        );

    \I__796\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7903\
        );

    \I__795\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7900\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__7903\,
            I => \N__7895\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__7900\,
            I => \N__7891\
        );

    \I__792\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7888\
        );

    \I__791\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7884\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__7895\,
            I => \N__7879\
        );

    \I__789\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7876\
        );

    \I__788\ : Span4Mux_h
    port map (
            O => \N__7891\,
            I => \N__7873\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__7888\,
            I => \N__7870\
        );

    \I__786\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7867\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__7884\,
            I => \N__7864\
        );

    \I__784\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7859\
        );

    \I__783\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7859\
        );

    \I__782\ : Odrv4
    port map (
            O => \N__7879\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__7876\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__7873\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__7870\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__7867\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__777\ : Odrv4
    port map (
            O => \N__7864\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__7859\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1\
        );

    \I__775\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7838\
        );

    \I__774\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7835\
        );

    \I__773\ : InMux
    port map (
            O => \N__7842\,
            I => \N__7827\
        );

    \I__772\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7824\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__7838\,
            I => \N__7821\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__7835\,
            I => \N__7818\
        );

    \I__769\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7815\
        );

    \I__768\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7810\
        );

    \I__767\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7810\
        );

    \I__766\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7805\
        );

    \I__765\ : InMux
    port map (
            O => \N__7830\,
            I => \N__7805\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__7827\,
            I => \N__7802\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__7824\,
            I => \N__7799\
        );

    \I__762\ : Span4Mux_h
    port map (
            O => \N__7821\,
            I => \N__7791\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__7818\,
            I => \N__7791\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__7815\,
            I => \N__7791\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__7810\,
            I => \N__7788\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7781\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__7802\,
            I => \N__7781\
        );

    \I__756\ : Span4Mux_h
    port map (
            O => \N__7799\,
            I => \N__7781\
        );

    \I__755\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7778\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__7791\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2\
        );

    \I__753\ : Odrv12
    port map (
            O => \N__7788\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__7781\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__7778\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2\
        );

    \I__750\ : InMux
    port map (
            O => \N__7769\,
            I => \N__7766\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__7766\,
            I => \N__7762\
        );

    \I__748\ : InMux
    port map (
            O => \N__7765\,
            I => \N__7759\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__7762\,
            I => \this_vga_signals.mult1_un54_sum_axb2_0\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__7759\,
            I => \this_vga_signals.mult1_un54_sum_axb2_0\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__7754\,
            I => \this_vga_signals.mult1_un40_sum_axb1_cascade_\
        );

    \I__744\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7747\
        );

    \I__743\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7744\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__7747\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_0\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__7744\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_0\
        );

    \I__740\ : InMux
    port map (
            O => \N__7739\,
            I => \N__7736\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__7733\,
            I => \this_vga_signals.g0_5_1\
        );

    \I__737\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7724\
        );

    \I__736\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7724\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__7724\,
            I => \N__7720\
        );

    \I__734\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7717\
        );

    \I__733\ : Odrv4
    port map (
            O => \N__7720\,
            I => \this_vga_signals.mult1_un47_sum_c2_0\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__7717\,
            I => \this_vga_signals.mult1_un47_sum_c2_0\
        );

    \I__731\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7709\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__7709\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_x1\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__7706\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_x0_cascade_\
        );

    \I__728\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__7700\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__7697\,
            I => \this_vga_signals.mult1_un54_sum_i_1_cascade_\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__7694\,
            I => \this_vga_signals.un11_address_2_5_cascade_\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__7691\,
            I => \this_vga_signals.mult1_un54_sum_i_x0_3_cascade_\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__722\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7681\
        );

    \I__721\ : InMux
    port map (
            O => \N__7684\,
            I => \N__7678\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__7681\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__7678\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__718\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7669\
        );

    \I__717\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7666\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__7669\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__7666\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__714\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7655\
        );

    \I__713\ : InMux
    port map (
            O => \N__7660\,
            I => \N__7655\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__7655\,
            I => \N__7651\
        );

    \I__711\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7648\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__7651\,
            I => \N__7645\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__7648\,
            I => \N__7642\
        );

    \I__708\ : Odrv4
    port map (
            O => \N__7645\,
            I => \this_vga_signals.d_N_8_0\
        );

    \I__707\ : Odrv12
    port map (
            O => \N__7642\,
            I => \this_vga_signals.d_N_8_0\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__7637\,
            I => \this_vga_signals.un11_address_1_5_cascade_\
        );

    \I__705\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__7631\,
            I => \this_vga_signals.g0_11_1\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__702\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7622\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__7622\,
            I => \this_vga_signals.g0_6_0\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__7619\,
            I => \this_vga_signals.g2_1_0_cascade_\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__7616\,
            I => \this_vga_signals.g3_cascade_\
        );

    \I__698\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__7610\,
            I => \this_vga_signals.g2_4_0\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__7607\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_2_N_2L1_cascade_\
        );

    \I__695\ : InMux
    port map (
            O => \N__7604\,
            I => \N__7598\
        );

    \I__694\ : InMux
    port map (
            O => \N__7603\,
            I => \N__7598\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__7598\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__692\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7592\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__7586\,
            I => \this_vga_signals.un11_address_0_5\
        );

    \I__688\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__686\ : Odrv4
    port map (
            O => \N__7577\,
            I => \this_vga_signals.vsync_1_0_a3_4\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__684\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__7565\,
            I => \this_vga_signals.if_N_15_mux\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__7562\,
            I => \this_vga_signals.if_m13_ns_1_cascade_\
        );

    \I__680\ : InMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__7556\,
            I => \N__7552\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__7555\,
            I => \N__7549\
        );

    \I__677\ : Span4Mux_h
    port map (
            O => \N__7552\,
            I => \N__7545\
        );

    \I__676\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7540\
        );

    \I__675\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7540\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__7545\,
            I => \this_vga_signals.if_m13_ns\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__7540\,
            I => \this_vga_signals.if_m13_ns\
        );

    \I__672\ : InMux
    port map (
            O => \N__7535\,
            I => \N__7532\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__7532\,
            I => \this_vga_signals.if_N_7\
        );

    \I__670\ : InMux
    port map (
            O => \N__7529\,
            I => \N__7526\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7526\,
            I => \this_vga_signals.d_N_9_0\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__7523\,
            I => \this_vga_signals.rgb_1_4_cascade_\
        );

    \I__667\ : InMux
    port map (
            O => \N__7520\,
            I => \N__7516\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__7519\,
            I => \N__7513\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__7516\,
            I => \N__7509\
        );

    \I__664\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7504\
        );

    \I__663\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7504\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__7509\,
            I => \N__7499\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__7504\,
            I => \N__7499\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__7499\,
            I => \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIETZ0Z844\
        );

    \I__659\ : InMux
    port map (
            O => \N__7496\,
            I => \N__7493\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__7493\,
            I => \this_vga_signals.d_N_5_0\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__656\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__7481\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__7478\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__651\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__7469\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_i_x1\
        );

    \I__649\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__7460\,
            I => \this_vga_signals.g1\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__7457\,
            I => \this_vga_signals.g3_0_2_cascade_\
        );

    \I__645\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__7451\,
            I => \this_vga_signals.if_N_3_0_i_1\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__7448\,
            I => \this_vga_signals.mult1_un54_sum_ac0_3_c_0_cascade_\
        );

    \I__642\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__7442\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_1\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__7439\,
            I => \this_vga_signals.mult1_un47_sum_ac0_1_cascade_\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__7436\,
            I => \this_vga_signals.rgb_1_2_cascade_\
        );

    \I__638\ : InMux
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__7427\,
            I => \this_vga_signals.if_i3_mux_0_0\
        );

    \I__635\ : InMux
    port map (
            O => \N__7424\,
            I => \N__7420\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__7423\,
            I => \N__7417\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__7420\,
            I => \N__7414\
        );

    \I__632\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7411\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__7414\,
            I => \this_vga_signals.if_i3_mux_2\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__7411\,
            I => \this_vga_signals.if_i3_mux_2\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__7406\,
            I => \this_vga_signals.g2_1_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__7400\,
            I => \this_vga_signals.g2_1\
        );

    \I__626\ : InMux
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__7394\,
            I => \this_vga_signals.mult1_un54_sum_ac0_1_1_0\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__7391\,
            I => \N__7388\
        );

    \I__623\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7385\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__7385\,
            I => \this_vga_signals.g0_5_0_1\
        );

    \I__621\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__7379\,
            I => \this_vga_signals.g3_0_2_0\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__7376\,
            I => \this_vga_signals.g2_cascade_\
        );

    \I__618\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7370\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__7370\,
            I => \this_vga_signals.g0_3_0_0\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__7367\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_2_0_cascade_\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__614\ : InMux
    port map (
            O => \N__7361\,
            I => \N__7358\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__7358\,
            I => \this_vga_signals.if_m1_3\
        );

    \I__612\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7352\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__7352\,
            I => \this_vga_signals.if_N_4_2\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__7349\,
            I => \this_vga_signals.if_i4_mux_0_1_cascade_\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__7346\,
            I => \this_vga_signals.vsync_1_0_a3_5_cascade_\
        );

    \I__608\ : IoInMux
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__606\ : Span12Mux_s10_v
    port map (
            O => \N__7337\,
            I => \N__7334\
        );

    \I__605\ : Odrv12
    port map (
            O => \N__7334\,
            I => this_vga_signals_vsync_1_i
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__7331\,
            I => \this_vga_signals.if_m13_0_ns_1_cascade_\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__7328\,
            I => \this_vga_signals.if_i3_mux_0_0_cascade_\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__7325\,
            I => \N__7322\
        );

    \I__601\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7319\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__7319\,
            I => \this_vga_signals.if_m13_0_ns_1\
        );

    \I__599\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7313\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__597\ : Odrv12
    port map (
            O => \N__7310\,
            I => \this_vga_signals.if_i3_mux_0_0_0\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__7307\,
            I => \this_vga_signals.if_m8_0_ns_1_cascade_\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__7304\,
            I => \this_vga_signals.g1_1_cascade_\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__7301\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__7298\,
            I => \this_vga_signals.g1_cascade_\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__7295\,
            I => \this_vga_signals.if_m1_3_cascade_\
        );

    \I__591\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7280\
        );

    \I__590\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7280\
        );

    \I__589\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7280\
        );

    \I__588\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7280\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__7274\,
            I => \N__7271\
        );

    \I__584\ : Span12Mux_h
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__583\ : Span12Mux_v
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__582\ : Odrv12
    port map (
            O => \N__7265\,
            I => rst_n_c
        );

    \I__581\ : InMux
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__7259\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__7256\,
            I => \this_vga_signals.if_i3_mux_2_0_cascade_\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__7253\,
            I => \this_vga_signals.if_m2_8_0_cascade_\
        );

    \I__577\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__7247\,
            I => \this_vga_signals.if_m8_0_ns_1\
        );

    \I__575\ : InMux
    port map (
            O => \N__7244\,
            I => \N__7241\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__7241\,
            I => \this_vga_signals.rgb_cnst_i_1Z0Z_5\
        );

    \I__573\ : IoInMux
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__571\ : Span4Mux_s1_h
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__570\ : Span4Mux_h
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__569\ : Span4Mux_v
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__7223\,
            I => rgb_c_5
        );

    \I__567\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7217\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__7217\,
            I => \N__7214\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__7214\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIAV48E1Z0Z_9\
        );

    \I__564\ : IoInMux
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__562\ : IoSpan4Mux
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__561\ : IoSpan4Mux
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__560\ : Span4Mux_s2_h
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__7196\,
            I => rgb_c_3
        );

    \I__558\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7189\
        );

    \I__557\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7186\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__7189\,
            I => \this_vga_signals.N_379_0\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__7186\,
            I => \this_vga_signals.N_379_0\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__7181\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIA99QRZ0Z_9_cascade_\
        );

    \I__553\ : IoInMux
    port map (
            O => \N__7178\,
            I => \N__7175\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__7175\,
            I => \N__7172\
        );

    \I__551\ : Span4Mux_s3_h
    port map (
            O => \N__7172\,
            I => \N__7169\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__7169\,
            I => rgb_c_1
        );

    \I__549\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__7163\,
            I => \this_vga_signals.rgb_cnst_i_0_5\
        );

    \I__547\ : IoInMux
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__7157\,
            I => \N__7153\
        );

    \I__545\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7150\
        );

    \I__544\ : IoSpan4Mux
    port map (
            O => \N__7153\,
            I => \N__7147\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__7150\,
            I => \N__7144\
        );

    \I__542\ : Sp12to4
    port map (
            O => \N__7147\,
            I => \N__7141\
        );

    \I__541\ : Span4Mux_v
    port map (
            O => \N__7144\,
            I => \N__7138\
        );

    \I__540\ : Span12Mux_s6_h
    port map (
            O => \N__7141\,
            I => \N__7135\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__7138\,
            I => \N__7132\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__7135\,
            I => \N_11_0\
        );

    \I__537\ : Odrv4
    port map (
            O => \N__7132\,
            I => \N_11_0\
        );

    \I__536\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7124\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__7124\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__534\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7118\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__7118\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__532\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7112\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__7112\,
            I => \N__7109\
        );

    \I__530\ : Odrv4
    port map (
            O => \N__7109\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \I__529\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__7103\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__527\ : IoInMux
    port map (
            O => \N__7100\,
            I => \N__7097\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__525\ : Odrv12
    port map (
            O => \N__7094\,
            I => \N_33\
        );

    \I__524\ : IoInMux
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__522\ : Odrv12
    port map (
            O => \N__7085\,
            I => \N_11\
        );

    \I__521\ : IoInMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__519\ : Span4Mux_s1_h
    port map (
            O => \N__7076\,
            I => \N__7073\
        );

    \I__518\ : Span4Mux_v
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__517\ : Span4Mux_v
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__516\ : Span4Mux_h
    port map (
            O => \N__7067\,
            I => \N__7064\
        );

    \I__515\ : Odrv4
    port map (
            O => \N__7064\,
            I => rgb_c_0
        );

    \I__514\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7058\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__7058\,
            I => \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1Z0Z_9\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__7055\,
            I => \this_vga_signals.rgb_cnst_i_1Z0Z_3_cascade_\
        );

    \I__511\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__7049\,
            I => port_clk_c
        );

    \I__509\ : IoInMux
    port map (
            O => \N__7046\,
            I => \N__7043\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__507\ : Span4Mux_s0_h
    port map (
            O => \N__7040\,
            I => \N__7037\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__7037\,
            I => \this_vga_signals.N_469_0\
        );

    \I__505\ : IoInMux
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__7031\,
            I => port_rw_c_i
        );

    \I__503\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__7025\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \IN_MUX_bfv_12_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_24_0_\
        );

    \IN_MUX_bfv_12_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_12_25_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_current_address_q_cry_7\,
            carryinitout => \bfn_15_22_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIVV6F6_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9515\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_608_g\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIR7M7_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7046\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_469_0_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7052\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIR7M7_9_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11706\,
            in2 => \_gnd_net_\,
            in3 => \N__8651\,
            lcout => \this_vga_signals.N_469_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_rw_obuf_RNO_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => port_rw_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7106\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7028\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7115\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_0_9_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9281\,
            lcout => \N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIEC104_0_9_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7156\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI18GF6U3_9_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14091\,
            in1 => \N__7061\,
            in2 => \_gnd_net_\,
            in3 => \N__12926\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1_9_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000000000"
        )
    port map (
            in0 => \N__10413\,
            in1 => \N__13774\,
            in2 => \N__12988\,
            in3 => \N__20309\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_cnst_i_1_3_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011101111"
        )
    port map (
            in0 => \N__15904\,
            in1 => \N__10420\,
            in2 => \N__13787\,
            in3 => \N__13007\,
            lcout => OPEN,
            ltout => \this_vga_signals.rgb_cnst_i_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIAV48E1_9_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001000000"
        )
    port map (
            in0 => \N__10436\,
            in1 => \N__7192\,
            in2 => \N__7055\,
            in3 => \N__13775\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNIAV48E1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGGSVD_9_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__13008\,
            in1 => \N__13788\,
            in2 => \_gnd_net_\,
            in3 => \N__20331\,
            lcout => \this_vga_signals.N_379_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_cnst_i_1_5_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101111001111"
        )
    port map (
            in0 => \N__10421\,
            in1 => \N__15905\,
            in2 => \N__13793\,
            in3 => \N__13009\,
            lcout => \this_vga_signals.rgb_cnst_i_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI9UBTOU3_9_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__7244\,
            in1 => \N__14092\,
            in2 => \N__14849\,
            in3 => \N__7166\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIDP942V3_9_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14093\,
            in1 => \N__7220\,
            in2 => \_gnd_net_\,
            in3 => \N__13055\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIA99QR_9_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000010"
        )
    port map (
            in0 => \N__7193\,
            in1 => \N__10411\,
            in2 => \N__13010\,
            in3 => \N__15903\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_esr_RNIA99QRZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNID3EMFU3_9_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14084\,
            in2 => \N__7181\,
            in3 => \N__11540\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_9_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__10412\,
            in1 => \N__13006\,
            in2 => \N__13792\,
            in3 => \N__20330\,
            lcout => \this_vga_signals.rgb_cnst_i_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7289\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIEC104_9_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9167\,
            in1 => \N__9593\,
            in2 => \_gnd_net_\,
            in3 => \N__9260\,
            lcout => \N_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__7290\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7127\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7291\,
            in2 => \_gnd_net_\,
            in3 => \N__7121\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__7292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7262\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_3_1_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010010100101"
        )
    port map (
            in0 => \N__9821\,
            in1 => \N__7559\,
            in2 => \N__11464\,
            in3 => \N__7520\,
            lcout => \this_vga_signals.g0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_26_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__9365\,
            in1 => \N__7250\,
            in2 => \_gnd_net_\,
            in3 => \N__9794\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_i3_mux_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_24_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110000"
        )
    port map (
            in0 => \N__7316\,
            in1 => \N__8240\,
            in2 => \N__7256\,
            in3 => \N__18342\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_5_2_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011010"
        )
    port map (
            in0 => \N__8239\,
            in1 => \_gnd_net_\,
            in2 => \N__9392\,
            in3 => \N__9795\,
            lcout => \this_vga_signals.g0_5_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m2_8_0_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101100110"
        )
    port map (
            in0 => \N__9793\,
            in1 => \N__9364\,
            in2 => \_gnd_net_\,
            in3 => \N__8238\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m2_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m2_8_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7887\,
            in2 => \N__7253\,
            in3 => \N__7841\,
            lcout => \this_vga_signals.if_N_3_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8585\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18212\,
            ce => \N__8674\,
            sr => \N__8647\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8558\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18212\,
            ce => \N__8674\,
            sr => \N__8647\
        );

    \this_vga_signals.un16_address_if_m8_0_ns_1_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101100100100"
        )
    port map (
            in0 => \N__9740\,
            in1 => \N__9357\,
            in2 => \N__9250\,
            in3 => \N__9472\,
            lcout => \this_vga_signals.if_m8_0_ns_1\,
            ltout => \this_vga_signals.if_m8_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m8_0_ns_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001011010"
        )
    port map (
            in0 => \N__9358\,
            in1 => \_gnd_net_\,
            in2 => \N__7307\,
            in3 => \N__9832\,
            lcout => \this_vga_signals.if_i3_mux_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g1_1_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9833\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11426\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_14_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110100101"
        )
    port map (
            in0 => \N__9359\,
            in1 => \N__7894\,
            in2 => \N__7304\,
            in3 => \N__7831\,
            lcout => \this_vga_signals.if_N_3_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_1_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100011101"
        )
    port map (
            in0 => \N__8384\,
            in1 => \N__9223\,
            in2 => \N__7490\,
            in3 => \N__9739\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1\,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g1_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__7830\,
            in1 => \_gnd_net_\,
            in2 => \N__7301\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.g1\,
            ltout => \this_vga_signals.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_22_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__9360\,
            in1 => \N__11427\,
            in2 => \N__7298\,
            in3 => \N__9834\,
            lcout => \this_vga_signals.if_N_3_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m1_3_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__9379\,
            in1 => \N__8229\,
            in2 => \_gnd_net_\,
            in3 => \N__8284\,
            lcout => \this_vga_signals.if_m1_3\,
            ltout => \this_vga_signals.if_m1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m3_1_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__9727\,
            in1 => \_gnd_net_\,
            in2 => \N__7295\,
            in3 => \N__9228\,
            lcout => \this_vga_signals.if_N_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__9378\,
            in1 => \N__8228\,
            in2 => \_gnd_net_\,
            in3 => \N__8283\,
            lcout => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m7_1_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000001"
        )
    port map (
            in0 => \N__9728\,
            in1 => \N__9473\,
            in2 => \N__7364\,
            in3 => \N__9229\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_i4_mux_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m8_1_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011100100"
        )
    port map (
            in0 => \N__9474\,
            in1 => \N__7355\,
            in2 => \N__7349\,
            in3 => \N__18297\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8753\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18220\,
            ce => \N__8675\,
            sr => \N__8646\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI2GCG1_7_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11395\,
            in1 => \N__12169\,
            in2 => \N__9402\,
            in3 => \N__9711\,
            lcout => OPEN,
            ltout => \this_vga_signals.vsync_1_0_a3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7583\,
            in1 => \N__9471\,
            in2 => \N__7346\,
            in3 => \N__12476\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m13_0_ns_1_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9470\,
            in1 => \N__9227\,
            in2 => \_gnd_net_\,
            in3 => \N__9710\,
            lcout => \this_vga_signals.if_m13_0_ns_1\,
            ltout => \this_vga_signals.if_m13_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m13_0_ns_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110101100101"
        )
    port map (
            in0 => \N__9830\,
            in1 => \N__9380\,
            in2 => \N__7331\,
            in3 => \N__7660\,
            lcout => \this_vga_signals.if_i3_mux_0_0\,
            ltout => \this_vga_signals.if_i3_mux_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_15_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101000100"
        )
    port map (
            in0 => \N__11394\,
            in1 => \N__7424\,
            in2 => \N__7328\,
            in3 => \N__18322\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_34_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110101100101"
        )
    port map (
            in0 => \N__9831\,
            in1 => \N__9381\,
            in2 => \N__7325\,
            in3 => \N__7661\,
            lcout => \this_vga_signals.if_i3_mux_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m11_1_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__7673\,
            in1 => \N__8371\,
            in2 => \N__7688\,
            in3 => \N__8454\,
            lcout => \this_vga_signals.if_N_15_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_9_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8745\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18227\,
            ce => \N__8680\,
            sr => \N__8642\
        );

    \this_vga_signals.un16_address_g2_3_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7899\,
            in2 => \_gnd_net_\,
            in3 => \N__7842\,
            lcout => \this_vga_signals.g2_1\,
            ltout => \this_vga_signals.g2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g3_0_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11409\,
            in1 => \N__9852\,
            in2 => \N__7406\,
            in3 => \N__8990\,
            lcout => \this_vga_signals.g3_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001111011"
        )
    port map (
            in0 => \N__7403\,
            in1 => \N__7397\,
            in2 => \N__7391\,
            in3 => \N__17321\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_13_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000011110000"
        )
    port map (
            in0 => \N__17322\,
            in1 => \N__7382\,
            in2 => \N__7376\,
            in3 => \N__7373\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_12_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17111\,
            in1 => \N__8144\,
            in2 => \N__7367\,
            in3 => \N__11146\,
            lcout => \this_vga_signals.N_3_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_0_N_3L3_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12330\,
            in2 => \N__17160\,
            in3 => \N__11145\,
            lcout => \this_vga_signals.g0_i_0_N_3L3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x2_2_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101011010"
        )
    port map (
            in0 => \N__11512\,
            in1 => \N__12516\,
            in2 => \N__11456\,
            in3 => \N__12552\,
            lcout => \this_vga_signals.g0_i_x2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g4_0_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__11417\,
            in1 => \N__7445\,
            in2 => \N__12363\,
            in3 => \N__10901\,
            lcout => \this_vga_signals.g4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_5_1_0_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000101010101"
        )
    port map (
            in0 => \N__9090\,
            in1 => \N__9138\,
            in2 => \N__9018\,
            in3 => \N__18341\,
            lcout => \this_vga_signals.g0_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_c2_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111110101"
        )
    port map (
            in0 => \N__8103\,
            in1 => \N__7882\,
            in2 => \N__9015\,
            in3 => \N__7832\,
            lcout => \this_vga_signals.mult1_un47_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_0_0_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000101010101"
        )
    port map (
            in0 => \N__9089\,
            in1 => \N__9136\,
            in2 => \N__9017\,
            in3 => \N__18340\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_c2_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__8105\,
            in1 => \N__7961\,
            in2 => \_gnd_net_\,
            in3 => \N__8001\,
            lcout => \this_vga_signals.mult1_un54_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_1_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000001010"
        )
    port map (
            in0 => \N__8104\,
            in1 => \N__7883\,
            in2 => \N__9016\,
            in3 => \N__7833\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un47_sum_ac0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_ac0_3_d_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__9000\,
            in1 => \N__9137\,
            in2 => \N__7439\,
            in3 => \N__18339\,
            lcout => \this_vga_signals.mult1_un47_sum_ac0_3_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_i_3_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__8222\,
            in1 => \N__9790\,
            in2 => \N__7555\,
            in3 => \N__7512\,
            lcout => \this_vga_signals.rgb_1_2\,
            ltout => \this_vga_signals.rgb_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18336\,
            in1 => \N__8943\,
            in2 => \N__7436\,
            in3 => \N__7723\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__8224\,
            in1 => \N__7433\,
            in2 => \N__7423\,
            in3 => \N__18335\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g3_0_2_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9792\,
            in1 => \N__7466\,
            in2 => \N__11463\,
            in3 => \N__8944\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_19_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__7595\,
            in1 => \N__8003\,
            in2 => \N__7457\,
            in3 => \N__17310\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_3_c_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_18_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001101"
        )
    port map (
            in0 => \N__17311\,
            in1 => \N__7454\,
            in2 => \N__7448\,
            in3 => \N__7964\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABC21_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000111"
        )
    port map (
            in0 => \N__8221\,
            in1 => \N__8289\,
            in2 => \N__9391\,
            in3 => \N__9732\,
            lcout => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIABCZ0Z21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un47_sum_axbxc3_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000111"
        )
    port map (
            in0 => \N__9791\,
            in1 => \N__7548\,
            in2 => \N__7519\,
            in3 => \N__8223\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIG8C01_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100001100000"
        )
    port map (
            in0 => \N__8412\,
            in1 => \N__8326\,
            in2 => \N__9485\,
            in3 => \N__8461\,
            lcout => \this_vga_signals.d_N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8513\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18213\,
            ce => \N__8676\,
            sr => \N__8645\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8581\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18213\,
            ce => \N__8676\,
            sr => \N__8645\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8534\,
            lcout => \this_vga_signals.M_vcounter_q_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18213\,
            ce => \N__8676\,
            sr => \N__8645\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8752\,
            lcout => \this_vga_signals.M_vcounter_q_9_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18213\,
            ce => \N__8676\,
            sr => \N__8645\
        );

    \this_vga_signals.un16_address_if_m13_ns_1_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101110111"
        )
    port map (
            in0 => \N__8462\,
            in1 => \N__7654\,
            in2 => \N__7574\,
            in3 => \N__8288\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m13_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m13_ns_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101000100"
        )
    port map (
            in0 => \N__9390\,
            in1 => \N__7535\,
            in2 => \N__7562\,
            in3 => \N__18296\,
            lcout => \this_vga_signals.if_m13_ns\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m6_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100110010011"
        )
    port map (
            in0 => \N__8327\,
            in1 => \N__9469\,
            in2 => \N__8291\,
            in3 => \N__8413\,
            lcout => \this_vga_signals.if_N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_ns_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14337\,
            in2 => \N__7475\,
            in3 => \N__7798\,
            lcout => \this_vga_signals.rgb_1_4\,
            ltout => \this_vga_signals.rgb_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIET844_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7529\,
            in2 => \N__7523\,
            in3 => \N__7496\,
            lcout => \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIETZ0Z844\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111111"
        )
    port map (
            in0 => \N__8321\,
            in1 => \N__8411\,
            in2 => \N__8380\,
            in3 => \N__8453\,
            lcout => \this_vga_signals.d_N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_0_2_1_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8064\,
            in1 => \N__7604\,
            in2 => \N__8047\,
            in3 => \N__8020\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1\,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_i_x1_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011100100"
        )
    port map (
            in0 => \N__9211\,
            in1 => \N__8362\,
            in2 => \N__7478\,
            in3 => \N__9697\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_i_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_N_2L1_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__8063\,
            in1 => \N__7603\,
            in2 => \N__8046\,
            in3 => \N__8019\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_2_N_2L1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_ac0_3_2_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110001111"
        )
    port map (
            in0 => \N__8320\,
            in1 => \N__8410\,
            in2 => \N__7607\,
            in3 => \N__8452\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8512\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18215\,
            ce => \N__8677\,
            sr => \N__8643\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8574\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18221\,
            ce => \N__8679\,
            sr => \N__8641\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18221\,
            ce => \N__8679\,
            sr => \N__8641\
        );

    \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8505\,
            lcout => \this_vga_signals.M_vcounter_q_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18221\,
            ce => \N__8679\,
            sr => \N__8641\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8550\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18221\,
            ce => \N__8679\,
            sr => \N__8641\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8551\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18221\,
            ce => \N__8679\,
            sr => \N__8641\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8529\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18221\,
            ce => \N__8679\,
            sr => \N__8641\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_5_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11270\,
            in2 => \_gnd_net_\,
            in3 => \N__9874\,
            lcout => \this_vga_signals.un11_address_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIA9V41_9_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9261\,
            in1 => \N__12258\,
            in2 => \_gnd_net_\,
            in3 => \N__9875\,
            lcout => \this_vga_signals.vsync_1_0_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNII2LG_7_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__7684\,
            in1 => \N__7672\,
            in2 => \_gnd_net_\,
            in3 => \N__8363\,
            lcout => \this_vga_signals.d_N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_11_1_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__9860\,
            in1 => \N__9406\,
            in2 => \N__11460\,
            in3 => \N__9143\,
            lcout => \this_vga_signals.g0_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_11_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20323\,
            in2 => \_gnd_net_\,
            in3 => \N__17168\,
            lcout => this_vram_mem_radreg_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18196\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNILIQM_0_5_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11428\,
            in2 => \_gnd_net_\,
            in3 => \N__9859\,
            lcout => OPEN,
            ltout => \this_vga_signals.un11_address_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_6_0_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001010000"
        )
    port map (
            in0 => \N__9019\,
            in1 => \N__7907\,
            in2 => \N__7637\,
            in3 => \N__7843\,
            lcout => \this_vga_signals.g0_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_11_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011100"
        )
    port map (
            in0 => \N__7634\,
            in1 => \N__9092\,
            in2 => \N__7628\,
            in3 => \N__18358\,
            lcout => OPEN,
            ltout => \this_vga_signals.g2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g3_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000110011"
        )
    port map (
            in0 => \N__7613\,
            in1 => \N__11169\,
            in2 => \N__7619\,
            in3 => \N__17102\,
            lcout => OPEN,
            ltout => \this_vga_signals.g3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_0_i_a4_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000001"
        )
    port map (
            in0 => \N__8804\,
            in1 => \N__12336\,
            in2 => \N__7616\,
            in3 => \N__11462\,
            lcout => \this_vga_signals.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g2_4_0_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11331\,
            in2 => \_gnd_net_\,
            in3 => \N__11504\,
            lcout => \this_vga_signals.g2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_0_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__7769\,
            in1 => \N__7703\,
            in2 => \_gnd_net_\,
            in3 => \N__17320\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g1_8_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12459\,
            in1 => \N__12140\,
            in2 => \_gnd_net_\,
            in3 => \N__11028\,
            lcout => \this_vga_signals.g1_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc1_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101011010"
        )
    port map (
            in0 => \N__11503\,
            in1 => \N__12508\,
            in2 => \N__11408\,
            in3 => \N__12548\,
            lcout => \this_vga_signals.mult1_un54_sum_i_1\,
            ltout => \this_vga_signals.mult1_un54_sum_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x2_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12139\,
            in2 => \N__7697\,
            in3 => \N__17101\,
            lcout => \this_vga_signals.g0_i_x2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_1_N_3L3_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__11505\,
            in1 => \N__17118\,
            in2 => \_gnd_net_\,
            in3 => \N__10899\,
            lcout => \this_vga_signals.g0_1_N_3L3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_RNIJVJM_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8237\,
            lcout => OPEN,
            ltout => \this_vga_signals.un11_address_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_5_1_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001010000"
        )
    port map (
            in0 => \N__9013\,
            in1 => \N__7906\,
            in2 => \N__7694\,
            in3 => \N__7844\,
            lcout => \this_vga_signals.g0_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_x0_3_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001100111001"
        )
    port map (
            in0 => \N__7963\,
            in1 => \N__7750\,
            in2 => \N__7985\,
            in3 => \N__17299\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_i_x0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_i_ns_3_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__17300\,
            in1 => \N__7751\,
            in2 => \N__7691\,
            in3 => \N__7942\,
            lcout => this_vga_signals_un16_address_if_generate_plus_mult1_un54_sum_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_c_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__8102\,
            in1 => \N__7765\,
            in2 => \N__17319\,
            in3 => \N__8002\,
            lcout => \this_vga_signals.mult1_un54_sum_ac0_3_c\,
            ltout => \this_vga_signals.mult1_un54_sum_ac0_3_c_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001101"
        )
    port map (
            in0 => \N__17298\,
            in1 => \N__7984\,
            in2 => \N__7967\,
            in3 => \N__7962\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_1_N_5L8_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010001"
        )
    port map (
            in0 => \N__7943\,
            in1 => \N__7934\,
            in2 => \N__7922\,
            in3 => \N__17301\,
            lcout => \this_vga_signals.g0_1_N_5L8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb2_0_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100111000011"
        )
    port map (
            in0 => \N__7898\,
            in1 => \N__8090\,
            in2 => \N__9020\,
            in3 => \N__7834\,
            lcout => \this_vga_signals.mult1_un54_sum_axb2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un40_sum_axb1_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8119\,
            in2 => \_gnd_net_\,
            in3 => \N__8894\,
            lcout => \this_vga_signals.mult1_un40_sum_axb1\,
            ltout => \this_vga_signals.mult1_un40_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_0_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9011\,
            in1 => \N__7730\,
            in2 => \N__7754\,
            in3 => \N__18337\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_5_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__7739\,
            in1 => \N__11496\,
            in2 => \N__11457\,
            in3 => \N__12509\,
            lcout => \this_vga_signals.if_N_13_i_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9010\,
            in1 => \N__7729\,
            in2 => \N__17318\,
            in3 => \N__18338\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_1_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__7712\,
            in1 => \_gnd_net_\,
            in2 => \N__7706\,
            in3 => \N__9135\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_35_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11413\,
            in2 => \N__8147\,
            in3 => \N__12297\,
            lcout => \this_vga_signals.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIL7SG_4_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__8066\,
            in1 => \N__8325\,
            in2 => \N__8290\,
            in3 => \N__8460\,
            lcout => \this_vga_signals.un11_address_c4_i\,
            ltout => \this_vga_signals.un11_address_c4_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_1_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010101101001"
        )
    port map (
            in0 => \N__8091\,
            in1 => \N__9475\,
            in2 => \N__8132\,
            in3 => \N__8474\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_5_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_4_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8125\,
            in1 => \N__8891\,
            in2 => \N__8129\,
            in3 => \N__18303\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_5_4\,
            ltout => \this_vga_signals.mult1_un54_sum_axb1_5_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un54_sum_axb1_5_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111010010"
        )
    port map (
            in0 => \N__8892\,
            in1 => \N__8126\,
            in2 => \N__8108\,
            in3 => \N__8986\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8218\,
            lcout => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8701\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18208\,
            ce => \N__8678\,
            sr => \N__8644\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8700\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18208\,
            ce => \N__8678\,
            sr => \N__8644\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIOJB1_5_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8065\,
            in2 => \N__8048\,
            in3 => \N__8021\,
            lcout => \this_vga_signals.SUM_2_i_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_0_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8323\,
            in1 => \N__8367\,
            in2 => \N__8414\,
            in3 => \N__8446\,
            lcout => \this_vga_signals.SUM_2_i_a4_a0_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIJK9S_8_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__9465\,
            in1 => \N__8486\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_vga_signals.SUM_2_i_a4_1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIJ3MB6_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__8473\,
            in1 => \N__8165\,
            in2 => \N__8480\,
            in3 => \N__8153\,
            lcout => \this_vga_signals.SUM_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_7_rep1_esr_RNIHIQV_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__8447\,
            in1 => \_gnd_net_\,
            in2 => \N__8379\,
            in3 => \N__8324\,
            lcout => OPEN,
            ltout => \this_vga_signals.un11_address_c5_a0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPM1_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111101110000"
        )
    port map (
            in0 => \N__8281\,
            in1 => \N__8220\,
            in2 => \N__8477\,
            in3 => \N__9257\,
            lcout => \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI1LPMZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_9_rep1_esr_RNIELM41_1_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8448\,
            in1 => \N__8409\,
            in2 => \N__8378\,
            in3 => \N__8322\,
            lcout => \this_vga_signals.SUM_2_i_a4_0_a0_2_3\,
            ltout => \this_vga_signals.SUM_2_i_a4_0_a0_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUK2_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110000"
        )
    port map (
            in0 => \N__8282\,
            in1 => \N__8219\,
            in2 => \N__8174\,
            in3 => \N__8171\,
            lcout => \this_vga_signals.SUM_2_i_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIQJ31_9_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__9258\,
            in1 => \N__9709\,
            in2 => \N__9484\,
            in3 => \N__8159\,
            lcout => \this_vga_signals.SUM_2_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11686\,
            in1 => \N__9901\,
            in2 => \N__9575\,
            in3 => \N__9574\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__18216\,
            ce => 'H',
            sr => \N__8640\
        );

    \this_vga_signals.M_vcounter_q_1_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11688\,
            in1 => \N__12441\,
            in2 => \_gnd_net_\,
            in3 => \N__8597\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__18216\,
            ce => 'H',
            sr => \N__8640\
        );

    \this_vga_signals.M_vcounter_q_2_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11687\,
            in1 => \N__12108\,
            in2 => \_gnd_net_\,
            in3 => \N__8594\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__18216\,
            ce => 'H',
            sr => \N__8640\
        );

    \this_vga_signals.M_vcounter_q_3_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11689\,
            in1 => \N__12257\,
            in2 => \_gnd_net_\,
            in3 => \N__8591\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__18216\,
            ce => 'H',
            sr => \N__8640\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11289\,
            in2 => \_gnd_net_\,
            in3 => \N__8588\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9873\,
            in3 => \N__8561\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9410\,
            in3 => \N__8537\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9721\,
            in2 => \_gnd_net_\,
            in3 => \N__8516\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9497\,
            in2 => \_gnd_net_\,
            in3 => \N__8489\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9259\,
            in2 => \_gnd_net_\,
            in3 => \N__8756\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIAA7K1_9_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__8708\,
            in1 => \N__10702\,
            in2 => \N__10778\,
            in3 => \N__10741\,
            lcout => \N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIC1AR_4_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__10511\,
            in1 => \N__10639\,
            in2 => \_gnd_net_\,
            in3 => \N__10595\,
            lcout => \this_vga_signals.hsync_1_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8702\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18223\,
            ce => \N__8681\,
            sr => \N__8639\
        );

    \this_vga_signals.rgb_cnst_i_o2_0_4_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13750\,
            in2 => \N__10410\,
            in3 => \N__12959\,
            lcout => \this_vga_signals.N_381_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_cnst_i_a5_0_4_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__15881\,
            in1 => \N__10392\,
            in2 => \N__13769\,
            in3 => \N__12958\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIS1MK91_9_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__20324\,
            in1 => \N__8609\,
            in2 => \N__8603\,
            in3 => \N__15880\,
            lcout => \this_vga_signals.N_371_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIUDBJI_0_9_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__10376\,
            in1 => \N__12987\,
            in2 => \N__13770\,
            in3 => \N__20289\,
            lcout => OPEN,
            ltout => \this_vga_signals.rgb_cnst_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIO6OD01_9_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__12986\,
            in1 => \N__13751\,
            in2 => \N__8600\,
            in3 => \N__15902\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_esr_RNIO6OD01Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIR0T9KU3_9_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14077\,
            in2 => \N__8831\,
            in3 => \N__12908\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x2_5_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16083\,
            in1 => \N__16121\,
            in2 => \N__8816\,
            in3 => \N__8795\,
            lcout => \this_vga_signals.g0_i_x2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_o2_1_x2_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10914\,
            in3 => \N__10964\,
            lcout => \this_vga_signals.N_10_i\,
            ltout => \this_vga_signals.N_10_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x2_5_1_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110100110"
        )
    port map (
            in0 => \N__17116\,
            in1 => \N__12335\,
            in2 => \N__8798\,
            in3 => \N__11451\,
            lcout => \this_vga_signals.g0_i_x2_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g4_0_0_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__10906\,
            in1 => \N__12332\,
            in2 => \N__11465\,
            in3 => \N__10966\,
            lcout => OPEN,
            ltout => \this_vga_signals.g4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g4_1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111101"
        )
    port map (
            in0 => \N__17117\,
            in1 => \N__8789\,
            in2 => \N__8780\,
            in3 => \N__11144\,
            lcout => \this_vga_signals.g4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_0_N_5L7_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000100000"
        )
    port map (
            in0 => \N__8777\,
            in1 => \N__8768\,
            in2 => \N__12170\,
            in3 => \N__16082\,
            lcout => \this_vga_signals.g0_i_0_N_5L7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x2_0_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12331\,
            in1 => \N__11450\,
            in2 => \_gnd_net_\,
            in3 => \N__10902\,
            lcout => \this_vga_signals.g0_i_x2_1_1\,
            ltout => \this_vga_signals.g0_i_x2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x1_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__11143\,
            in1 => \N__10965\,
            in2 => \N__8759\,
            in3 => \N__17115\,
            lcout => \this_vga_signals.g0_i_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17158\,
            in3 => \N__11147\,
            lcout => this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1,
            ltout => \this_vga_signals_un16_address_if_generate_plus_mult1_un61_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_0_i_a4_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__12333\,
            in1 => \N__9149\,
            in2 => \N__8861\,
            in3 => \N__16057\,
            lcout => \this_vga_signals.N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x0_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000010100"
        )
    port map (
            in0 => \N__10967\,
            in1 => \N__11148\,
            in2 => \N__17159\,
            in3 => \N__8858\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_ns_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8852\,
            in2 => \N__8846\,
            in3 => \N__16056\,
            lcout => \this_vga_signals.mult1_un68_sum_ac0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g1_1_1_a3_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10968\,
            in1 => \N__11455\,
            in2 => \_gnd_net_\,
            in3 => \N__10900\,
            lcout => \this_vga_signals.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m3_4_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17103\,
            in2 => \N__11005\,
            in3 => \N__11027\,
            lcout => this_vga_signals_un16_address_if_i1_mux_0,
            ltout => \this_vga_signals_un16_address_if_i1_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x2_0_i_o3_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__17110\,
            in1 => \_gnd_net_\,
            in2 => \N__8843\,
            in3 => \N__11149\,
            lcout => \this_vga_signals.N_6_i\,
            ltout => \this_vga_signals.N_6_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g1_0_a3_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001001001101"
        )
    port map (
            in0 => \N__12334\,
            in1 => \N__12168\,
            in2 => \N__8840\,
            in3 => \N__8837\,
            lcout => \this_vga_signals.g1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_axb1_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__10883\,
            in1 => \_gnd_net_\,
            in2 => \N__10971\,
            in3 => \N__11437\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m5_0_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__12304\,
            in1 => \N__10880\,
            in2 => \N__11461\,
            in3 => \N__10949\,
            lcout => \this_vga_signals.if_N_1_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_0_i_x2_1_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__10882\,
            in1 => \_gnd_net_\,
            in2 => \N__10970\,
            in3 => \N__11436\,
            lcout => \this_vga_signals.N_11_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_25_1_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100110011111"
        )
    port map (
            in0 => \N__9012\,
            in1 => \N__9142\,
            in2 => \N__9110\,
            in3 => \N__18359\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_25_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_25_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101101001"
        )
    port map (
            in0 => \N__9101\,
            in1 => \N__8870\,
            in2 => \N__9095\,
            in3 => \N__9091\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_13_i_i_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_9_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001010001000"
        )
    port map (
            in0 => \N__9050\,
            in1 => \N__11190\,
            in2 => \N__9053\,
            in3 => \N__17132\,
            lcout => \this_vga_signals.g2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g2_0_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000100001"
        )
    port map (
            in0 => \N__10881\,
            in1 => \N__12305\,
            in2 => \N__10969\,
            in3 => \N__11435\,
            lcout => \this_vga_signals.g2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIVRQGTU3_9_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14090\,
            in1 => \N__13082\,
            in2 => \_gnd_net_\,
            in3 => \N__9044\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIE9LD1_7_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000010011"
        )
    port map (
            in0 => \N__9861\,
            in1 => \N__9405\,
            in2 => \N__11418\,
            in3 => \N__9742\,
            lcout => OPEN,
            ltout => \this_vga_signals.un11_address_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_3_0_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110100110"
        )
    port map (
            in0 => \N__11348\,
            in1 => \N__9014\,
            in2 => \N__8897\,
            in3 => \N__8893\,
            lcout => \this_vga_signals.g0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__12440\,
            in1 => \N__9897\,
            in2 => \N__12138\,
            in3 => \N__12247\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_28_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_8_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__9650\,
            in1 => \N__9404\,
            in2 => \N__9521\,
            in3 => \N__9496\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIVV6F6_9_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11660\,
            in1 => \N__9570\,
            in2 => \N__9518\,
            in3 => \N__9263\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNIVV6F6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clock.M_counter_q_1_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15257\,
            in1 => \N__13040\,
            in2 => \_gnd_net_\,
            in3 => \N__9550\,
            lcout => \this_pixel_clock.M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIROQM_7_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9495\,
            in2 => \_gnd_net_\,
            in3 => \N__9743\,
            lcout => OPEN,
            ltout => \this_vga_signals.rgb297_i_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICM2P1_6_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__11406\,
            in1 => \N__9862\,
            in2 => \N__9413\,
            in3 => \N__9403\,
            lcout => \this_vga_signals.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI38HR1_5_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__9863\,
            in1 => \N__9287\,
            in2 => \_gnd_net_\,
            in3 => \N__11407\,
            lcout => \this_vga_signals.CO0_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clock.M_counter_q_RNIJR071_1_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15256\,
            in1 => \N__13039\,
            in2 => \_gnd_net_\,
            in3 => \N__9549\,
            lcout => \M_counter_q_RNIJR071_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__10772\,
            in1 => \N__10705\,
            in2 => \_gnd_net_\,
            in3 => \N__10739\,
            lcout => \this_vga_signals.N_33_0\,
            ltout => \this_vga_signals.N_33_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICLUO4_9_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9262\,
            in1 => \N__9163\,
            in2 => \N__9152\,
            in3 => \N__9589\,
            lcout => \this_vga_signals.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIF4AR_7_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10637\,
            in1 => \N__10738\,
            in2 => \_gnd_net_\,
            in3 => \N__10593\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI704B1_9_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__10706\,
            in1 => \_gnd_net_\,
            in2 => \N__9578\,
            in3 => \N__10773\,
            lcout => \N_23_0\,
            ltout => \N_23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clock.M_counter_q_RNIQR4I2_1_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15306\,
            in1 => \N__13038\,
            in2 => \N__9554\,
            in3 => \N__9551\,
            lcout => \M_counter_q_RNIQR4I2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11747\,
            in2 => \N__11618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_24_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11702\,
            in1 => \N__10325\,
            in2 => \_gnd_net_\,
            in3 => \N__9536\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__18217\,
            ce => 'H',
            sr => \N__11582\
        );

    \this_vga_signals.M_hcounter_q_3_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11699\,
            in1 => \N__10548\,
            in2 => \_gnd_net_\,
            in3 => \N__9533\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__18217\,
            ce => 'H',
            sr => \N__11582\
        );

    \this_vga_signals.M_hcounter_q_4_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11703\,
            in1 => \N__10510\,
            in2 => \_gnd_net_\,
            in3 => \N__9530\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__18217\,
            ce => 'H',
            sr => \N__11582\
        );

    \this_vga_signals.M_hcounter_q_5_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11700\,
            in1 => \N__10638\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__18217\,
            ce => 'H',
            sr => \N__11582\
        );

    \this_vga_signals.M_hcounter_q_6_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11704\,
            in1 => \N__10594\,
            in2 => \_gnd_net_\,
            in3 => \N__9524\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__18217\,
            ce => 'H',
            sr => \N__11582\
        );

    \this_vga_signals.M_hcounter_q_7_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11701\,
            in1 => \N__10740\,
            in2 => \_gnd_net_\,
            in3 => \N__9638\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__18217\,
            ce => 'H',
            sr => \N__11582\
        );

    \this_vga_signals.M_hcounter_q_8_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11705\,
            in1 => \N__10774\,
            in2 => \_gnd_net_\,
            in3 => \N__9635\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__18217\,
            ce => 'H',
            sr => \N__11582\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10701\,
            in2 => \_gnd_net_\,
            in3 => \N__9632\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18222\,
            ce => \N__10466\,
            sr => \N__11577\
        );

    \this_vga_signals.un16_address_g0_10_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010010000010"
        )
    port map (
            in0 => \N__16060\,
            in1 => \N__16136\,
            in2 => \N__12365\,
            in3 => \N__12055\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_30_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__12178\,
            in1 => \N__9629\,
            in2 => \N__9620\,
            in3 => \N__9617\,
            lcout => \this_vga_signals.N_9_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m2_0_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16058\,
            in1 => \N__11183\,
            in2 => \N__12364\,
            in3 => \N__17181\,
            lcout => \this_vga_signals.if_N_3_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_x2_1_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9611\,
            in1 => \N__16059\,
            in2 => \N__16146\,
            in3 => \N__10802\,
            lcout => \this_vga_signals.g0_i_x2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_1_0_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100101000"
        )
    port map (
            in0 => \N__12056\,
            in1 => \N__12356\,
            in2 => \N__16147\,
            in3 => \N__16061\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__12180\,
            in1 => \N__9602\,
            in2 => \N__9596\,
            in3 => \N__11077\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_i_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000010100"
        )
    port map (
            in0 => \N__12179\,
            in1 => \N__10112\,
            in2 => \N__10106\,
            in3 => \N__12475\,
            lcout => \this_vga_signals.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_7_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__10103\,
            in1 => \N__9911\,
            in2 => \N__10097\,
            in3 => \N__9938\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI3CNE3O2_9_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20291\,
            in1 => \N__10085\,
            in2 => \N__10079\,
            in3 => \N__10808\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_0_N_4L5_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9959\,
            in2 => \_gnd_net_\,
            in3 => \N__11076\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_0_N_4L5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_0_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010000010"
        )
    port map (
            in0 => \N__9881\,
            in1 => \N__9953\,
            in2 => \N__9947\,
            in3 => \N__9944\,
            lcout => \this_vga_signals.if_i4_mux_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g1_7_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10838\,
            in1 => \N__9932\,
            in2 => \N__9926\,
            in3 => \N__17164\,
            lcout => \this_vga_signals.g1_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_0_N_2L1_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12460\,
            in2 => \_gnd_net_\,
            in3 => \N__9905\,
            lcout => \this_vga_signals.g0_i_0_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIU721_7_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11438\,
            in1 => \N__9867\,
            in2 => \_gnd_net_\,
            in3 => \N__9741\,
            lcout => \this_vga_signals.M_vcounter_d_1_sqmuxa_i_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI39EPS4_9_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__10124\,
            in1 => \N__10142\,
            in2 => \N__20290\,
            in3 => \N__10130\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_m1_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10330\,
            in2 => \_gnd_net_\,
            in3 => \N__20148\,
            lcout => \this_vga_signals.mult1_un82_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_m7_0_x4_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101001010110"
        )
    port map (
            in0 => \N__10277\,
            in1 => \N__10331\,
            in2 => \N__17779\,
            in3 => \N__10551\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_8_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_m7_0_m2_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110001110"
        )
    port map (
            in0 => \N__11610\,
            in1 => \N__11746\,
            in2 => \N__10151\,
            in3 => \N__10148\,
            lcout => \this_vga_signals.mult1_un89_sum_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_m7_0_m2_0_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100101101111"
        )
    port map (
            in0 => \N__17769\,
            in1 => \N__10549\,
            in2 => \N__10334\,
            in3 => \N__10283\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un82_sum_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_0_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10550\,
            in1 => \N__17770\,
            in2 => \N__10136\,
            in3 => \N__10276\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_0\,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un89_sum_axbxc3_2_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__17774\,
            in1 => \N__10333\,
            in2 => \N__10133\,
            in3 => \N__10552\,
            lcout => \this_vga_signals.mult1_un89_sum_axbxc3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_c2_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010111011"
        )
    port map (
            in0 => \N__10332\,
            in1 => \N__11745\,
            in2 => \_gnd_net_\,
            in3 => \N__20149\,
            lcout => \this_vga_signals.mult1_un82_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101111010100"
        )
    port map (
            in0 => \N__10553\,
            in1 => \N__17775\,
            in2 => \N__10326\,
            in3 => \N__10118\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un54_sum_c3_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101000101"
        )
    port map (
            in0 => \N__10664\,
            in1 => \N__10655\,
            in2 => \N__10640\,
            in3 => \N__10592\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc1_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10636\,
            in2 => \N__10349\,
            in3 => \N__10508\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc1\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axbxc3_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__11901\,
            in1 => \N__11871\,
            in2 => \N__10346\,
            in3 => \N__10475\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un68_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_c3_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001110001"
        )
    port map (
            in0 => \N__10309\,
            in1 => \N__10535\,
            in2 => \N__10343\,
            in3 => \N__10275\,
            lcout => \this_vga_signals.mult1_un75_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__11872\,
            in1 => \N__10340\,
            in2 => \N__11903\,
            in3 => \N__10474\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_m7_0_o4_1_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101110001"
        )
    port map (
            in0 => \N__10308\,
            in1 => \N__11736\,
            in2 => \N__10286\,
            in3 => \N__10274\,
            lcout => \this_vga_signals.if_N_9_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_axb1_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__10509\,
            in1 => \N__11897\,
            in2 => \_gnd_net_\,
            in3 => \N__11870\,
            lcout => \this_vga_signals.mult1_un68_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111010111"
        )
    port map (
            in0 => \N__10771\,
            in1 => \N__10737\,
            in2 => \N__10704\,
            in3 => \N__10591\,
            lcout => \this_vga_signals.SUM_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000101111111"
        )
    port map (
            in0 => \N__10588\,
            in1 => \N__10689\,
            in2 => \N__10742\,
            in3 => \N__10769\,
            lcout => \this_vga_signals.SUM_3\,
            ltout => \this_vga_signals.SUM_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_1_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011111111111"
        )
    port map (
            in0 => \N__10506\,
            in1 => \N__10631\,
            in2 => \N__10781\,
            in3 => \N__10589\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110101000010"
        )
    port map (
            in0 => \N__10770\,
            in1 => \N__10733\,
            in2 => \N__10703\,
            in3 => \N__10587\,
            lcout => \this_vga_signals.N_34\,
            ltout => \this_vga_signals.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_1_0_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100011111"
        )
    port map (
            in0 => \N__10630\,
            in1 => \N__10505\,
            in2 => \N__10658\,
            in3 => \N__10653\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un61_sum_axbxc3_2_2_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100000"
        )
    port map (
            in0 => \N__10654\,
            in1 => \N__10632\,
            in2 => \N__10598\,
            in3 => \N__10590\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_address_if_generate_plus_mult1_un68_sum_c2_0_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111011101"
        )
    port map (
            in0 => \N__10534\,
            in1 => \N__10507\,
            in2 => \N__10478\,
            in3 => \N__11896\,
            lcout => \this_vga_signals.mult1_un68_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11567\,
            in2 => \_gnd_net_\,
            in3 => \N__11693\,
            lcout => \this_vga_signals.N_469_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_RNI18AF_4_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__12824\,
            in1 => \N__12841\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => debug_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_cnst_i_a5_0_0_3_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__15816\,
            in1 => \N__18943\,
            in2 => \N__15879\,
            in3 => \N__18404\,
            lcout => \this_vga_signals.rgb_cnst_i_a5_0_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIETEJ4_2_11_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18944\,
            in1 => \N__18397\,
            in2 => \_gnd_net_\,
            in3 => \N__15800\,
            lcout => \M_this_vram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m3_5_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17180\,
            in1 => \N__10832\,
            in2 => \N__12398\,
            in3 => \N__11043\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m5_4_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010111"
        )
    port map (
            in0 => \N__12181\,
            in1 => \N__12473\,
            in2 => \N__10820\,
            in3 => \N__10817\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m5_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIC40KO51_3_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10793\,
            in1 => \N__11057\,
            in2 => \N__10811\,
            in3 => \N__12057\,
            lcout => \this_vga_signals.g1_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_o2_1_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__10980\,
            in1 => \N__12348\,
            in2 => \N__11458\,
            in3 => \N__10915\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_1_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__11422\,
            in1 => \N__10916\,
            in2 => \_gnd_net_\,
            in3 => \N__17178\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_axb2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axb2_0_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12347\,
            in1 => \N__11173\,
            in2 => \N__10796\,
            in3 => \N__10981\,
            lcout => \this_vga_signals.mult1_un68_sum_axb2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIRV8NA3_3_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11174\,
            in1 => \N__12349\,
            in2 => \_gnd_net_\,
            in3 => \N__17179\,
            lcout => \this_vga_signals.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_m2_5_0_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16086\,
            in1 => \N__10787\,
            in2 => \_gnd_net_\,
            in3 => \N__16140\,
            lcout => \this_vga_signals.if_m2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un68_sum_axbxc3_0_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12394\,
            in1 => \N__11044\,
            in2 => \_gnd_net_\,
            in3 => \N__17162\,
            lcout => \this_vga_signals.mult1_un68_sum_axbxc3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_1_1_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17163\,
            in1 => \N__12351\,
            in2 => \_gnd_net_\,
            in3 => \N__11192\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_21_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001000"
        )
    port map (
            in0 => \N__16085\,
            in1 => \N__12172\,
            in2 => \N__11096\,
            in3 => \N__12058\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_ac0_3_d_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_17_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__11093\,
            in1 => \N__12578\,
            in2 => \N__11084\,
            in3 => \N__11081\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_o2_0_0_x2_0_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11191\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17161\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_i_o2_0_0_x2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_o2_0_0_o4_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110111010100"
        )
    port map (
            in0 => \N__12171\,
            in1 => \N__12352\,
            in2 => \N__11060\,
            in3 => \N__16084\,
            lcout => \this_vga_signals.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_i_3_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001100110110"
        )
    port map (
            in0 => \N__17187\,
            in1 => \N__11193\,
            in2 => \N__11051\,
            in3 => \N__11006\,
            lcout => rgb_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_if_generate_plus_mult1_un61_sum_c2_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__11442\,
            in1 => \N__10987\,
            in2 => \N__12354\,
            in3 => \N__10912\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_o2_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__11443\,
            in1 => \N__10988\,
            in2 => \N__12355\,
            in3 => \N__10913\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_0_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__12593\,
            in1 => \N__15576\,
            in2 => \N__11912\,
            in3 => \N__16327\,
            lcout => \M_current_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18201\,
            ce => 'H',
            sr => \N__15321\
        );

    \M_current_address_q_RNO_0_0_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__16460\,
            in1 => \N__12627\,
            in2 => \N__17622\,
            in3 => \N__16326\,
            lcout => \N_401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIKNO0B_9_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__20266\,
            in1 => \N__11902\,
            in2 => \_gnd_net_\,
            in3 => \N__11873\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_1_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11707\,
            in2 => \N__11614\,
            in3 => \N__11735\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18214\,
            ce => 'H',
            sr => \N__11578\
        );

    \this_vga_signals.M_hcounter_q_0_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__11708\,
            in1 => \N__11606\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18214\,
            ce => 'H',
            sr => \N__11578\
        );

    \this_vga_signals.un16_address_g0_1_N_7L13_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12350\,
            in1 => \N__11194\,
            in2 => \_gnd_net_\,
            in3 => \N__17197\,
            lcout => \this_vga_signals.g0_1_N_7L13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_bm_1_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14889\,
            in1 => \N__14006\,
            in2 => \_gnd_net_\,
            in3 => \N__13066\,
            lcout => \this_vga_signals.rgb_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11531\,
            lcout => \this_delay_clk.M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18189\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_23_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__12563\,
            in1 => \N__11513\,
            in2 => \N__11459\,
            in3 => \N__12527\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_N_13_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_20_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011110101"
        )
    port map (
            in0 => \N__17198\,
            in1 => \_gnd_net_\,
            in2 => \N__11198\,
            in3 => \N__11195\,
            lcout => \this_vga_signals.if_N_16_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_1_N_6L11_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011001011001"
        )
    port map (
            in0 => \N__12572\,
            in1 => \N__12562\,
            in2 => \N__12523\,
            in3 => \N__12485\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_N_6L11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_1_N_8L15_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010001000010"
        )
    port map (
            in0 => \N__12173\,
            in1 => \N__12474\,
            in2 => \N__12401\,
            in3 => \N__12390\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_N_8L15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_1_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010101001"
        )
    port map (
            in0 => \N__12174\,
            in1 => \N__12374\,
            in2 => \N__12368\,
            in3 => \N__16087\,
            lcout => \this_vga_signals.if_N_6_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_vga_signals_address_a0_b_0_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__16142\,
            in1 => \N__16093\,
            in2 => \_gnd_net_\,
            in3 => \N__17879\,
            lcout => a0_b_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_i_o2_0_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101110001110"
        )
    port map (
            in0 => \N__12353\,
            in1 => \N__16141\,
            in2 => \N__12182\,
            in3 => \N__16088\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un68_sum_c2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un16_address_g0_0_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16089\,
            in1 => \N__12059\,
            in2 => \N__12032\,
            in3 => \N__12029\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI10UUE23_9_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000100"
        )
    port map (
            in0 => \N__20473\,
            in1 => \N__20298\,
            in2 => \N__12023\,
            in3 => \N__20449\,
            lcout => \M_this_vga_signals_address_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12857\,
            lcout => \this_start_data_delay_M_last_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIMM211_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101110"
        )
    port map (
            in0 => \N__15558\,
            in1 => \N__16301\,
            in2 => \N__12746\,
            in3 => \N__12800\,
            lcout => \N_312_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_RNIBJQQ_4_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__12744\,
            in1 => \N__12856\,
            in2 => \_gnd_net_\,
            in3 => \N__12822\,
            lcout => \N_349_0\,
            ltout => \N_349_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_8_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16302\,
            in1 => \N__16636\,
            in2 => \N__12860\,
            in3 => \N__13870\,
            lcout => \N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_RNI18AF_0_4_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12855\,
            in2 => \_gnd_net_\,
            in3 => \N__12821\,
            lcout => debug_0,
            ltout => \debug_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_address_ibuf_RNIR5I81_7_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__12794\,
            in1 => \N__12770\,
            in2 => \N__12749\,
            in3 => \N__12745\,
            lcout => \M_state_q_ns_0_a3_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_0_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12628\,
            in2 => \N__12608\,
            in3 => \N__12607\,
            lcout => \M_current_address_q_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \un1_M_current_address_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_1_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13135\,
            in2 => \_gnd_net_\,
            in3 => \N__12587\,
            lcout => \M_current_address_q_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_0\,
            carryout => \un1_M_current_address_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_2_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15619\,
            in2 => \_gnd_net_\,
            in3 => \N__12584\,
            lcout => \M_current_address_q_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_1\,
            carryout => \un1_M_current_address_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_3_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13407\,
            in2 => \_gnd_net_\,
            in3 => \N__12581\,
            lcout => \M_current_address_q_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_2\,
            carryout => \un1_M_current_address_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_4_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14575\,
            in2 => \_gnd_net_\,
            in3 => \N__12887\,
            lcout => \M_current_address_q_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_3\,
            carryout => \un1_M_current_address_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_5_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13270\,
            in2 => \_gnd_net_\,
            in3 => \N__12884\,
            lcout => \M_current_address_q_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_4\,
            carryout => \un1_M_current_address_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_6_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15358\,
            in2 => \_gnd_net_\,
            in3 => \N__12881\,
            lcout => \M_current_address_q_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_5\,
            carryout => \un1_M_current_address_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_7_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14716\,
            in2 => \_gnd_net_\,
            in3 => \N__12878\,
            lcout => \M_current_address_q_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_6\,
            carryout => \un1_M_current_address_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_8_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13866\,
            in2 => \_gnd_net_\,
            in3 => \N__12875\,
            lcout => \M_current_address_q_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \un1_M_current_address_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_9_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15127\,
            in2 => \_gnd_net_\,
            in3 => \N__12872\,
            lcout => \M_current_address_q_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_8\,
            carryout => \un1_M_current_address_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_10_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13543\,
            in2 => \_gnd_net_\,
            in3 => \N__12869\,
            lcout => \M_current_address_q_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_9\,
            carryout => \un1_M_current_address_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_11_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19390\,
            in2 => \_gnd_net_\,
            in3 => \N__12866\,
            lcout => \M_current_address_q_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_10\,
            carryout => \un1_M_current_address_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_12_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19544\,
            in2 => \_gnd_net_\,
            in3 => \N__12863\,
            lcout => \M_current_address_q_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_current_address_q_cry_11\,
            carryout => \un1_M_current_address_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_1_13_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19462\,
            in2 => \_gnd_net_\,
            in3 => \N__13043\,
            lcout => \M_current_address_q_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clock.M_counter_q_0_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15308\,
            in2 => \_gnd_net_\,
            in3 => \N__13032\,
            lcout => \this_pixel_clock.M_counter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_1_11_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18974\,
            in1 => \N__18485\,
            in2 => \_gnd_net_\,
            in3 => \N__15836\,
            lcout => \M_this_vram_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_bm_0_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12896\,
            in1 => \N__14479\,
            in2 => \_gnd_net_\,
            in3 => \N__14904\,
            lcout => \this_vga_signals.rgb_bmZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_bm_2_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14905\,
            in1 => \N__14480\,
            in2 => \_gnd_net_\,
            in3 => \N__13100\,
            lcout => \this_vga_signals.rgb_bmZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m7_am_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101110"
        )
    port map (
            in0 => \N__16768\,
            in1 => \N__16931\,
            in2 => \N__17006\,
            in3 => \N__16847\,
            lcout => OPEN,
            ltout => \m7_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m7_ns_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14948\,
            in2 => \N__12899\,
            in3 => \N__13112\,
            lcout => m7_ns,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m28_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100101000"
        )
    port map (
            in0 => \N__16846\,
            in1 => \N__17002\,
            in2 => \N__16934\,
            in3 => \N__16767\,
            lcout => OPEN,
            ltout => \m28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m29_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__14947\,
            in1 => \_gnd_net_\,
            in2 => \N__12890\,
            in3 => \N__14513\,
            lcout => m29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m32_am_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000101001000"
        )
    port map (
            in0 => \N__16999\,
            in1 => \N__16843\,
            in2 => \N__16932\,
            in3 => \N__16762\,
            lcout => OPEN,
            ltout => \m32_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m32_ns_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__14938\,
            in1 => \_gnd_net_\,
            in2 => \N__13115\,
            in3 => \N__13106\,
            lcout => m32_ns,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m7_bm_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011000000"
        )
    port map (
            in0 => \N__17001\,
            in1 => \N__16845\,
            in2 => \N__16933\,
            in3 => \N__16766\,
            lcout => m7_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m32_bm_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101010010"
        )
    port map (
            in0 => \N__16844\,
            in1 => \N__17000\,
            in2 => \N__16769\,
            in3 => \N__16924\,
            lcout => m32_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_11_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__19382\,
            in1 => \N__16436\,
            in2 => \N__16310\,
            in3 => \N__13828\,
            lcout => \N_412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m42_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14890\,
            in1 => \N__13099\,
            in2 => \_gnd_net_\,
            in3 => \N__14498\,
            lcout => rgb_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_5_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__16285\,
            in1 => \N__13269\,
            in2 => \N__13696\,
            in3 => \N__16450\,
            lcout => \N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_RNO_1_1_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16437\,
            in2 => \_gnd_net_\,
            in3 => \N__15529\,
            lcout => \N_352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.rgb_bm_3_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14447\,
            in1 => \N__14891\,
            in2 => \_gnd_net_\,
            in3 => \N__13070\,
            lcout => \this_vga_signals.rgb_bmZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_10_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__13542\,
            in1 => \N__16438\,
            in2 => \N__18050\,
            in3 => \N__16286\,
            lcout => \N_411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_3_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__16284\,
            in1 => \N__18049\,
            in2 => \N__13408\,
            in3 => \N__16449\,
            lcout => \N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_12_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__19545\,
            in1 => \N__16451\,
            in2 => \N__13697\,
            in3 => \N__16294\,
            lcout => OPEN,
            ltout => \N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_12_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__16295\,
            in1 => \N__15575\,
            in2 => \N__13664\,
            in3 => \N__13661\,
            lcout => \M_current_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18192\,
            ce => 'H',
            sr => \N__15323\
        );

    \M_current_address_q_10_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__15573\,
            in1 => \N__16296\,
            in2 => \N__13655\,
            in3 => \N__13646\,
            lcout => \M_current_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18192\,
            ce => 'H',
            sr => \N__15323\
        );

    \M_current_address_q_3_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__15574\,
            in1 => \N__16297\,
            in2 => \N__13523\,
            in3 => \N__13514\,
            lcout => \M_current_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18192\,
            ce => 'H',
            sr => \N__15323\
        );

    \M_current_address_q_5_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__13382\,
            in1 => \N__15555\,
            in2 => \N__13376\,
            in3 => \N__16298\,
            lcout => \M_current_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18192\,
            ce => 'H',
            sr => \N__15323\
        );

    \M_current_address_q_RNO_0_1_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__16462\,
            in1 => \N__13134\,
            in2 => \N__16635\,
            in3 => \N__16312\,
            lcout => OPEN,
            ltout => \N_402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_1_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__15569\,
            in1 => \N__16328\,
            in2 => \N__13250\,
            in3 => \N__13247\,
            lcout => \M_current_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18195\,
            ce => 'H',
            sr => \N__15307\
        );

    \M_current_address_q_8_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111010000100"
        )
    port map (
            in0 => \N__16314\,
            in1 => \N__13991\,
            in2 => \N__15578\,
            in3 => \N__13985\,
            lcout => \M_current_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18195\,
            ce => 'H',
            sr => \N__15307\
        );

    \M_current_address_q_11_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110101001000"
        )
    port map (
            in0 => \N__16313\,
            in1 => \N__13844\,
            in2 => \N__15577\,
            in3 => \N__13835\,
            lcout => \M_current_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18195\,
            ce => 'H',
            sr => \N__15307\
        );

    \M_current_address_q_RNO_0_4_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__16311\,
            in1 => \N__14568\,
            in2 => \N__13829\,
            in3 => \N__16461\,
            lcout => \N_405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_9_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__16321\,
            in1 => \N__15565\,
            in2 => \N__15107\,
            in3 => \N__13799\,
            lcout => \M_current_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18200\,
            ce => 'H',
            sr => \N__15312\
        );

    \this_vram.mem_radreg_RNIETEJ4_1_11_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__15841\,
            in1 => \N__18737\,
            in2 => \N__18518\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vram_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb291_cry_0_c_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14018\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => rgb291_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb291_cry_1_c_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14150\,
            in2 => \N__14978\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => rgb291_cry_0,
            carryout => rgb291_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb291_cry_2_c_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15773\,
            in2 => \N__14182\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => rgb291_cry_1,
            carryout => rgb291_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb291_cry_3_c_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14024\,
            in2 => \N__14183\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => rgb291_cry_2,
            carryout => rgb291,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI4ODS4_9_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20329\,
            in2 => \_gnd_net_\,
            in3 => \N__14096\,
            lcout => \this_vga_signals.rgb_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_0_11_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15838\,
            in1 => \N__18973\,
            in2 => \_gnd_net_\,
            in3 => \N__18484\,
            lcout => \mem_radreg_RNIMTEJ4_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIETEJ4_0_11_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18396\,
            in1 => \N__18936\,
            in2 => \_gnd_net_\,
            in3 => \N__15837\,
            lcout => \mem_radreg_RNIETEJ4_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m44_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011010000"
        )
    port map (
            in0 => \N__16908\,
            in1 => \N__16986\,
            in2 => \N__16842\,
            in3 => \N__16747\,
            lcout => OPEN,
            ltout => \m44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m46_bm_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__14512\,
            in1 => \_gnd_net_\,
            in2 => \N__14012\,
            in3 => \N__14951\,
            lcout => m46_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m22_am_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010110000"
        )
    port map (
            in0 => \N__16984\,
            in1 => \N__16906\,
            in2 => \N__16760\,
            in3 => \N__16825\,
            lcout => OPEN,
            ltout => \m22_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m22_ns_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__13997\,
            in1 => \_gnd_net_\,
            in2 => \N__14009\,
            in3 => \N__14937\,
            lcout => m22_ns,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m22_bm_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101100"
        )
    port map (
            in0 => \N__16985\,
            in1 => \N__16907\,
            in2 => \N__16761\,
            in3 => \N__16826\,
            lcout => m22_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m24_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100001001000"
        )
    port map (
            in0 => \N__16809\,
            in1 => \N__16970\,
            in2 => \N__16740\,
            in3 => \N__16887\,
            lcout => m24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m40_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101001"
        )
    port map (
            in0 => \N__16971\,
            in1 => \N__16810\,
            in2 => \N__16905\,
            in3 => \N__16727\,
            lcout => OPEN,
            ltout => \m40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m41_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__14492\,
            in1 => \_gnd_net_\,
            in2 => \N__14501\,
            in3 => \N__14936\,
            lcout => m41,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m10_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111100"
        )
    port map (
            in0 => \N__16968\,
            in1 => \N__16807\,
            in2 => \N__16903\,
            in3 => \N__16722\,
            lcout => m10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI1UGICK_9_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__14465\,
            in1 => \N__17873\,
            in2 => \_gnd_net_\,
            in3 => \N__17169\,
            lcout => rgb_1_axb_0,
            ltout => \rgb_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m15_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14491\,
            in2 => \N__14483\,
            in3 => \N__15767\,
            lcout => m15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m19_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110001000"
        )
    port map (
            in0 => \N__16969\,
            in1 => \N__16808\,
            in2 => \N__16904\,
            in3 => \N__16723\,
            lcout => m19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_1_cry_0_0_c_RNO_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101011000000"
        )
    port map (
            in0 => \N__17869\,
            in1 => \N__14461\,
            in2 => \N__17878\,
            in3 => \N__17199\,
            lcout => \rgb_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m37_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14949\,
            in1 => \N__14962\,
            in2 => \_gnd_net_\,
            in3 => \N__16687\,
            lcout => m37,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m46_am_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16688\,
            in1 => \N__14963\,
            in2 => \_gnd_net_\,
            in3 => \N__14950\,
            lcout => OPEN,
            ltout => \m46_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m46_ns_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14906\,
            in2 => \N__14861\,
            in3 => \N__14858\,
            lcout => rgb_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_1_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__15325\,
            in1 => \N__14834\,
            in2 => \N__14549\,
            in3 => \N__16643\,
            lcout => \M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_0_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110010"
        )
    port map (
            in0 => \N__16241\,
            in1 => \N__15326\,
            in2 => \N__14522\,
            in3 => \N__16453\,
            lcout => \M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_RNIMM211_1_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16452\,
            in1 => \N__15522\,
            in2 => \_gnd_net_\,
            in3 => \N__16240\,
            lcout => \M_this_vram_write_en_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_7_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__14712\,
            in1 => \N__16473\,
            in2 => \N__16325\,
            in3 => \N__17623\,
            lcout => OPEN,
            ltout => \N_408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_7_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__16299\,
            in1 => \N__15557\,
            in2 => \N__14828\,
            in3 => \N__14825\,
            lcout => \M_current_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18197\,
            ce => 'H',
            sr => \N__15324\
        );

    \M_current_address_q_4_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__15556\,
            in1 => \N__16300\,
            in2 => \N__14693\,
            in3 => \N__14684\,
            lcout => \M_current_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18197\,
            ce => 'H',
            sr => \N__15324\
        );

    \M_state_q_RNO_0_0_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__16678\,
            in1 => \N__14545\,
            in2 => \N__19964\,
            in3 => \N__15530\,
            lcout => \N_351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_2_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__15606\,
            in1 => \N__16317\,
            in2 => \N__16478\,
            in3 => \N__19771\,
            lcout => OPEN,
            ltout => \N_403_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_2_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__16318\,
            in1 => \N__15564\,
            in2 => \N__15725\,
            in3 => \N__15722\,
            lcout => \M_current_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18202\,
            ce => 'H',
            sr => \N__15322\
        );

    \M_current_address_q_13_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__15562\,
            in1 => \N__16319\,
            in2 => \N__16160\,
            in3 => \N__15587\,
            lcout => \M_current_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18202\,
            ce => 'H',
            sr => \N__15322\
        );

    \M_current_address_q_RNO_0_6_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__16316\,
            in1 => \N__15345\,
            in2 => \N__16376\,
            in3 => \N__16477\,
            lcout => OPEN,
            ltout => \N_407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_6_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__15563\,
            in1 => \N__16320\,
            in2 => \N__15473\,
            in3 => \N__15470\,
            lcout => \M_current_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18202\,
            ce => 'H',
            sr => \N__15322\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICJRF0D_9_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17201\,
            lcout => \M_vcounter_q_esr_RNICJRF0D_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_9_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__15126\,
            in1 => \N__16472\,
            in2 => \N__19772\,
            in3 => \N__16315\,
            lcout => \N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIRM6F7_9_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__20262\,
            in1 => \N__15098\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIETEJ4_11_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18514\,
            in1 => \N__18736\,
            in2 => \_gnd_net_\,
            in3 => \N__15842\,
            lcout => \mem_radreg_RNIETEJ4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_2_11_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15840\,
            in1 => \N__19067\,
            in2 => \_gnd_net_\,
            in3 => \N__18821\,
            lcout => \M_this_vram_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNIMTEJ4_11_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18820\,
            in1 => \N__19066\,
            in2 => \_gnd_net_\,
            in3 => \N__15839\,
            lcout => \mem_radreg_RNIMTEJ4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIB9J4TN_9_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001001000"
        )
    port map (
            in0 => \N__17846\,
            in1 => \N__17170\,
            in2 => \N__17865\,
            in3 => \N__17351\,
            lcout => \M_vcounter_q_esr_RNIB9J4TN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m14_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100110100"
        )
    port map (
            in0 => \N__16880\,
            in1 => \N__16967\,
            in2 => \N__16824\,
            in3 => \N__16721\,
            lcout => m14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_1_cry_0_0_c_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15761\,
            in2 => \N__17021\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => rgb_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_1_cry_0_0_c_RNIFFTTT41_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15755\,
            in2 => \N__15749\,
            in3 => \N__15737\,
            lcout => rgb_1_3,
            ltout => OPEN,
            carryin => rgb_1_cry_0,
            carryout => rgb_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_1_cry_1_0_c_RNIPTLTE01_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17012\,
            in2 => \N__17795\,
            in3 => \N__15734\,
            lcout => rgb_1_4,
            ltout => OPEN,
            carryin => rgb_1_cry_1,
            carryout => rgb_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_1_cry_2_0_c_RNISLC8LA_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17885\,
            in2 => \_gnd_net_\,
            in3 => \N__15731\,
            lcout => rgb_1_5,
            ltout => OPEN,
            carryin => rgb_1_cry_2,
            carryout => rgb_1_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_1_6_THRU_LUT4_0_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15728\,
            lcout => \rgb_1_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_1_cry_0_0_c_RNO_0_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17832\,
            in2 => \_gnd_net_\,
            in3 => \N__17200\,
            lcout => \rgb_1_cry_0_0_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI1H9RHL_9_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101011000000"
        )
    port map (
            in0 => \N__17833\,
            in1 => \N__18363\,
            in2 => \N__17853\,
            in3 => \N__17350\,
            lcout => \M_vcounter_q_esr_RNI1H9RHL_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_2_5_0__m36_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110101111110"
        )
    port map (
            in0 => \N__16966\,
            in1 => \N__16879\,
            in2 => \N__16823\,
            in3 => \N__16720\,
            lcout => m36,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_state_q_RNO_0_1_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__16679\,
            in1 => \N__16655\,
            in2 => \N__19963\,
            in3 => \N__16287\,
            lcout => \M_state_q_ns_0_a3_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNI2PEE1_1_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16637\,
            in2 => \_gnd_net_\,
            in3 => \N__19251\,
            lcout => \M_this_vram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_current_address_q_RNO_0_13_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__19432\,
            in1 => \N__16471\,
            in2 => \N__16375\,
            in3 => \N__16309\,
            lcout => \N_414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIRN34U9_9_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20325\,
            in1 => \N__16148\,
            in2 => \_gnd_net_\,
            in3 => \N__16094\,
            lcout => \M_this_vga_signals_address_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIRB7JA_9_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17647\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15919\,
            lcout => \rgbZ0Z_1\,
            ltout => \rgbZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI2RH6LA_9_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__18370\,
            in1 => \_gnd_net_\,
            in2 => \N__17888\,
            in3 => \_gnd_net_\,
            lcout => \M_vcounter_q_esr_RNI2RH6LA_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIVLNKSA_9_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17339\,
            lcout => \M_vcounter_q_esr_RNIVLNKSA_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIN383L_9_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20308\,
            in2 => \_gnd_net_\,
            in3 => \N__17783\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNI1OEE1_0_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17627\,
            in2 => \_gnd_net_\,
            in3 => \N__19297\,
            lcout => \M_this_vram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIFAVQ5_9_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20310\,
            in2 => \_gnd_net_\,
            in3 => \N__17498\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_wclke_3_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__19595\,
            in1 => \N__19391\,
            in2 => \N__19499\,
            in3 => \N__19309\,
            lcout => \this_vram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_12_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20338\,
            in2 => \_gnd_net_\,
            in3 => \N__17349\,
            lcout => \this_vram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_wclke_3_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19579\,
            in1 => \N__19394\,
            in2 => \N__19500\,
            in3 => \N__19310\,
            lcout => \this_vram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNISOI11_0_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17219\,
            in1 => \N__19871\,
            in2 => \_gnd_net_\,
            in3 => \N__18533\,
            lcout => \this_vram.mem_mem_0_1_RNISOI11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5OL72_0_12_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18877\,
            in1 => \N__18680\,
            in2 => \_gnd_net_\,
            in3 => \N__18653\,
            lcout => \this_vram.mem_N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5GH72_12_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18593\,
            in1 => \N__18494\,
            in2 => \_gnd_net_\,
            in3 => \N__18866\,
            lcout => \this_vram.mem_N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_wclke_3_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__19312\,
            in1 => \N__19496\,
            in2 => \N__19601\,
            in3 => \N__19393\,
            lcout => \this_vram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_wclke_3_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19596\,
            in1 => \N__19392\,
            in2 => \N__19502\,
            in3 => \N__19311\,
            lcout => \this_vram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI1GH72_12_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18851\,
            in1 => \N__19799\,
            in2 => \_gnd_net_\,
            in3 => \N__19937\,
            lcout => \this_vram_mem_N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_13_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20339\,
            in2 => \_gnd_net_\,
            in3 => \N__18371\,
            lcout => \this_vram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNI4REE1_3_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18045\,
            in2 => \_gnd_net_\,
            in3 => \N__19276\,
            lcout => \M_this_vram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_0_LC_24_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17915\,
            in1 => \N__17903\,
            in2 => \_gnd_net_\,
            in3 => \N__19878\,
            lcout => \this_vram.mem_mem_0_0_RNIQOI11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_0_LC_24_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19879\,
            in1 => \N__18776\,
            in2 => \_gnd_net_\,
            in3 => \N__18764\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_0_RNIU0N11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI1GH72_0_12_LC_24_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__18746\,
            in1 => \_gnd_net_\,
            in2 => \N__18740\,
            in3 => \N__18878\,
            lcout => \this_vram.mem_N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_RNISSK11_0_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18707\,
            in1 => \N__19872\,
            in2 => \_gnd_net_\,
            in3 => \N__18695\,
            lcout => \this_vram.mem_mem_1_0_RNISSK11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_0_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18674\,
            in1 => \N__19877\,
            in2 => \_gnd_net_\,
            in3 => \N__18668\,
            lcout => \this_vram.mem_mem_3_0_RNI05P11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_0_RNISSK11_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__18647\,
            in1 => \_gnd_net_\,
            in2 => \N__19880\,
            in3 => \N__18635\,
            lcout => \this_vram.mem_mem_1_0_RNISSKZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNI01N11_0_LC_24_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18620\,
            in1 => \N__19876\,
            in2 => \_gnd_net_\,
            in3 => \N__18611\,
            lcout => \this_vram.mem_mem_2_1_RNI01N11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_1_RNISOI11_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18587\,
            in1 => \N__19868\,
            in2 => \_gnd_net_\,
            in3 => \N__18572\,
            lcout => \this_vram.mem_mem_0_1_RNISOIZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNIUSK11_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19869\,
            in1 => \N__18560\,
            in2 => \_gnd_net_\,
            in3 => \N__18548\,
            lcout => \this_vram.mem_mem_1_1_RNIUSKZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_1_RNI01N11_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19103\,
            in1 => \N__19094\,
            in2 => \_gnd_net_\,
            in3 => \N__19870\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_2_1_RNI01NZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5GH72_0_12_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18876\,
            in1 => \_gnd_net_\,
            in2 => \N__19076\,
            in3 => \N__19073\,
            lcout => \this_vram.mem_N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_1_1_RNIUSK11_0_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19046\,
            in1 => \N__19031\,
            in2 => \_gnd_net_\,
            in3 => \N__19841\,
            lcout => \this_vram.mem_mem_1_1_RNIUSK11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI25P11_0_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19842\,
            in1 => \_gnd_net_\,
            in2 => \N__19016\,
            in3 => \N__19007\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_3_1_RNI25P11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OL72_12_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18865\,
            in1 => \_gnd_net_\,
            in2 => \N__18986\,
            in3 => \N__18983\,
            lcout => \this_vram.mem_N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI5OL72_12_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18953\,
            in1 => \N__19907\,
            in2 => \_gnd_net_\,
            in3 => \N__18863\,
            lcout => \this_vram_mem_N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_1_RNI25P11_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18911\,
            in1 => \N__18905\,
            in2 => \_gnd_net_\,
            in3 => \N__19843\,
            lcout => OPEN,
            ltout => \this_vram.mem_mem_3_1_RNI25PZ0Z11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_radreg_RNI9OL72_0_12_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__18887\,
            in1 => \_gnd_net_\,
            in2 => \N__18881\,
            in3 => \N__18864\,
            lcout => \this_vram.mem_N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_2_0_RNIU0N11_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19822\,
            in1 => \N__18803\,
            in2 => \_gnd_net_\,
            in3 => \N__18788\,
            lcout => \this_vram.mem_mem_2_0_RNIU0NZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_3_0_RNI05P11_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19931\,
            in1 => \N__19823\,
            in2 => \_gnd_net_\,
            in3 => \N__19916\,
            lcout => \this_vram.mem_mem_3_0_RNI05PZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_0_0_RNIQOI11_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19901\,
            in1 => \N__19886\,
            in2 => \_gnd_net_\,
            in3 => \N__19821\,
            lcout => \this_vram.mem_mem_0_0_RNIQOIZ0Z11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_4_0_wclke_3_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19597\,
            in1 => \N__19402\,
            in2 => \N__19501\,
            in3 => \N__19316\,
            lcout => \this_vram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_data_ibuf_RNI3QEE1_2_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19767\,
            in2 => \_gnd_net_\,
            in3 => \N__19277\,
            lcout => \M_this_vram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_5_0_wclke_3_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19580\,
            in1 => \N__19403\,
            in2 => \N__19498\,
            in3 => \N__19313\,
            lcout => \this_vram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_7_0_wclke_3_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19315\,
            in1 => \N__19581\,
            in2 => \N__19497\,
            in3 => \N__19386\,
            lcout => \this_vram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vram.mem_mem_6_0_wclke_3_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19582\,
            in1 => \N__19480\,
            in2 => \N__19401\,
            in3 => \N__19314\,
            lcout => \this_vram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI51C6S_9_LC_24_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20332\,
            in2 => \_gnd_net_\,
            in3 => \N__20167\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNID2F8IP1_9_LC_24_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20333\,
            in1 => \N__20480\,
            in2 => \_gnd_net_\,
            in3 => \N__20459\,
            lcout => \M_this_vga_signals_address_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIGD3HC3_9_LC_24_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20334\,
            in1 => \N__20168\,
            in2 => \_gnd_net_\,
            in3 => \N__20135\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_address_ibuf_RNIPG5P_5_LC_32_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__20024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20018\,
            lcout => \M_state_q_ns_0_a3_0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \port_address_ibuf_RNI7ITU1_2_LC_32_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20006\,
            in1 => \N__19994\,
            in2 => \N__19982\,
            in3 => \N__19973\,
            lcout => \M_state_q_ns_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
