// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     Jun 20 2021 15:53:16

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    write_address,
    write_data,
    rgb,
    write_en,
    vsync,
    vblank,
    rst_n,
    hsync,
    hblank,
    clk);

    input [14:0] write_address;
    input [5:0] write_data;
    output [5:0] rgb;
    input write_en;
    output vsync;
    output vblank;
    input rst_n;
    output hsync;
    output hblank;
    input clk;

    wire N__15245;
    wire N__15244;
    wire N__15243;
    wire N__15234;
    wire N__15233;
    wire N__15232;
    wire N__15225;
    wire N__15224;
    wire N__15223;
    wire N__15216;
    wire N__15215;
    wire N__15214;
    wire N__15207;
    wire N__15206;
    wire N__15205;
    wire N__15198;
    wire N__15197;
    wire N__15196;
    wire N__15189;
    wire N__15188;
    wire N__15187;
    wire N__15180;
    wire N__15179;
    wire N__15178;
    wire N__15171;
    wire N__15170;
    wire N__15169;
    wire N__15162;
    wire N__15161;
    wire N__15160;
    wire N__15153;
    wire N__15152;
    wire N__15151;
    wire N__15144;
    wire N__15143;
    wire N__15142;
    wire N__15135;
    wire N__15134;
    wire N__15133;
    wire N__15126;
    wire N__15125;
    wire N__15124;
    wire N__15117;
    wire N__15116;
    wire N__15115;
    wire N__15108;
    wire N__15107;
    wire N__15106;
    wire N__15099;
    wire N__15098;
    wire N__15097;
    wire N__15090;
    wire N__15089;
    wire N__15088;
    wire N__15081;
    wire N__15080;
    wire N__15079;
    wire N__15072;
    wire N__15071;
    wire N__15070;
    wire N__15063;
    wire N__15062;
    wire N__15061;
    wire N__15054;
    wire N__15053;
    wire N__15052;
    wire N__15045;
    wire N__15044;
    wire N__15043;
    wire N__15036;
    wire N__15035;
    wire N__15034;
    wire N__15027;
    wire N__15026;
    wire N__15025;
    wire N__15018;
    wire N__15017;
    wire N__15016;
    wire N__15009;
    wire N__15008;
    wire N__15007;
    wire N__15000;
    wire N__14999;
    wire N__14998;
    wire N__14991;
    wire N__14990;
    wire N__14989;
    wire N__14982;
    wire N__14981;
    wire N__14980;
    wire N__14973;
    wire N__14972;
    wire N__14971;
    wire N__14964;
    wire N__14963;
    wire N__14962;
    wire N__14955;
    wire N__14954;
    wire N__14953;
    wire N__14946;
    wire N__14945;
    wire N__14944;
    wire N__14927;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14919;
    wire N__14914;
    wire N__14911;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14899;
    wire N__14896;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14885;
    wire N__14882;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14870;
    wire N__14865;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14847;
    wire N__14846;
    wire N__14845;
    wire N__14844;
    wire N__14839;
    wire N__14836;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14817;
    wire N__14814;
    wire N__14809;
    wire N__14804;
    wire N__14803;
    wire N__14802;
    wire N__14801;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14793;
    wire N__14790;
    wire N__14785;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14775;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14767;
    wire N__14764;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14738;
    wire N__14735;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14698;
    wire N__14697;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14680;
    wire N__14677;
    wire N__14676;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14659;
    wire N__14656;
    wire N__14651;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14639;
    wire N__14636;
    wire N__14631;
    wire N__14630;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14615;
    wire N__14614;
    wire N__14613;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14586;
    wire N__14583;
    wire N__14578;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14566;
    wire N__14565;
    wire N__14562;
    wire N__14557;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14521;
    wire N__14518;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14479;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14471;
    wire N__14468;
    wire N__14467;
    wire N__14466;
    wire N__14465;
    wire N__14464;
    wire N__14463;
    wire N__14462;
    wire N__14457;
    wire N__14456;
    wire N__14455;
    wire N__14454;
    wire N__14453;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14436;
    wire N__14435;
    wire N__14432;
    wire N__14431;
    wire N__14426;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14408;
    wire N__14407;
    wire N__14406;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14372;
    wire N__14365;
    wire N__14362;
    wire N__14361;
    wire N__14358;
    wire N__14357;
    wire N__14354;
    wire N__14349;
    wire N__14344;
    wire N__14339;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14311;
    wire N__14306;
    wire N__14299;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14247;
    wire N__14242;
    wire N__14239;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14177;
    wire N__14176;
    wire N__14175;
    wire N__14174;
    wire N__14173;
    wire N__14172;
    wire N__14171;
    wire N__14170;
    wire N__14169;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14161;
    wire N__14158;
    wire N__14157;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14145;
    wire N__14142;
    wire N__14141;
    wire N__14140;
    wire N__14139;
    wire N__14134;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14097;
    wire N__14096;
    wire N__14095;
    wire N__14092;
    wire N__14087;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14071;
    wire N__14066;
    wire N__14063;
    wire N__14058;
    wire N__14055;
    wire N__14050;
    wire N__14047;
    wire N__14042;
    wire N__14035;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13993;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13864;
    wire N__13861;
    wire N__13860;
    wire N__13859;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13821;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13805;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13781;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13760;
    wire N__13759;
    wire N__13758;
    wire N__13757;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13726;
    wire N__13725;
    wire N__13724;
    wire N__13723;
    wire N__13722;
    wire N__13721;
    wire N__13720;
    wire N__13719;
    wire N__13718;
    wire N__13717;
    wire N__13716;
    wire N__13715;
    wire N__13714;
    wire N__13713;
    wire N__13712;
    wire N__13711;
    wire N__13710;
    wire N__13709;
    wire N__13708;
    wire N__13707;
    wire N__13706;
    wire N__13705;
    wire N__13704;
    wire N__13703;
    wire N__13702;
    wire N__13701;
    wire N__13700;
    wire N__13699;
    wire N__13698;
    wire N__13697;
    wire N__13696;
    wire N__13695;
    wire N__13694;
    wire N__13693;
    wire N__13692;
    wire N__13691;
    wire N__13690;
    wire N__13689;
    wire N__13688;
    wire N__13687;
    wire N__13686;
    wire N__13685;
    wire N__13684;
    wire N__13683;
    wire N__13682;
    wire N__13681;
    wire N__13680;
    wire N__13679;
    wire N__13678;
    wire N__13677;
    wire N__13676;
    wire N__13675;
    wire N__13674;
    wire N__13673;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13669;
    wire N__13668;
    wire N__13667;
    wire N__13666;
    wire N__13665;
    wire N__13664;
    wire N__13663;
    wire N__13662;
    wire N__13661;
    wire N__13660;
    wire N__13659;
    wire N__13658;
    wire N__13657;
    wire N__13656;
    wire N__13655;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13447;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13403;
    wire N__13402;
    wire N__13401;
    wire N__13400;
    wire N__13397;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13383;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13378;
    wire N__13375;
    wire N__13372;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13354;
    wire N__13353;
    wire N__13352;
    wire N__13349;
    wire N__13348;
    wire N__13347;
    wire N__13344;
    wire N__13341;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13301;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13291;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13279;
    wire N__13278;
    wire N__13277;
    wire N__13276;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13266;
    wire N__13265;
    wire N__13262;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13239;
    wire N__13238;
    wire N__13237;
    wire N__13230;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13210;
    wire N__13209;
    wire N__13208;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13194;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13173;
    wire N__13172;
    wire N__13171;
    wire N__13162;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13150;
    wire N__13149;
    wire N__13148;
    wire N__13147;
    wire N__13146;
    wire N__13143;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13131;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13114;
    wire N__13111;
    wire N__13110;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13086;
    wire N__13085;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13071;
    wire N__13068;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13049;
    wire N__13042;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13030;
    wire N__13029;
    wire N__13026;
    wire N__13025;
    wire N__13022;
    wire N__13021;
    wire N__13018;
    wire N__13017;
    wire N__13016;
    wire N__13007;
    wire N__12998;
    wire N__12997;
    wire N__12994;
    wire N__12993;
    wire N__12990;
    wire N__12983;
    wire N__12980;
    wire N__12979;
    wire N__12964;
    wire N__12961;
    wire N__12956;
    wire N__12955;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12938;
    wire N__12935;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12912;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12897;
    wire N__12894;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12868;
    wire N__12865;
    wire N__12858;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12540;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12520;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12498;
    wire N__12491;
    wire N__12490;
    wire N__12489;
    wire N__12486;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12474;
    wire N__12471;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12382;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12355;
    wire N__12352;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12289;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12271;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12239;
    wire N__12236;
    wire N__12235;
    wire N__12230;
    wire N__12227;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12191;
    wire N__12188;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12176;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12164;
    wire N__12163;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12143;
    wire N__12140;
    wire N__12139;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12126;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12111;
    wire N__12110;
    wire N__12109;
    wire N__12108;
    wire N__12107;
    wire N__12102;
    wire N__12099;
    wire N__12090;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12076;
    wire N__12071;
    wire N__12070;
    wire N__12067;
    wire N__12066;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12016;
    wire N__12015;
    wire N__12012;
    wire N__12011;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11990;
    wire N__11987;
    wire N__11986;
    wire N__11985;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11936;
    wire N__11935;
    wire N__11934;
    wire N__11933;
    wire N__11930;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11908;
    wire N__11907;
    wire N__11906;
    wire N__11905;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11846;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11810;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11798;
    wire N__11797;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11784;
    wire N__11779;
    wire N__11776;
    wire N__11771;
    wire N__11770;
    wire N__11769;
    wire N__11768;
    wire N__11767;
    wire N__11764;
    wire N__11757;
    wire N__11754;
    wire N__11747;
    wire N__11746;
    wire N__11745;
    wire N__11744;
    wire N__11741;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11723;
    wire N__11714;
    wire N__11713;
    wire N__11712;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11690;
    wire N__11687;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11486;
    wire N__11485;
    wire N__11482;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11259;
    wire N__11256;
    wire N__11255;
    wire N__11252;
    wire N__11251;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11221;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11022;
    wire N__11019;
    wire N__11018;
    wire N__11015;
    wire N__11014;
    wire N__11011;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10984;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10963;
    wire N__10962;
    wire N__10961;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10949;
    wire N__10946;
    wire N__10937;
    wire N__10934;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10923;
    wire N__10922;
    wire N__10919;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10898;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10870;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10862;
    wire N__10859;
    wire N__10854;
    wire N__10849;
    wire N__10844;
    wire N__10843;
    wire N__10842;
    wire N__10839;
    wire N__10838;
    wire N__10835;
    wire N__10834;
    wire N__10831;
    wire N__10828;
    wire N__10823;
    wire N__10820;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10798;
    wire N__10797;
    wire N__10794;
    wire N__10793;
    wire N__10792;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10738;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10730;
    wire N__10729;
    wire N__10728;
    wire N__10727;
    wire N__10724;
    wire N__10719;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10681;
    wire N__10680;
    wire N__10677;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10640;
    wire N__10637;
    wire N__10636;
    wire N__10633;
    wire N__10632;
    wire N__10631;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10616;
    wire N__10613;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10591;
    wire N__10590;
    wire N__10589;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10577;
    wire N__10574;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10540;
    wire N__10539;
    wire N__10536;
    wire N__10531;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10519;
    wire N__10516;
    wire N__10515;
    wire N__10510;
    wire N__10507;
    wire N__10502;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10497;
    wire N__10496;
    wire N__10493;
    wire N__10484;
    wire N__10479;
    wire N__10472;
    wire N__10471;
    wire N__10466;
    wire N__10465;
    wire N__10464;
    wire N__10463;
    wire N__10462;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10454;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10443;
    wire N__10440;
    wire N__10435;
    wire N__10428;
    wire N__10423;
    wire N__10418;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10309;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10294;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10283;
    wire N__10282;
    wire N__10281;
    wire N__10274;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10251;
    wire N__10246;
    wire N__10243;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10231;
    wire N__10230;
    wire N__10225;
    wire N__10222;
    wire N__10217;
    wire N__10216;
    wire N__10215;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10203;
    wire N__10202;
    wire N__10199;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9730;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9715;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9433;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8803;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8733;
    wire N__8732;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8716;
    wire N__8713;
    wire N__8712;
    wire N__8707;
    wire N__8704;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8644;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8526;
    wire N__8521;
    wire N__8518;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8451;
    wire N__8446;
    wire N__8443;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8338;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7888;
    wire N__7887;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7877;
    wire N__7874;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7771;
    wire N__7770;
    wire N__7767;
    wire N__7766;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7738;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7713;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7666;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7647;
    wire N__7640;
    wire N__7637;
    wire N__7628;
    wire N__7625;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7615;
    wire N__7614;
    wire N__7611;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7580;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7548;
    wire N__7545;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7519;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7467;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5157;
    wire N__5156;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5144;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5125;
    wire N__5124;
    wire N__5119;
    wire N__5118;
    wire N__5117;
    wire N__5114;
    wire N__5113;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5086;
    wire N__5079;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5054;
    wire N__5051;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5043;
    wire N__5038;
    wire N__5037;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5029;
    wire N__5026;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5003;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4972;
    wire N__4963;
    wire N__4958;
    wire N__4955;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4945;
    wire N__4944;
    wire N__4941;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4927;
    wire N__4926;
    wire N__4921;
    wire N__4920;
    wire N__4919;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4882;
    wire N__4879;
    wire N__4878;
    wire N__4875;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4856;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4832;
    wire N__4829;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4817;
    wire N__4816;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4808;
    wire N__4805;
    wire N__4804;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4785;
    wire N__4784;
    wire N__4779;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4765;
    wire N__4760;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4744;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire write_data_c_5;
    wire write_data_c_4;
    wire write_data_c_3;
    wire write_data_c_2;
    wire write_data_c_1;
    wire write_data_c_0;
    wire write_address_c_9;
    wire write_address_c_8;
    wire write_address_c_7;
    wire write_address_c_6;
    wire write_address_c_5;
    wire write_address_c_4;
    wire write_address_c_3;
    wire write_address_c_2;
    wire write_address_c_10;
    wire write_address_c_1;
    wire write_address_c_0;
    wire VCCG0;
    wire this_vga_signals_N_170_i;
    wire this_vga_signals_N_171_i;
    wire rgb5_i;
    wire vsync_c;
    wire this_vga_signals_N_94_i;
    wire \this_vram.mem_out_bus0_0 ;
    wire \this_vram.mem_out_bus1_0 ;
    wire \this_vram.mem_out_bus0_2 ;
    wire \this_vram.mem_out_bus1_2 ;
    wire \this_vram.mem_out_bus0_3 ;
    wire \this_vram.mem_out_bus1_3 ;
    wire \this_vram.mem_out_bus0_4 ;
    wire \this_vram.mem_out_bus1_4 ;
    wire \this_vram.mem_out_bus1_5 ;
    wire \this_vram.mem_out_bus0_5 ;
    wire \this_vram.mem_out_bus3_0 ;
    wire \this_vram.mem_out_bus2_0 ;
    wire \this_vram.mem_mem_0_0_RNILGFZ0Z11 ;
    wire \this_vram.mem_mem_2_0_RNIPOJZ0Z11_cascade_ ;
    wire \this_vram.mem_N_2362 ;
    wire \this_vram.mem_N_2364_cascade_ ;
    wire M_this_vram_read_data_0;
    wire \this_vram.mem_out_bus3_3 ;
    wire \this_vram.mem_out_bus2_3 ;
    wire \this_vram.mem_mem_0_1_RNINGF11Z0Z_0 ;
    wire \this_vram.mem_mem_2_1_RNIROJ11Z0Z_0_cascade_ ;
    wire \this_vram.mem_out_bus4_3 ;
    wire \this_vram.mem_out_bus6_3 ;
    wire \this_vram.mem_mem_4_1_RNI14P11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_2336_cascade_ ;
    wire \this_vram.mem_N_2335 ;
    wire \this_vram.mem_out_bus3_2 ;
    wire \this_vram.mem_out_bus2_2 ;
    wire \this_vram.mem_mem_2_1_RNIROJZ0Z11_cascade_ ;
    wire \this_vram.mem_mem_0_1_RNINGFZ0Z11 ;
    wire \this_vram.mem_out_bus3_5 ;
    wire \this_vram.mem_out_bus2_5 ;
    wire \this_vram.mem_mem_0_2_RNIPGF11Z0Z_0 ;
    wire \this_vram.mem_mem_2_2_RNITOJ11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_2371_cascade_ ;
    wire \this_vram.mem_out_bus2_4 ;
    wire \this_vram.mem_out_bus3_4 ;
    wire \this_vram.mem_mem_0_2_RNIPGFZ0Z11 ;
    wire \this_vram.mem_mem_2_2_RNITOJZ0Z11_cascade_ ;
    wire \this_vram.mem_N_2326_cascade_ ;
    wire \this_vram.mem_N_2373 ;
    wire M_this_vram_read_data_5;
    wire \this_vram.mem_N_2328 ;
    wire M_this_vram_read_data_4;
    wire \this_vram.mem_N_2337 ;
    wire M_this_vram_read_data_3;
    wire \this_vram.mem_out_bus0_1 ;
    wire \this_vram.mem_out_bus1_1 ;
    wire \this_vram.mem_out_bus3_1 ;
    wire \this_vram.mem_out_bus2_1 ;
    wire \this_vram.mem_mem_0_0_RNILGF11Z0Z_0 ;
    wire \this_vram.mem_mem_2_0_RNIPOJ11Z0Z_0_cascade_ ;
    wire \this_vram.mem_out_bus6_0 ;
    wire \this_vram.mem_out_bus4_0 ;
    wire \this_vram.mem_WE_27 ;
    wire \this_vram.mem_out_bus5_0 ;
    wire \this_vram.mem_out_bus7_0 ;
    wire \this_vram.mem_mem_5_0_RNI18RZ0Z11_cascade_ ;
    wire \this_vram.mem_mem_4_0_RNIV3PZ0Z11 ;
    wire \this_vram.mem_N_2363 ;
    wire \this_vram.mem_N_2344 ;
    wire \this_vram.mem_N_2346 ;
    wire \this_vram.mem_G_25_0_cascade_ ;
    wire M_this_vram_read_data_2;
    wire \this_vram.mem_WE_21 ;
    wire \this_vram.mem_N_2327 ;
    wire \this_vram.mem_N_2353 ;
    wire \this_vram.mem_N_2355_cascade_ ;
    wire \this_vram.mem_G_25_0 ;
    wire M_this_vram_read_data_1;
    wire \this_vram.mem_out_bus4_4 ;
    wire \this_vram.mem_out_bus6_4 ;
    wire \this_vram.mem_mem_4_2_RNI34PZ0Z11 ;
    wire \this_vram.mem_WE_18 ;
    wire \this_vram.mem_out_bus6_1 ;
    wire \this_vram.mem_out_bus4_1 ;
    wire \this_vram.mem_out_bus5_1 ;
    wire \this_vram.mem_out_bus7_1 ;
    wire \this_vram.mem_mem_4_0_RNIV3P11Z0Z_0 ;
    wire \this_vram.mem_mem_5_0_RNI18R11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_2354 ;
    wire \this_vram.mem_WE_24 ;
    wire \this_vram.mem_out_bus4_2 ;
    wire \this_vram.mem_out_bus6_2 ;
    wire \this_vram.mem_mem_4_1_RNI14PZ0Z11_cascade_ ;
    wire \this_vram.mem_N_2345 ;
    wire \this_vram.mem_WE_15 ;
    wire \this_vga_signals.m24_0_1_cascade_ ;
    wire \this_vga_signals.N_25_cascade_ ;
    wire \this_vga_signals.m24_0_1_0 ;
    wire \this_vga_signals.m27_0_o2_1 ;
    wire \this_vga_signals.m27_0_0_cascade_ ;
    wire \this_vga_signals.i9_mux_cascade_ ;
    wire \this_vga_signals.N_40 ;
    wire M_this_vga_signals_address_7;
    wire bfn_13_15_0_;
    wire M_this_vga_signals_address_8;
    wire \this_vga_signals.address_1_cry_0 ;
    wire M_this_vga_signals_address_9;
    wire \this_vga_signals.address_1_cry_1 ;
    wire M_this_vga_signals_address_10;
    wire \this_vga_signals.address_1_cry_2 ;
    wire \this_vga_signals.address_1_cry_3 ;
    wire \this_vga_signals.address_1_cry_4 ;
    wire \this_vram.mem_radregZ0Z_13 ;
    wire \this_vga_signals.address_1_cry_5 ;
    wire \this_vga_signals.address_1_cry_6 ;
    wire \this_vram.mem_radregZ0Z_14 ;
    wire M_this_vga_signals_address_5;
    wire bfn_13_17_0_;
    wire M_this_vga_signals_address_6;
    wire \this_vga_signals.address_1_0_cry_0 ;
    wire \this_vga_signals.address_1 ;
    wire \this_vga_signals.address_1_0_cry_1 ;
    wire \this_vga_signals.address_1_0_3 ;
    wire \this_vga_signals.address_1_0_cry_2 ;
    wire \this_vga_signals.address_1_0_4 ;
    wire \this_vga_signals.address_1_0_cry_3 ;
    wire \this_vga_signals.address_1_0_5 ;
    wire \this_vga_signals.address_1_0_cry_4 ;
    wire \this_vga_signals.address_1_0_6 ;
    wire \this_vga_signals.address_1_0_cry_5 ;
    wire \this_vga_signals.address_1_0_7 ;
    wire \this_vga_signals.address_1_0_cry_6 ;
    wire \this_vga_signals.address_1_0_8 ;
    wire bfn_13_18_0_;
    wire \this_vga_signals.address_1_0_8_THRU_CO ;
    wire \this_vga_signals.m27_0_o2_0_3 ;
    wire \this_vga_signals.N_36 ;
    wire \this_vga_signals.m27_0_a2_1_5 ;
    wire \this_vga_signals.m27_0_a2_1_5_cascade_ ;
    wire \this_vga_signals.N_68_cascade_ ;
    wire \this_vga_signals.m27_0_a2_1_4 ;
    wire \this_vga_signals.M_vcounter_q_0_i_a2_0_0 ;
    wire \this_vga_signals.M_vstate_qZ0Z_0 ;
    wire \this_vga_signals.M_vstate_qZ0Z_1 ;
    wire \this_vga_signals.m24_0_0 ;
    wire bfn_14_15_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_14_16_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_9 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_10 ;
    wire \this_vga_signals.M_hstate_q_ns_i_i_1_0 ;
    wire \this_vga_signals.N_76_cascade_ ;
    wire \this_vga_signals.N_29_cascade_ ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire bfn_14_18_0_;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_0 ;
    wire \this_vga_signals.address_1_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_7 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_7 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_8 ;
    wire bfn_14_19_0_;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8 ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_0_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_1_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_2_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_3_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_4_THRU_CO ;
    wire GNDG0;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_5_THRU_CO ;
    wire \this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_6_THRU_CO ;
    wire \this_vga_signals.N_68 ;
    wire bfn_14_20_0_;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire N_112_g;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_hstate_qZ0Z_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_10 ;
    wire M_this_vga_signals_address_2;
    wire M_this_vga_signals_address_3;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.N_37_cascade_ ;
    wire \this_vga_signals.M_hstate_q_ns_i_i_2_0 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.M_hcounter_qZ0Z_11 ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.M_hstate_d_0_sqmuxa_0_a2_0_a2_0_cascade_ ;
    wire \this_vga_signals.N_169_4 ;
    wire \this_vga_signals.M_hstate_d_0_sqmuxa ;
    wire \this_vga_signals.N_169 ;
    wire \this_vga_signals.N_42 ;
    wire \this_vga_signals.N_46 ;
    wire \this_vga_signals.N_83 ;
    wire \this_vga_signals.M_hstate_qZ0Z_1 ;
    wire \this_vga_signals.N_27 ;
    wire M_this_reset_cond_out_0;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire clk_c_g;
    wire \this_vram.mem_out_bus6_5 ;
    wire \this_vram.mem_out_bus4_5 ;
    wire \this_vram.mem_mem_4_2_RNI34P11Z0Z_0_cascade_ ;
    wire \this_vram.mem_N_2372 ;
    wire \this_vram.mem_WE_12 ;
    wire CONSTANT_ONE_NET;
    wire \this_vram.mem_out_bus9_5 ;
    wire \this_vram.mem_out_bus8_5 ;
    wire \this_vram.mem_mem_8_2_RNI9H021Z0Z_0 ;
    wire \this_vram.mem_out_bus5_2 ;
    wire \this_vram.mem_out_bus7_2 ;
    wire \this_vram.mem_mem_5_1_RNI38RZ0Z11 ;
    wire \this_vram.mem_out_bus5_3 ;
    wire \this_vram.mem_out_bus7_3 ;
    wire \this_vram.mem_mem_5_1_RNI38R11Z0Z_0 ;
    wire \this_vram.mem_WE_9 ;
    wire \this_vram.mem_out_bus7_4 ;
    wire \this_vram.mem_out_bus5_4 ;
    wire \this_vram.mem_mem_5_2_RNI58RZ0Z11 ;
    wire \this_vram.mem_out_bus7_5 ;
    wire \this_vram.mem_radregZ0Z_12 ;
    wire \this_vram.mem_out_bus5_5 ;
    wire \this_vram.mem_mem_5_2_RNI58R11Z0Z_0 ;
    wire \this_vram.mem_WE_6 ;
    wire \this_vram.mem_out_bus9_0 ;
    wire \this_vram.mem_out_bus8_0 ;
    wire \this_vram.mem_mem_8_0_RNI5HZ0Z021 ;
    wire \this_vram.mem_out_bus8_1 ;
    wire \this_vram.mem_out_bus9_1 ;
    wire \this_vram.mem_mem_8_0_RNI5H021Z0Z_0 ;
    wire \this_vram.mem_out_bus8_2 ;
    wire \this_vram.mem_out_bus9_2 ;
    wire \this_vram.mem_mem_8_1_RNI7HZ0Z021 ;
    wire \this_vram.mem_N_27 ;
    wire \this_vram.mem_WE_0 ;
    wire write_address_c_13;
    wire write_address_c_12;
    wire \this_vram.mem_N_29 ;
    wire write_address_c_14;
    wire write_address_c_11;
    wire \this_vram.mem_N_29_cascade_ ;
    wire write_en_c;
    wire \this_vram.mem_WE_3 ;
    wire \this_vram.mem_out_bus9_3 ;
    wire \this_vram.mem_out_bus8_3 ;
    wire \this_vram.mem_mem_8_1_RNI7H021Z0Z_0 ;
    wire \this_vram.mem_radregZ0Z_11 ;
    wire \this_vram.mem_out_bus8_4 ;
    wire \this_vram.mem_out_bus9_4 ;
    wire \this_vram.mem_mem_8_2_RNI9HZ0Z021 ;
    wire _gnd_net_;

    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,\this_vram.mem_out_bus0_1 ,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,\this_vram.mem_out_bus0_0 ,dangling_wire_11,dangling_wire_12,dangling_wire_13}),
            .RADDR({N__9071,N__9290,N__9500,N__9707,N__9968,N__10175,N__11210,N__11447,N__11678,N__12464,N__12725}),
            .WADDR({N__5789,N__7460,N__7253,N__7043,N__6833,N__6623,N__6410,N__6203,N__5993,N__5582,N__5378}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,N__7758,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__7610,dangling_wire_41,dangling_wire_42,dangling_wire_43}),
            .RCLKE(),
            .RCLK(N__13655),
            .RE(N__13208),
            .WCLKE(N__8459),
            .WCLK(N__13656),
            .WE(N__13146));
    defparam \this_vram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,\this_vram.mem_out_bus0_3 ,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,\this_vram.mem_out_bus0_2 ,dangling_wire_55,dangling_wire_56,dangling_wire_57}),
            .RADDR({N__9064,N__9283,N__9494,N__9701,N__9962,N__10169,N__11204,N__11441,N__11672,N__12458,N__12719}),
            .WADDR({N__5783,N__7454,N__7247,N__7037,N__6827,N__6617,N__6404,N__6197,N__5987,N__5576,N__5372}),
            .MASK({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .WDATA({dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,N__4954,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,N__4832,dangling_wire_85,dangling_wire_86,dangling_wire_87}),
            .RCLKE(),
            .RCLK(N__13659),
            .RE(N__13171),
            .WCLKE(N__8458),
            .WCLK(N__13660),
            .WE(N__13131));
    defparam \this_vram.mem_mem_0_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_0_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_0_2_physical  (
            .RDATA({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,\this_vram.mem_out_bus0_5 ,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,\this_vram.mem_out_bus0_4 ,dangling_wire_99,dangling_wire_100,dangling_wire_101}),
            .RADDR({N__9052,N__9271,N__9488,N__9695,N__9956,N__10163,N__11198,N__11435,N__11666,N__12451,N__12713}),
            .WADDR({N__5777,N__7448,N__7240,N__7031,N__6821,N__6611,N__6398,N__6191,N__5977,N__5570,N__5362}),
            .MASK({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .WDATA({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__5124,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,N__5002,dangling_wire_129,dangling_wire_130,dangling_wire_131}),
            .RCLKE(),
            .RCLK(N__13663),
            .RE(N__13016),
            .WCLKE(N__8451),
            .WCLK(N__13664),
            .WE(N__13110));
    defparam \this_vram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,\this_vram.mem_out_bus1_1 ,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,\this_vram.mem_out_bus1_0 ,dangling_wire_143,dangling_wire_144,dangling_wire_145}),
            .RADDR({N__9040,N__9259,N__9478,N__9685,N__9946,N__10153,N__11191,N__11428,N__11660,N__12439,N__12703}),
            .WADDR({N__5767,N__7442,N__7228,N__7021,N__6815,N__6605,N__6391,N__6184,N__5965,N__5564,N__5350}),
            .MASK({dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161}),
            .WDATA({dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__7765,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,N__7580,dangling_wire_173,dangling_wire_174,dangling_wire_175}),
            .RCLKE(),
            .RCLK(N__13667),
            .RE(N__13194),
            .WCLKE(N__8534),
            .WCLK(N__13668),
            .WE(N__13114));
    defparam \this_vram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,\this_vram.mem_out_bus1_3 ,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,\this_vram.mem_out_bus1_2 ,dangling_wire_187,dangling_wire_188,dangling_wire_189}),
            .RADDR({N__9028,N__9247,N__9466,N__9673,N__9934,N__10141,N__11179,N__11416,N__11650,N__12427,N__12691}),
            .WADDR({N__5755,N__7432,N__7216,N__7009,N__6805,N__6595,N__6379,N__6172,N__5953,N__5557,N__5338}),
            .MASK({dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205}),
            .WDATA({dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,N__4940,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,N__4828,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .RCLKE(),
            .RCLK(N__13675),
            .RE(N__13265),
            .WCLKE(N__8533),
            .WCLK(N__13674),
            .WE(N__13172));
    defparam \this_vram.mem_mem_1_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_1_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_1_2_physical  (
            .RDATA({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,\this_vram.mem_out_bus1_5 ,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,\this_vram.mem_out_bus1_4 ,dangling_wire_231,dangling_wire_232,dangling_wire_233}),
            .RADDR({N__9016,N__9235,N__9454,N__9661,N__9922,N__10129,N__11167,N__11404,N__11638,N__12415,N__12679}),
            .WADDR({N__5743,N__7420,N__7204,N__6997,N__6793,N__6583,N__6367,N__6160,N__5941,N__5545,N__5326}),
            .MASK({dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249}),
            .WDATA({dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,N__5113,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,N__5003,dangling_wire_261,dangling_wire_262,dangling_wire_263}),
            .RCLKE(),
            .RCLK(N__13683),
            .RE(N__13266),
            .WCLKE(N__8526),
            .WCLK(N__13684),
            .WE(N__13173));
    defparam \this_vram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,\this_vram.mem_out_bus2_1 ,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,\this_vram.mem_out_bus2_0 ,dangling_wire_275,dangling_wire_276,dangling_wire_277}),
            .RADDR({N__9004,N__9223,N__9442,N__9649,N__9910,N__10117,N__11155,N__11392,N__11626,N__12403,N__12667}),
            .WADDR({N__5731,N__7408,N__7192,N__6985,N__6781,N__6571,N__6355,N__6148,N__5929,N__5533,N__5314}),
            .MASK({dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293}),
            .WDATA({dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,N__7738,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,N__7590,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .RCLKE(),
            .RCLK(N__13690),
            .RE(N__13237),
            .WCLKE(N__8342),
            .WCLK(N__13691),
            .WE(N__13238));
    defparam \this_vram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,\this_vram.mem_out_bus2_3 ,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,\this_vram.mem_out_bus2_2 ,dangling_wire_319,dangling_wire_320,dangling_wire_321}),
            .RADDR({N__8992,N__9211,N__9430,N__9637,N__9898,N__10105,N__11143,N__11380,N__11614,N__12391,N__12655}),
            .WADDR({N__5719,N__7396,N__7180,N__6973,N__6769,N__6559,N__6343,N__6136,N__5917,N__5521,N__5302}),
            .MASK({dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337}),
            .WDATA({dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,N__4927,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,N__4816,dangling_wire_349,dangling_wire_350,dangling_wire_351}),
            .RCLKE(),
            .RCLK(N__13696),
            .RE(N__13332),
            .WCLKE(N__8338),
            .WCLK(N__13697),
            .WE(N__13239));
    defparam \this_vram.mem_mem_2_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_2_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_2_2_physical  (
            .RDATA({dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,\this_vram.mem_out_bus2_5 ,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,\this_vram.mem_out_bus2_4 ,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .RADDR({N__8980,N__9199,N__9418,N__9625,N__9886,N__10093,N__11131,N__11368,N__11602,N__12379,N__12643}),
            .WADDR({N__5707,N__7384,N__7168,N__6961,N__6757,N__6547,N__6331,N__6124,N__5905,N__5509,N__5290}),
            .MASK({dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381}),
            .WDATA({dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,N__5112,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,N__5036,dangling_wire_393,dangling_wire_394,dangling_wire_395}),
            .RCLKE(),
            .RCLK(N__13700),
            .RE(N__13379),
            .WCLKE(N__8337),
            .WCLK(N__13701),
            .WE(N__13300));
    defparam \this_vram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,\this_vram.mem_out_bus3_1 ,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,\this_vram.mem_out_bus3_0 ,dangling_wire_407,dangling_wire_408,dangling_wire_409}),
            .RADDR({N__8968,N__9187,N__9406,N__9613,N__9874,N__10081,N__11119,N__11356,N__11590,N__12367,N__12631}),
            .WADDR({N__5695,N__7372,N__7156,N__6949,N__6745,N__6535,N__6319,N__6112,N__5893,N__5497,N__5278}),
            .MASK({dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425}),
            .WDATA({dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,N__7748,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,N__7565,dangling_wire_437,dangling_wire_438,dangling_wire_439}),
            .RCLKE(),
            .RCLK(N__13704),
            .RE(N__13380),
            .WCLKE(N__8643),
            .WCLK(N__13705),
            .WE(N__13301));
    defparam \this_vram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,\this_vram.mem_out_bus3_3 ,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,\this_vram.mem_out_bus3_2 ,dangling_wire_451,dangling_wire_452,dangling_wire_453}),
            .RADDR({N__8956,N__9175,N__9394,N__9601,N__9862,N__10069,N__11107,N__11344,N__11578,N__12355,N__12619}),
            .WADDR({N__5683,N__7360,N__7144,N__6937,N__6733,N__6523,N__6307,N__6100,N__5881,N__5485,N__5266}),
            .MASK({dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469}),
            .WDATA({dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,N__4907,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,N__4808,dangling_wire_481,dangling_wire_482,dangling_wire_483}),
            .RCLKE(),
            .RCLK(N__13708),
            .RE(N__13352),
            .WCLKE(N__8644),
            .WCLK(N__13709),
            .WE(N__13353));
    defparam \this_vram.mem_mem_3_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_3_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_3_2_physical  (
            .RDATA({dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,\this_vram.mem_out_bus3_5 ,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,\this_vram.mem_out_bus3_4 ,dangling_wire_495,dangling_wire_496,dangling_wire_497}),
            .RADDR({N__8944,N__9163,N__9382,N__9589,N__9850,N__10057,N__11095,N__11332,N__11566,N__12343,N__12607}),
            .WADDR({N__5671,N__7348,N__7132,N__6925,N__6721,N__6511,N__6295,N__6088,N__5869,N__5473,N__5254}),
            .MASK({dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513}),
            .WDATA({dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,N__5117,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,N__5025,dangling_wire_525,dangling_wire_526,dangling_wire_527}),
            .RCLKE(),
            .RCLK(N__13712),
            .RE(N__13378),
            .WCLKE(N__8648),
            .WCLK(N__13713),
            .WE(N__13354));
    defparam \this_vram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,\this_vram.mem_out_bus4_1 ,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,\this_vram.mem_out_bus4_0 ,dangling_wire_539,dangling_wire_540,dangling_wire_541}),
            .RADDR({N__8932,N__9151,N__9370,N__9577,N__9838,N__10045,N__11083,N__11320,N__11554,N__12331,N__12595}),
            .WADDR({N__5659,N__7336,N__7120,N__6913,N__6709,N__6499,N__6283,N__6076,N__5857,N__5461,N__5242}),
            .MASK({dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557}),
            .WDATA({dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,N__7713,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,N__7533,dangling_wire_569,dangling_wire_570,dangling_wire_571}),
            .RCLKE(),
            .RCLK(N__13716),
            .RE(N__13384),
            .WCLKE(N__8802),
            .WCLK(N__13717),
            .WE(N__13385));
    defparam \this_vram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,\this_vram.mem_out_bus4_3 ,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,\this_vram.mem_out_bus4_2 ,dangling_wire_583,dangling_wire_584,dangling_wire_585}),
            .RADDR({N__8920,N__9139,N__9358,N__9565,N__9826,N__10033,N__11071,N__11308,N__11542,N__12319,N__12583}),
            .WADDR({N__5647,N__7324,N__7108,N__6901,N__6697,N__6487,N__6271,N__6064,N__5845,N__5449,N__5230}),
            .MASK({dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601}),
            .WDATA({dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,N__4926,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,N__4784,dangling_wire_613,dangling_wire_614,dangling_wire_615}),
            .RCLKE(),
            .RCLK(N__13720),
            .RE(N__13396),
            .WCLKE(N__8803),
            .WCLK(N__13721),
            .WE(N__13386));
    defparam \this_vram.mem_mem_4_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_4_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_4_2_physical  (
            .RDATA({dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,\this_vram.mem_out_bus4_5 ,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,\this_vram.mem_out_bus4_4 ,dangling_wire_627,dangling_wire_628,dangling_wire_629}),
            .RADDR({N__8908,N__9127,N__9346,N__9553,N__9814,N__10021,N__11059,N__11296,N__11530,N__12307,N__12571}),
            .WADDR({N__5635,N__7312,N__7096,N__6889,N__6685,N__6475,N__6259,N__6052,N__5833,N__5437,N__5218}),
            .MASK({dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645}),
            .WDATA({dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,N__5118,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,N__5037,dangling_wire_657,dangling_wire_658,dangling_wire_659}),
            .RCLKE(),
            .RCLK(N__13724),
            .RE(N__13400),
            .WCLKE(N__8807),
            .WCLK(N__13725),
            .WE(N__13401));
    defparam \this_vram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,\this_vram.mem_out_bus5_1 ,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,\this_vram.mem_out_bus5_0 ,dangling_wire_671,dangling_wire_672,dangling_wire_673}),
            .RADDR({N__8896,N__9115,N__9334,N__9541,N__9802,N__10009,N__11047,N__11284,N__11518,N__12295,N__12559}),
            .WADDR({N__5623,N__7300,N__7084,N__6877,N__6673,N__6463,N__6247,N__6040,N__5821,N__5425,N__5206}),
            .MASK({dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689}),
            .WDATA({dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,N__7712,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,N__7509,dangling_wire_701,dangling_wire_702,dangling_wire_703}),
            .RCLKE(),
            .RCLK(N__13726),
            .RE(N__13403),
            .WCLKE(N__13446),
            .WCLK(N__13727),
            .WE(N__13402));
    defparam \this_vram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,\this_vram.mem_out_bus5_3 ,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,\this_vram.mem_out_bus5_2 ,dangling_wire_715,dangling_wire_716,dangling_wire_717}),
            .RADDR({N__9067,N__9286,N__9487,N__9694,N__9955,N__10162,N__11194,N__11431,N__11659,N__12454,N__12712}),
            .WADDR({N__5776,N__7441,N__7243,N__7030,N__6814,N__6604,N__6394,N__6187,N__5986,N__5560,N__5371}),
            .MASK({dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733}),
            .WDATA({dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,N__4955,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,N__4815,dangling_wire_745,dangling_wire_746,dangling_wire_747}),
            .RCLKE(),
            .RCLK(N__13657),
            .RE(N__13049),
            .WCLKE(N__13451),
            .WCLK(N__13658),
            .WE(N__12997));
    defparam \this_vram.mem_mem_5_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_5_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_5_2_physical  (
            .RDATA({dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,\this_vram.mem_out_bus5_5 ,dangling_wire_752,dangling_wire_753,dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,dangling_wire_758,\this_vram.mem_out_bus5_4 ,dangling_wire_759,dangling_wire_760,dangling_wire_761}),
            .RADDR({N__9055,N__9274,N__9475,N__9682,N__9943,N__10150,N__11182,N__11419,N__11647,N__12442,N__12700}),
            .WADDR({N__5764,N__7429,N__7231,N__7018,N__6802,N__6592,N__6382,N__6175,N__5974,N__5548,N__5359}),
            .MASK({dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,dangling_wire_767,dangling_wire_768,dangling_wire_769,dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777}),
            .WDATA({dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,N__5171,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785,dangling_wire_786,dangling_wire_787,dangling_wire_788,N__5029,dangling_wire_789,dangling_wire_790,dangling_wire_791}),
            .RCLKE(),
            .RCLK(N__13661),
            .RE(N__12979),
            .WCLKE(N__13447),
            .WCLK(N__13662),
            .WE(N__12993));
    defparam \this_vram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,\this_vram.mem_out_bus6_1 ,dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,dangling_wire_802,\this_vram.mem_out_bus6_0 ,dangling_wire_803,dangling_wire_804,dangling_wire_805}),
            .RADDR({N__9043,N__9262,N__9463,N__9670,N__9931,N__10138,N__11170,N__11407,N__11635,N__12430,N__12688}),
            .WADDR({N__5752,N__7417,N__7219,N__7006,N__6790,N__6580,N__6370,N__6163,N__5962,N__5536,N__5347}),
            .MASK({dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,dangling_wire_811,dangling_wire_812,dangling_wire_813,dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821}),
            .WDATA({dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,N__7772,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,N__7628,dangling_wire_833,dangling_wire_834,dangling_wire_835}),
            .RCLKE(),
            .RCLK(N__13665),
            .RE(N__12897),
            .WCLKE(N__14255),
            .WCLK(N__13666),
            .WE(N__12934));
    defparam \this_vram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,\this_vram.mem_out_bus6_3 ,dangling_wire_840,dangling_wire_841,dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,dangling_wire_846,\this_vram.mem_out_bus6_2 ,dangling_wire_847,dangling_wire_848,dangling_wire_849}),
            .RADDR({N__9031,N__9250,N__9451,N__9658,N__9919,N__10126,N__11158,N__11395,N__11623,N__12418,N__12676}),
            .WADDR({N__5740,N__7405,N__7207,N__6994,N__6778,N__6568,N__6358,N__6151,N__5950,N__5524,N__5335}),
            .MASK({dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,dangling_wire_855,dangling_wire_856,dangling_wire_857,dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865}),
            .WDATA({dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,N__4944,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873,dangling_wire_874,dangling_wire_875,dangling_wire_876,N__4804,dangling_wire_877,dangling_wire_878,dangling_wire_879}),
            .RCLKE(),
            .RCLK(N__13670),
            .RE(N__12954),
            .WCLKE(N__14254),
            .WCLK(N__13671),
            .WE(N__13030));
    defparam \this_vram.mem_mem_6_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_6_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_6_2_physical  (
            .RDATA({dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,\this_vram.mem_out_bus6_5 ,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889,dangling_wire_890,\this_vram.mem_out_bus6_4 ,dangling_wire_891,dangling_wire_892,dangling_wire_893}),
            .RADDR({N__9019,N__9238,N__9439,N__9646,N__9907,N__10114,N__11146,N__11383,N__11611,N__12406,N__12664}),
            .WADDR({N__5728,N__7393,N__7195,N__6982,N__6766,N__6556,N__6346,N__6139,N__5938,N__5512,N__5323}),
            .MASK({dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,dangling_wire_899,dangling_wire_900,dangling_wire_901,dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909}),
            .WDATA({dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,N__5164,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917,dangling_wire_918,dangling_wire_919,dangling_wire_920,N__5050,dangling_wire_921,dangling_wire_922,dangling_wire_923}),
            .RCLKE(),
            .RCLK(N__13680),
            .RE(N__12955),
            .WCLKE(N__14247),
            .WCLK(N__13679),
            .WE(N__13087));
    defparam \this_vram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,\this_vram.mem_out_bus7_1 ,dangling_wire_928,dangling_wire_929,dangling_wire_930,dangling_wire_931,dangling_wire_932,dangling_wire_933,dangling_wire_934,\this_vram.mem_out_bus7_0 ,dangling_wire_935,dangling_wire_936,dangling_wire_937}),
            .RADDR({N__9007,N__9226,N__9427,N__9634,N__9895,N__10102,N__11134,N__11371,N__11599,N__12394,N__12652}),
            .WADDR({N__5716,N__7381,N__7183,N__6970,N__6754,N__6544,N__6334,N__6127,N__5926,N__5500,N__5311}),
            .MASK({dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,dangling_wire_943,dangling_wire_944,dangling_wire_945,dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953}),
            .WDATA({dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,N__7771,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961,dangling_wire_962,dangling_wire_963,dangling_wire_964,N__7624,dangling_wire_965,dangling_wire_966,dangling_wire_967}),
            .RCLKE(),
            .RCLK(N__13686),
            .RE(N__13149),
            .WCLKE(N__13994),
            .WCLK(N__13687),
            .WE(N__13088));
    defparam \this_vram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,\this_vram.mem_out_bus7_3 ,dangling_wire_972,dangling_wire_973,dangling_wire_974,dangling_wire_975,dangling_wire_976,dangling_wire_977,dangling_wire_978,\this_vram.mem_out_bus7_2 ,dangling_wire_979,dangling_wire_980,dangling_wire_981}),
            .RADDR({N__8995,N__9214,N__9415,N__9622,N__9883,N__10090,N__11122,N__11359,N__11587,N__12382,N__12640}),
            .WADDR({N__5704,N__7369,N__7171,N__6958,N__6742,N__6532,N__6322,N__6115,N__5914,N__5488,N__5299}),
            .MASK({dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,dangling_wire_987,dangling_wire_988,dangling_wire_989,dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997}),
            .WDATA({dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,N__4920,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005,dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,N__4778,dangling_wire_1009,dangling_wire_1010,dangling_wire_1011}),
            .RCLKE(),
            .RCLK(N__13694),
            .RE(N__13150),
            .WCLKE(N__13993),
            .WCLK(N__13695),
            .WE(N__13147));
    defparam \this_vram.mem_mem_7_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_7_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_7_2_physical  (
            .RDATA({dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,\this_vram.mem_out_bus7_5 ,dangling_wire_1016,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019,dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,\this_vram.mem_out_bus7_4 ,dangling_wire_1023,dangling_wire_1024,dangling_wire_1025}),
            .RADDR({N__8983,N__9202,N__9403,N__9610,N__9871,N__10078,N__11110,N__11347,N__11575,N__12370,N__12628}),
            .WADDR({N__5692,N__7357,N__7159,N__6946,N__6730,N__6520,N__6310,N__6103,N__5902,N__5476,N__5287}),
            .MASK({dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033,dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041}),
            .WDATA({dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,N__5157,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049,dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,N__5043,dangling_wire_1053,dangling_wire_1054,dangling_wire_1055}),
            .RCLKE(),
            .RCLK(N__13698),
            .RE(N__13209),
            .WCLKE(N__13992),
            .WCLK(N__13699),
            .WE(N__13148));
    defparam \this_vram.mem_mem_8_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_8_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_8_0_physical  (
            .RDATA({dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,\this_vram.mem_out_bus8_1 ,dangling_wire_1060,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063,dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,\this_vram.mem_out_bus8_0 ,dangling_wire_1067,dangling_wire_1068,dangling_wire_1069}),
            .RADDR({N__8971,N__9190,N__9391,N__9598,N__9859,N__10066,N__11098,N__11335,N__11563,N__12358,N__12616}),
            .WADDR({N__5680,N__7345,N__7147,N__6934,N__6718,N__6508,N__6298,N__6091,N__5890,N__5464,N__5275}),
            .MASK({dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077,dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085}),
            .WDATA({dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,N__7766,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093,dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,N__7614,dangling_wire_1097,dangling_wire_1098,dangling_wire_1099}),
            .RCLKE(),
            .RCLK(N__13702),
            .RE(N__13210),
            .WCLKE(N__14543),
            .WCLK(N__13703),
            .WE(N__13276));
    defparam \this_vram.mem_mem_8_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_8_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_8_1_physical  (
            .RDATA({dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,\this_vram.mem_out_bus8_3 ,dangling_wire_1104,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107,dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,\this_vram.mem_out_bus8_2 ,dangling_wire_1111,dangling_wire_1112,dangling_wire_1113}),
            .RADDR({N__8959,N__9178,N__9379,N__9586,N__9847,N__10054,N__11086,N__11323,N__11551,N__12346,N__12604}),
            .WADDR({N__5668,N__7333,N__7135,N__6922,N__6706,N__6496,N__6286,N__6079,N__5878,N__5452,N__5263}),
            .MASK({dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121,dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129}),
            .WDATA({dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,N__4878,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137,dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,N__4765,dangling_wire_1141,dangling_wire_1142,dangling_wire_1143}),
            .RCLKE(),
            .RCLK(N__13706),
            .RE(N__13278),
            .WCLKE(N__14535),
            .WCLK(N__13707),
            .WE(N__13277));
    defparam \this_vram.mem_mem_8_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_8_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_8_2_physical  (
            .RDATA({dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,\this_vram.mem_out_bus8_5 ,dangling_wire_1148,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151,dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,\this_vram.mem_out_bus8_4 ,dangling_wire_1155,dangling_wire_1156,dangling_wire_1157}),
            .RADDR({N__8947,N__9166,N__9367,N__9574,N__9835,N__10042,N__11074,N__11311,N__11539,N__12334,N__12592}),
            .WADDR({N__5656,N__7321,N__7123,N__6910,N__6694,N__6484,N__6274,N__6067,N__5866,N__5440,N__5251}),
            .MASK({dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165,dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173}),
            .WDATA({dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,N__5144,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181,dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,N__5065,dangling_wire_1185,dangling_wire_1186,dangling_wire_1187}),
            .RCLKE(),
            .RCLK(N__13710),
            .RE(N__13279),
            .WCLKE(N__14542),
            .WCLK(N__13711),
            .WE(N__13339));
    defparam \this_vram.mem_mem_9_0_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_9_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_9_0_physical  (
            .RDATA({dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,\this_vram.mem_out_bus9_1 ,dangling_wire_1192,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195,dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,\this_vram.mem_out_bus9_0 ,dangling_wire_1199,dangling_wire_1200,dangling_wire_1201}),
            .RADDR({N__8935,N__9154,N__9355,N__9562,N__9823,N__10030,N__11062,N__11299,N__11527,N__12322,N__12580}),
            .WADDR({N__5644,N__7309,N__7111,N__6898,N__6682,N__6472,N__6262,N__6055,N__5854,N__5428,N__5239}),
            .MASK({dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209,dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217}),
            .WDATA({dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,N__7770,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225,dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,N__7600,dangling_wire_1229,dangling_wire_1230,dangling_wire_1231}),
            .RCLKE(),
            .RCLK(N__13714),
            .RE(N__13347),
            .WCLKE(N__14919),
            .WCLK(N__13715),
            .WE(N__13340));
    defparam \this_vram.mem_mem_9_1_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_9_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_9_1_physical  (
            .RDATA({dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,\this_vram.mem_out_bus9_3 ,dangling_wire_1236,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239,dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,\this_vram.mem_out_bus9_2 ,dangling_wire_1243,dangling_wire_1244,dangling_wire_1245}),
            .RADDR({N__8923,N__9142,N__9343,N__9550,N__9811,N__10018,N__11050,N__11287,N__11515,N__12310,N__12568}),
            .WADDR({N__5632,N__7297,N__7099,N__6886,N__6670,N__6460,N__6250,N__6043,N__5842,N__5416,N__5227}),
            .MASK({dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253,dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261}),
            .WDATA({dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,N__4919,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269,dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,N__4743,dangling_wire_1273,dangling_wire_1274,dangling_wire_1275}),
            .RCLKE(),
            .RCLK(N__13718),
            .RE(N__13348),
            .WCLKE(N__14926),
            .WCLK(N__13719),
            .WE(N__13381));
    defparam \this_vram.mem_mem_9_2_physical .WRITE_MODE=3;
    defparam \this_vram.mem_mem_9_2_physical .READ_MODE=3;
    SB_RAM40_4K \this_vram.mem_mem_9_2_physical  (
            .RDATA({dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,\this_vram.mem_out_bus9_5 ,dangling_wire_1280,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283,dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,\this_vram.mem_out_bus9_4 ,dangling_wire_1287,dangling_wire_1288,dangling_wire_1289}),
            .RADDR({N__8911,N__9130,N__9331,N__9538,N__9799,N__10006,N__11038,N__11275,N__11503,N__12298,N__12556}),
            .WADDR({N__5620,N__7285,N__7087,N__6874,N__6658,N__6448,N__6238,N__6031,N__5830,N__5404,N__5215}),
            .MASK({dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297,dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305}),
            .WDATA({dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,N__5156,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313,dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,N__5069,dangling_wire_1317,dangling_wire_1318,dangling_wire_1319}),
            .RCLKE(),
            .RCLK(N__13722),
            .RE(N__13383),
            .WCLKE(N__14927),
            .WCLK(N__13723),
            .WE(N__13382));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__15243),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__15245),
            .DIN(N__15244),
            .DOUT(N__15243),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__15245),
            .PADOUT(N__15244),
            .PADIN(N__15243),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__15234),
            .DIN(N__15233),
            .DOUT(N__15232),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__15234),
            .PADOUT(N__15233),
            .PADIN(N__15232),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7898),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__15225),
            .DIN(N__15224),
            .DOUT(N__15223),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__15225),
            .PADOUT(N__15224),
            .PADIN(N__15223),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7910),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuft_0_iopad (
            .OE(N__15216),
            .DIN(N__15215),
            .DOUT(N__15214),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO rgb_obuft_0_preio (
            .PADOEN(N__15216),
            .PADOUT(N__15215),
            .PADIN(N__15214),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7940),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__7892));
    IO_PAD rgb_obuft_1_iopad (
            .OE(N__15207),
            .DIN(N__15206),
            .DOUT(N__15205),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO rgb_obuft_1_preio (
            .PADOEN(N__15207),
            .PADOUT(N__15206),
            .PADIN(N__15205),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8699),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__7845));
    IO_PAD rgb_obuft_2_iopad (
            .OE(N__15198),
            .DIN(N__15197),
            .DOUT(N__15196),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO rgb_obuft_2_preio (
            .PADOEN(N__15198),
            .PADOUT(N__15197),
            .PADIN(N__15196),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8351),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__7846));
    IO_PAD rgb_obuft_3_iopad (
            .OE(N__15189),
            .DIN(N__15188),
            .DOUT(N__15187),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO rgb_obuft_3_preio (
            .PADOEN(N__15189),
            .PADOUT(N__15188),
            .PADIN(N__15187),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8216),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__7877));
    IO_PAD rgb_obuft_4_iopad (
            .OE(N__15180),
            .DIN(N__15179),
            .DOUT(N__15178),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO rgb_obuft_4_preio (
            .PADOEN(N__15180),
            .PADOUT(N__15179),
            .PADIN(N__15178),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8243),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__7888));
    IO_PAD rgb_obuft_5_iopad (
            .OE(N__15171),
            .DIN(N__15170),
            .DOUT(N__15169),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO rgb_obuft_5_preio (
            .PADOEN(N__15171),
            .PADOUT(N__15170),
            .PADIN(N__15169),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__8270),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__7887));
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__15162),
            .DIN(N__15161),
            .DOUT(N__15160),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__15162),
            .PADOUT(N__15161),
            .PADIN(N__15160),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__15153),
            .DIN(N__15152),
            .DOUT(N__15151),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__15153),
            .PADOUT(N__15152),
            .PADIN(N__15151),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7823),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__15144),
            .DIN(N__15143),
            .DOUT(N__15142),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__15144),
            .PADOUT(N__15143),
            .PADIN(N__15142),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__7829),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_0_iopad (
            .OE(N__15135),
            .DIN(N__15134),
            .DOUT(N__15133),
            .PACKAGEPIN(write_address[0]));
    defparam write_address_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_0_preio (
            .PADOEN(N__15135),
            .PADOUT(N__15134),
            .PADIN(N__15133),
            .CLOCKENABLE(),
            .DIN0(write_address_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_1_iopad (
            .OE(N__15126),
            .DIN(N__15125),
            .DOUT(N__15124),
            .PACKAGEPIN(write_address[1]));
    defparam write_address_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_1_preio (
            .PADOEN(N__15126),
            .PADOUT(N__15125),
            .PADIN(N__15124),
            .CLOCKENABLE(),
            .DIN0(write_address_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_10_iopad (
            .OE(N__15117),
            .DIN(N__15116),
            .DOUT(N__15115),
            .PACKAGEPIN(write_address[10]));
    defparam write_address_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_10_preio (
            .PADOEN(N__15117),
            .PADOUT(N__15116),
            .PADIN(N__15115),
            .CLOCKENABLE(),
            .DIN0(write_address_c_10),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_11_iopad (
            .OE(N__15108),
            .DIN(N__15107),
            .DOUT(N__15106),
            .PACKAGEPIN(write_address[11]));
    defparam write_address_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_11_preio (
            .PADOEN(N__15108),
            .PADOUT(N__15107),
            .PADIN(N__15106),
            .CLOCKENABLE(),
            .DIN0(write_address_c_11),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_12_iopad (
            .OE(N__15099),
            .DIN(N__15098),
            .DOUT(N__15097),
            .PACKAGEPIN(write_address[12]));
    defparam write_address_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_12_preio (
            .PADOEN(N__15099),
            .PADOUT(N__15098),
            .PADIN(N__15097),
            .CLOCKENABLE(),
            .DIN0(write_address_c_12),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_13_iopad (
            .OE(N__15090),
            .DIN(N__15089),
            .DOUT(N__15088),
            .PACKAGEPIN(write_address[13]));
    defparam write_address_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_13_preio (
            .PADOEN(N__15090),
            .PADOUT(N__15089),
            .PADIN(N__15088),
            .CLOCKENABLE(),
            .DIN0(write_address_c_13),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_14_iopad (
            .OE(N__15081),
            .DIN(N__15080),
            .DOUT(N__15079),
            .PACKAGEPIN(write_address[14]));
    defparam write_address_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_14_preio (
            .PADOEN(N__15081),
            .PADOUT(N__15080),
            .PADIN(N__15079),
            .CLOCKENABLE(),
            .DIN0(write_address_c_14),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_2_iopad (
            .OE(N__15072),
            .DIN(N__15071),
            .DOUT(N__15070),
            .PACKAGEPIN(write_address[2]));
    defparam write_address_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_2_preio (
            .PADOEN(N__15072),
            .PADOUT(N__15071),
            .PADIN(N__15070),
            .CLOCKENABLE(),
            .DIN0(write_address_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_3_iopad (
            .OE(N__15063),
            .DIN(N__15062),
            .DOUT(N__15061),
            .PACKAGEPIN(write_address[3]));
    defparam write_address_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_3_preio (
            .PADOEN(N__15063),
            .PADOUT(N__15062),
            .PADIN(N__15061),
            .CLOCKENABLE(),
            .DIN0(write_address_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_4_iopad (
            .OE(N__15054),
            .DIN(N__15053),
            .DOUT(N__15052),
            .PACKAGEPIN(write_address[4]));
    defparam write_address_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_4_preio (
            .PADOEN(N__15054),
            .PADOUT(N__15053),
            .PADIN(N__15052),
            .CLOCKENABLE(),
            .DIN0(write_address_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_5_iopad (
            .OE(N__15045),
            .DIN(N__15044),
            .DOUT(N__15043),
            .PACKAGEPIN(write_address[5]));
    defparam write_address_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_5_preio (
            .PADOEN(N__15045),
            .PADOUT(N__15044),
            .PADIN(N__15043),
            .CLOCKENABLE(),
            .DIN0(write_address_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_6_iopad (
            .OE(N__15036),
            .DIN(N__15035),
            .DOUT(N__15034),
            .PACKAGEPIN(write_address[6]));
    defparam write_address_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_6_preio (
            .PADOEN(N__15036),
            .PADOUT(N__15035),
            .PADIN(N__15034),
            .CLOCKENABLE(),
            .DIN0(write_address_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_7_iopad (
            .OE(N__15027),
            .DIN(N__15026),
            .DOUT(N__15025),
            .PACKAGEPIN(write_address[7]));
    defparam write_address_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_7_preio (
            .PADOEN(N__15027),
            .PADOUT(N__15026),
            .PADIN(N__15025),
            .CLOCKENABLE(),
            .DIN0(write_address_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_8_iopad (
            .OE(N__15018),
            .DIN(N__15017),
            .DOUT(N__15016),
            .PACKAGEPIN(write_address[8]));
    defparam write_address_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_8_preio (
            .PADOEN(N__15018),
            .PADOUT(N__15017),
            .PADIN(N__15016),
            .CLOCKENABLE(),
            .DIN0(write_address_c_8),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_address_ibuf_9_iopad (
            .OE(N__15009),
            .DIN(N__15008),
            .DOUT(N__15007),
            .PACKAGEPIN(write_address[9]));
    defparam write_address_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam write_address_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO write_address_ibuf_9_preio (
            .PADOEN(N__15009),
            .PADOUT(N__15008),
            .PADIN(N__15007),
            .CLOCKENABLE(),
            .DIN0(write_address_c_9),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_data_ibuf_0_iopad (
            .OE(N__15000),
            .DIN(N__14999),
            .DOUT(N__14998),
            .PACKAGEPIN(write_data[0]));
    defparam write_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam write_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO write_data_ibuf_0_preio (
            .PADOEN(N__15000),
            .PADOUT(N__14999),
            .PADIN(N__14998),
            .CLOCKENABLE(),
            .DIN0(write_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_data_ibuf_1_iopad (
            .OE(N__14991),
            .DIN(N__14990),
            .DOUT(N__14989),
            .PACKAGEPIN(write_data[1]));
    defparam write_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam write_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO write_data_ibuf_1_preio (
            .PADOEN(N__14991),
            .PADOUT(N__14990),
            .PADIN(N__14989),
            .CLOCKENABLE(),
            .DIN0(write_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_data_ibuf_2_iopad (
            .OE(N__14982),
            .DIN(N__14981),
            .DOUT(N__14980),
            .PACKAGEPIN(write_data[2]));
    defparam write_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam write_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO write_data_ibuf_2_preio (
            .PADOEN(N__14982),
            .PADOUT(N__14981),
            .PADIN(N__14980),
            .CLOCKENABLE(),
            .DIN0(write_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_data_ibuf_3_iopad (
            .OE(N__14973),
            .DIN(N__14972),
            .DOUT(N__14971),
            .PACKAGEPIN(write_data[3]));
    defparam write_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam write_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO write_data_ibuf_3_preio (
            .PADOEN(N__14973),
            .PADOUT(N__14972),
            .PADIN(N__14971),
            .CLOCKENABLE(),
            .DIN0(write_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_data_ibuf_4_iopad (
            .OE(N__14964),
            .DIN(N__14963),
            .DOUT(N__14962),
            .PACKAGEPIN(write_data[4]));
    defparam write_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam write_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO write_data_ibuf_4_preio (
            .PADOEN(N__14964),
            .PADOUT(N__14963),
            .PADIN(N__14962),
            .CLOCKENABLE(),
            .DIN0(write_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_data_ibuf_5_iopad (
            .OE(N__14955),
            .DIN(N__14954),
            .DOUT(N__14953),
            .PACKAGEPIN(write_data[5]));
    defparam write_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam write_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO write_data_ibuf_5_preio (
            .PADOEN(N__14955),
            .PADOUT(N__14954),
            .PADIN(N__14953),
            .CLOCKENABLE(),
            .DIN0(write_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD write_en_ibuf_iopad (
            .OE(N__14946),
            .DIN(N__14945),
            .DOUT(N__14944),
            .PACKAGEPIN(write_en));
    defparam write_en_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam write_en_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO write_en_ibuf_preio (
            .PADOEN(N__14946),
            .PADOUT(N__14945),
            .PADIN(N__14944),
            .CLOCKENABLE(),
            .DIN0(write_en_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CEMux I__3638 (
            .O(N__14927),
            .I(N__14923));
    CEMux I__3637 (
            .O(N__14926),
            .I(N__14920));
    LocalMux I__3636 (
            .O(N__14923),
            .I(N__14914));
    LocalMux I__3635 (
            .O(N__14920),
            .I(N__14914));
    CEMux I__3634 (
            .O(N__14919),
            .I(N__14911));
    Span4Mux_v I__3633 (
            .O(N__14914),
            .I(N__14906));
    LocalMux I__3632 (
            .O(N__14911),
            .I(N__14906));
    Span4Mux_v I__3631 (
            .O(N__14906),
            .I(N__14903));
    Odrv4 I__3630 (
            .O(N__14903),
            .I(\this_vram.mem_WE_0 ));
    InMux I__3629 (
            .O(N__14900),
            .I(N__14896));
    InMux I__3628 (
            .O(N__14899),
            .I(N__14892));
    LocalMux I__3627 (
            .O(N__14896),
            .I(N__14889));
    InMux I__3626 (
            .O(N__14895),
            .I(N__14886));
    LocalMux I__3625 (
            .O(N__14892),
            .I(N__14882));
    Span4Mux_v I__3624 (
            .O(N__14889),
            .I(N__14877));
    LocalMux I__3623 (
            .O(N__14886),
            .I(N__14877));
    InMux I__3622 (
            .O(N__14885),
            .I(N__14874));
    Span4Mux_v I__3621 (
            .O(N__14882),
            .I(N__14871));
    Span4Mux_h I__3620 (
            .O(N__14877),
            .I(N__14865));
    LocalMux I__3619 (
            .O(N__14874),
            .I(N__14865));
    Span4Mux_h I__3618 (
            .O(N__14871),
            .I(N__14861));
    InMux I__3617 (
            .O(N__14870),
            .I(N__14858));
    Span4Mux_v I__3616 (
            .O(N__14865),
            .I(N__14855));
    InMux I__3615 (
            .O(N__14864),
            .I(N__14852));
    Span4Mux_h I__3614 (
            .O(N__14861),
            .I(N__14847));
    LocalMux I__3613 (
            .O(N__14858),
            .I(N__14847));
    Sp12to4 I__3612 (
            .O(N__14855),
            .I(N__14839));
    LocalMux I__3611 (
            .O(N__14852),
            .I(N__14839));
    Span4Mux_v I__3610 (
            .O(N__14847),
            .I(N__14836));
    InMux I__3609 (
            .O(N__14846),
            .I(N__14831));
    InMux I__3608 (
            .O(N__14845),
            .I(N__14831));
    InMux I__3607 (
            .O(N__14844),
            .I(N__14828));
    Span12Mux_h I__3606 (
            .O(N__14839),
            .I(N__14825));
    Span4Mux_h I__3605 (
            .O(N__14836),
            .I(N__14822));
    LocalMux I__3604 (
            .O(N__14831),
            .I(N__14817));
    LocalMux I__3603 (
            .O(N__14828),
            .I(N__14817));
    Span12Mux_h I__3602 (
            .O(N__14825),
            .I(N__14814));
    Sp12to4 I__3601 (
            .O(N__14822),
            .I(N__14809));
    Span12Mux_v I__3600 (
            .O(N__14817),
            .I(N__14809));
    Odrv12 I__3599 (
            .O(N__14814),
            .I(write_address_c_13));
    Odrv12 I__3598 (
            .O(N__14809),
            .I(write_address_c_13));
    InMux I__3597 (
            .O(N__14804),
            .I(N__14797));
    InMux I__3596 (
            .O(N__14803),
            .I(N__14794));
    InMux I__3595 (
            .O(N__14802),
            .I(N__14790));
    InMux I__3594 (
            .O(N__14801),
            .I(N__14785));
    InMux I__3593 (
            .O(N__14800),
            .I(N__14785));
    LocalMux I__3592 (
            .O(N__14797),
            .I(N__14781));
    LocalMux I__3591 (
            .O(N__14794),
            .I(N__14778));
    InMux I__3590 (
            .O(N__14793),
            .I(N__14775));
    LocalMux I__3589 (
            .O(N__14790),
            .I(N__14771));
    LocalMux I__3588 (
            .O(N__14785),
            .I(N__14768));
    InMux I__3587 (
            .O(N__14784),
            .I(N__14764));
    Span4Mux_v I__3586 (
            .O(N__14781),
            .I(N__14757));
    Span4Mux_h I__3585 (
            .O(N__14778),
            .I(N__14757));
    LocalMux I__3584 (
            .O(N__14775),
            .I(N__14757));
    InMux I__3583 (
            .O(N__14774),
            .I(N__14754));
    Span4Mux_v I__3582 (
            .O(N__14771),
            .I(N__14751));
    Span4Mux_h I__3581 (
            .O(N__14768),
            .I(N__14748));
    InMux I__3580 (
            .O(N__14767),
            .I(N__14745));
    LocalMux I__3579 (
            .O(N__14764),
            .I(N__14738));
    Sp12to4 I__3578 (
            .O(N__14757),
            .I(N__14738));
    LocalMux I__3577 (
            .O(N__14754),
            .I(N__14738));
    Span4Mux_v I__3576 (
            .O(N__14751),
            .I(N__14735));
    Span4Mux_v I__3575 (
            .O(N__14748),
            .I(N__14730));
    LocalMux I__3574 (
            .O(N__14745),
            .I(N__14730));
    Span12Mux_v I__3573 (
            .O(N__14738),
            .I(N__14727));
    Sp12to4 I__3572 (
            .O(N__14735),
            .I(N__14724));
    Span4Mux_v I__3571 (
            .O(N__14730),
            .I(N__14721));
    Span12Mux_h I__3570 (
            .O(N__14727),
            .I(N__14718));
    Span12Mux_h I__3569 (
            .O(N__14724),
            .I(N__14715));
    Span4Mux_h I__3568 (
            .O(N__14721),
            .I(N__14712));
    Odrv12 I__3567 (
            .O(N__14718),
            .I(write_address_c_12));
    Odrv12 I__3566 (
            .O(N__14715),
            .I(write_address_c_12));
    Odrv4 I__3565 (
            .O(N__14712),
            .I(write_address_c_12));
    InMux I__3564 (
            .O(N__14705),
            .I(N__14702));
    LocalMux I__3563 (
            .O(N__14702),
            .I(\this_vram.mem_N_29 ));
    InMux I__3562 (
            .O(N__14699),
            .I(N__14690));
    InMux I__3561 (
            .O(N__14698),
            .I(N__14690));
    InMux I__3560 (
            .O(N__14697),
            .I(N__14690));
    LocalMux I__3559 (
            .O(N__14690),
            .I(N__14687));
    Span12Mux_v I__3558 (
            .O(N__14687),
            .I(N__14684));
    Odrv12 I__3557 (
            .O(N__14684),
            .I(write_address_c_14));
    CascadeMux I__3556 (
            .O(N__14681),
            .I(N__14677));
    InMux I__3555 (
            .O(N__14680),
            .I(N__14672));
    InMux I__3554 (
            .O(N__14677),
            .I(N__14669));
    InMux I__3553 (
            .O(N__14676),
            .I(N__14666));
    InMux I__3552 (
            .O(N__14675),
            .I(N__14663));
    LocalMux I__3551 (
            .O(N__14672),
            .I(N__14660));
    LocalMux I__3550 (
            .O(N__14669),
            .I(N__14656));
    LocalMux I__3549 (
            .O(N__14666),
            .I(N__14651));
    LocalMux I__3548 (
            .O(N__14663),
            .I(N__14651));
    Span4Mux_v I__3547 (
            .O(N__14660),
            .I(N__14647));
    InMux I__3546 (
            .O(N__14659),
            .I(N__14644));
    Span4Mux_v I__3545 (
            .O(N__14656),
            .I(N__14639));
    Span4Mux_v I__3544 (
            .O(N__14651),
            .I(N__14639));
    InMux I__3543 (
            .O(N__14650),
            .I(N__14636));
    Span4Mux_v I__3542 (
            .O(N__14647),
            .I(N__14631));
    LocalMux I__3541 (
            .O(N__14644),
            .I(N__14631));
    Sp12to4 I__3540 (
            .O(N__14639),
            .I(N__14626));
    LocalMux I__3539 (
            .O(N__14636),
            .I(N__14623));
    Span4Mux_v I__3538 (
            .O(N__14631),
            .I(N__14620));
    InMux I__3537 (
            .O(N__14630),
            .I(N__14615));
    InMux I__3536 (
            .O(N__14629),
            .I(N__14615));
    Span12Mux_h I__3535 (
            .O(N__14626),
            .I(N__14608));
    Sp12to4 I__3534 (
            .O(N__14623),
            .I(N__14608));
    Span4Mux_v I__3533 (
            .O(N__14620),
            .I(N__14605));
    LocalMux I__3532 (
            .O(N__14615),
            .I(N__14602));
    InMux I__3531 (
            .O(N__14614),
            .I(N__14597));
    InMux I__3530 (
            .O(N__14613),
            .I(N__14597));
    Span12Mux_v I__3529 (
            .O(N__14608),
            .I(N__14594));
    Sp12to4 I__3528 (
            .O(N__14605),
            .I(N__14591));
    Sp12to4 I__3527 (
            .O(N__14602),
            .I(N__14586));
    LocalMux I__3526 (
            .O(N__14597),
            .I(N__14586));
    Span12Mux_h I__3525 (
            .O(N__14594),
            .I(N__14583));
    Span12Mux_h I__3524 (
            .O(N__14591),
            .I(N__14578));
    Span12Mux_v I__3523 (
            .O(N__14586),
            .I(N__14578));
    Odrv12 I__3522 (
            .O(N__14583),
            .I(write_address_c_11));
    Odrv12 I__3521 (
            .O(N__14578),
            .I(write_address_c_11));
    CascadeMux I__3520 (
            .O(N__14573),
            .I(\this_vram.mem_N_29_cascade_ ));
    CascadeMux I__3519 (
            .O(N__14570),
            .I(N__14567));
    InMux I__3518 (
            .O(N__14567),
            .I(N__14562));
    InMux I__3517 (
            .O(N__14566),
            .I(N__14557));
    InMux I__3516 (
            .O(N__14565),
            .I(N__14557));
    LocalMux I__3515 (
            .O(N__14562),
            .I(N__14552));
    LocalMux I__3514 (
            .O(N__14557),
            .I(N__14552));
    Span12Mux_v I__3513 (
            .O(N__14552),
            .I(N__14549));
    Span12Mux_h I__3512 (
            .O(N__14549),
            .I(N__14546));
    Odrv12 I__3511 (
            .O(N__14546),
            .I(write_en_c));
    CEMux I__3510 (
            .O(N__14543),
            .I(N__14539));
    CEMux I__3509 (
            .O(N__14542),
            .I(N__14536));
    LocalMux I__3508 (
            .O(N__14539),
            .I(N__14532));
    LocalMux I__3507 (
            .O(N__14536),
            .I(N__14529));
    CEMux I__3506 (
            .O(N__14535),
            .I(N__14526));
    Span4Mux_h I__3505 (
            .O(N__14532),
            .I(N__14521));
    Span4Mux_h I__3504 (
            .O(N__14529),
            .I(N__14521));
    LocalMux I__3503 (
            .O(N__14526),
            .I(N__14518));
    Odrv4 I__3502 (
            .O(N__14521),
            .I(\this_vram.mem_WE_3 ));
    Odrv4 I__3501 (
            .O(N__14518),
            .I(\this_vram.mem_WE_3 ));
    InMux I__3500 (
            .O(N__14513),
            .I(N__14510));
    LocalMux I__3499 (
            .O(N__14510),
            .I(N__14507));
    Span4Mux_v I__3498 (
            .O(N__14507),
            .I(N__14504));
    Odrv4 I__3497 (
            .O(N__14504),
            .I(\this_vram.mem_out_bus9_3 ));
    InMux I__3496 (
            .O(N__14501),
            .I(N__14498));
    LocalMux I__3495 (
            .O(N__14498),
            .I(N__14495));
    Odrv4 I__3494 (
            .O(N__14495),
            .I(\this_vram.mem_out_bus8_3 ));
    InMux I__3493 (
            .O(N__14492),
            .I(N__14489));
    LocalMux I__3492 (
            .O(N__14489),
            .I(N__14486));
    Span12Mux_h I__3491 (
            .O(N__14486),
            .I(N__14483));
    Odrv12 I__3490 (
            .O(N__14483),
            .I(\this_vram.mem_mem_8_1_RNI7H021Z0Z_0 ));
    InMux I__3489 (
            .O(N__14480),
            .I(N__14471));
    InMux I__3488 (
            .O(N__14479),
            .I(N__14471));
    InMux I__3487 (
            .O(N__14478),
            .I(N__14468));
    InMux I__3486 (
            .O(N__14477),
            .I(N__14457));
    InMux I__3485 (
            .O(N__14476),
            .I(N__14457));
    LocalMux I__3484 (
            .O(N__14471),
            .I(N__14449));
    LocalMux I__3483 (
            .O(N__14468),
            .I(N__14446));
    InMux I__3482 (
            .O(N__14467),
            .I(N__14443));
    InMux I__3481 (
            .O(N__14466),
            .I(N__14440));
    InMux I__3480 (
            .O(N__14465),
            .I(N__14437));
    InMux I__3479 (
            .O(N__14464),
            .I(N__14432));
    InMux I__3478 (
            .O(N__14463),
            .I(N__14426));
    InMux I__3477 (
            .O(N__14462),
            .I(N__14426));
    LocalMux I__3476 (
            .O(N__14457),
            .I(N__14422));
    InMux I__3475 (
            .O(N__14456),
            .I(N__14419));
    InMux I__3474 (
            .O(N__14455),
            .I(N__14416));
    InMux I__3473 (
            .O(N__14454),
            .I(N__14413));
    InMux I__3472 (
            .O(N__14453),
            .I(N__14408));
    InMux I__3471 (
            .O(N__14452),
            .I(N__14408));
    Span4Mux_v I__3470 (
            .O(N__14449),
            .I(N__14395));
    Span4Mux_v I__3469 (
            .O(N__14446),
            .I(N__14395));
    LocalMux I__3468 (
            .O(N__14443),
            .I(N__14395));
    LocalMux I__3467 (
            .O(N__14440),
            .I(N__14395));
    LocalMux I__3466 (
            .O(N__14437),
            .I(N__14395));
    InMux I__3465 (
            .O(N__14436),
            .I(N__14392));
    InMux I__3464 (
            .O(N__14435),
            .I(N__14389));
    LocalMux I__3463 (
            .O(N__14432),
            .I(N__14386));
    InMux I__3462 (
            .O(N__14431),
            .I(N__14383));
    LocalMux I__3461 (
            .O(N__14426),
            .I(N__14380));
    InMux I__3460 (
            .O(N__14425),
            .I(N__14377));
    Span4Mux_v I__3459 (
            .O(N__14422),
            .I(N__14372));
    LocalMux I__3458 (
            .O(N__14419),
            .I(N__14372));
    LocalMux I__3457 (
            .O(N__14416),
            .I(N__14365));
    LocalMux I__3456 (
            .O(N__14413),
            .I(N__14365));
    LocalMux I__3455 (
            .O(N__14408),
            .I(N__14365));
    InMux I__3454 (
            .O(N__14407),
            .I(N__14362));
    InMux I__3453 (
            .O(N__14406),
            .I(N__14358));
    Span4Mux_v I__3452 (
            .O(N__14395),
            .I(N__14354));
    LocalMux I__3451 (
            .O(N__14392),
            .I(N__14349));
    LocalMux I__3450 (
            .O(N__14389),
            .I(N__14349));
    Span4Mux_v I__3449 (
            .O(N__14386),
            .I(N__14344));
    LocalMux I__3448 (
            .O(N__14383),
            .I(N__14344));
    Span4Mux_h I__3447 (
            .O(N__14380),
            .I(N__14339));
    LocalMux I__3446 (
            .O(N__14377),
            .I(N__14339));
    Span4Mux_v I__3445 (
            .O(N__14372),
            .I(N__14334));
    Span4Mux_v I__3444 (
            .O(N__14365),
            .I(N__14334));
    LocalMux I__3443 (
            .O(N__14362),
            .I(N__14331));
    InMux I__3442 (
            .O(N__14361),
            .I(N__14328));
    LocalMux I__3441 (
            .O(N__14358),
            .I(N__14325));
    InMux I__3440 (
            .O(N__14357),
            .I(N__14322));
    Sp12to4 I__3439 (
            .O(N__14354),
            .I(N__14319));
    Span12Mux_h I__3438 (
            .O(N__14349),
            .I(N__14316));
    Span4Mux_v I__3437 (
            .O(N__14344),
            .I(N__14311));
    Span4Mux_v I__3436 (
            .O(N__14339),
            .I(N__14311));
    Span4Mux_h I__3435 (
            .O(N__14334),
            .I(N__14306));
    Span4Mux_v I__3434 (
            .O(N__14331),
            .I(N__14306));
    LocalMux I__3433 (
            .O(N__14328),
            .I(N__14299));
    Span12Mux_v I__3432 (
            .O(N__14325),
            .I(N__14299));
    LocalMux I__3431 (
            .O(N__14322),
            .I(N__14299));
    Odrv12 I__3430 (
            .O(N__14319),
            .I(\this_vram.mem_radregZ0Z_11 ));
    Odrv12 I__3429 (
            .O(N__14316),
            .I(\this_vram.mem_radregZ0Z_11 ));
    Odrv4 I__3428 (
            .O(N__14311),
            .I(\this_vram.mem_radregZ0Z_11 ));
    Odrv4 I__3427 (
            .O(N__14306),
            .I(\this_vram.mem_radregZ0Z_11 ));
    Odrv12 I__3426 (
            .O(N__14299),
            .I(\this_vram.mem_radregZ0Z_11 ));
    CascadeMux I__3425 (
            .O(N__14288),
            .I(N__14285));
    InMux I__3424 (
            .O(N__14285),
            .I(N__14282));
    LocalMux I__3423 (
            .O(N__14282),
            .I(\this_vram.mem_out_bus8_4 ));
    InMux I__3422 (
            .O(N__14279),
            .I(N__14276));
    LocalMux I__3421 (
            .O(N__14276),
            .I(N__14273));
    Sp12to4 I__3420 (
            .O(N__14273),
            .I(N__14270));
    Odrv12 I__3419 (
            .O(N__14270),
            .I(\this_vram.mem_out_bus9_4 ));
    InMux I__3418 (
            .O(N__14267),
            .I(N__14264));
    LocalMux I__3417 (
            .O(N__14264),
            .I(N__14261));
    Span12Mux_h I__3416 (
            .O(N__14261),
            .I(N__14258));
    Odrv12 I__3415 (
            .O(N__14258),
            .I(\this_vram.mem_mem_8_2_RNI9HZ0Z021 ));
    CEMux I__3414 (
            .O(N__14255),
            .I(N__14251));
    CEMux I__3413 (
            .O(N__14254),
            .I(N__14248));
    LocalMux I__3412 (
            .O(N__14251),
            .I(N__14242));
    LocalMux I__3411 (
            .O(N__14248),
            .I(N__14242));
    CEMux I__3410 (
            .O(N__14247),
            .I(N__14239));
    Span4Mux_v I__3409 (
            .O(N__14242),
            .I(N__14234));
    LocalMux I__3408 (
            .O(N__14239),
            .I(N__14234));
    Span4Mux_v I__3407 (
            .O(N__14234),
            .I(N__14231));
    Span4Mux_h I__3406 (
            .O(N__14231),
            .I(N__14228));
    Odrv4 I__3405 (
            .O(N__14228),
            .I(\this_vram.mem_WE_9 ));
    InMux I__3404 (
            .O(N__14225),
            .I(N__14222));
    LocalMux I__3403 (
            .O(N__14222),
            .I(N__14219));
    Odrv4 I__3402 (
            .O(N__14219),
            .I(\this_vram.mem_out_bus7_4 ));
    InMux I__3401 (
            .O(N__14216),
            .I(N__14213));
    LocalMux I__3400 (
            .O(N__14213),
            .I(N__14210));
    Span4Mux_v I__3399 (
            .O(N__14210),
            .I(N__14207));
    Span4Mux_v I__3398 (
            .O(N__14207),
            .I(N__14204));
    Odrv4 I__3397 (
            .O(N__14204),
            .I(\this_vram.mem_out_bus5_4 ));
    InMux I__3396 (
            .O(N__14201),
            .I(N__14198));
    LocalMux I__3395 (
            .O(N__14198),
            .I(N__14195));
    Span4Mux_v I__3394 (
            .O(N__14195),
            .I(N__14192));
    Sp12to4 I__3393 (
            .O(N__14192),
            .I(N__14189));
    Span12Mux_h I__3392 (
            .O(N__14189),
            .I(N__14186));
    Odrv12 I__3391 (
            .O(N__14186),
            .I(\this_vram.mem_mem_5_2_RNI58RZ0Z11 ));
    InMux I__3390 (
            .O(N__14183),
            .I(N__14180));
    LocalMux I__3389 (
            .O(N__14180),
            .I(\this_vram.mem_out_bus7_5 ));
    InMux I__3388 (
            .O(N__14177),
            .I(N__14165));
    InMux I__3387 (
            .O(N__14176),
            .I(N__14162));
    InMux I__3386 (
            .O(N__14175),
            .I(N__14158));
    InMux I__3385 (
            .O(N__14174),
            .I(N__14153));
    InMux I__3384 (
            .O(N__14173),
            .I(N__14150));
    InMux I__3383 (
            .O(N__14172),
            .I(N__14145));
    InMux I__3382 (
            .O(N__14171),
            .I(N__14145));
    InMux I__3381 (
            .O(N__14170),
            .I(N__14142));
    InMux I__3380 (
            .O(N__14169),
            .I(N__14134));
    InMux I__3379 (
            .O(N__14168),
            .I(N__14134));
    LocalMux I__3378 (
            .O(N__14165),
            .I(N__14129));
    LocalMux I__3377 (
            .O(N__14162),
            .I(N__14129));
    InMux I__3376 (
            .O(N__14161),
            .I(N__14126));
    LocalMux I__3375 (
            .O(N__14158),
            .I(N__14123));
    InMux I__3374 (
            .O(N__14157),
            .I(N__14120));
    InMux I__3373 (
            .O(N__14156),
            .I(N__14117));
    LocalMux I__3372 (
            .O(N__14153),
            .I(N__14110));
    LocalMux I__3371 (
            .O(N__14150),
            .I(N__14110));
    LocalMux I__3370 (
            .O(N__14145),
            .I(N__14110));
    LocalMux I__3369 (
            .O(N__14142),
            .I(N__14107));
    InMux I__3368 (
            .O(N__14141),
            .I(N__14104));
    InMux I__3367 (
            .O(N__14140),
            .I(N__14101));
    InMux I__3366 (
            .O(N__14139),
            .I(N__14098));
    LocalMux I__3365 (
            .O(N__14134),
            .I(N__14092));
    Span4Mux_v I__3364 (
            .O(N__14129),
            .I(N__14087));
    LocalMux I__3363 (
            .O(N__14126),
            .I(N__14087));
    Span4Mux_h I__3362 (
            .O(N__14123),
            .I(N__14082));
    LocalMux I__3361 (
            .O(N__14120),
            .I(N__14082));
    LocalMux I__3360 (
            .O(N__14117),
            .I(N__14079));
    Span4Mux_v I__3359 (
            .O(N__14110),
            .I(N__14076));
    Span4Mux_h I__3358 (
            .O(N__14107),
            .I(N__14071));
    LocalMux I__3357 (
            .O(N__14104),
            .I(N__14071));
    LocalMux I__3356 (
            .O(N__14101),
            .I(N__14066));
    LocalMux I__3355 (
            .O(N__14098),
            .I(N__14066));
    InMux I__3354 (
            .O(N__14097),
            .I(N__14063));
    InMux I__3353 (
            .O(N__14096),
            .I(N__14058));
    InMux I__3352 (
            .O(N__14095),
            .I(N__14058));
    Span12Mux_v I__3351 (
            .O(N__14092),
            .I(N__14055));
    Span4Mux_h I__3350 (
            .O(N__14087),
            .I(N__14050));
    Span4Mux_h I__3349 (
            .O(N__14082),
            .I(N__14050));
    Span4Mux_v I__3348 (
            .O(N__14079),
            .I(N__14047));
    Span4Mux_h I__3347 (
            .O(N__14076),
            .I(N__14042));
    Span4Mux_v I__3346 (
            .O(N__14071),
            .I(N__14042));
    Span12Mux_h I__3345 (
            .O(N__14066),
            .I(N__14035));
    LocalMux I__3344 (
            .O(N__14063),
            .I(N__14035));
    LocalMux I__3343 (
            .O(N__14058),
            .I(N__14035));
    Odrv12 I__3342 (
            .O(N__14055),
            .I(\this_vram.mem_radregZ0Z_12 ));
    Odrv4 I__3341 (
            .O(N__14050),
            .I(\this_vram.mem_radregZ0Z_12 ));
    Odrv4 I__3340 (
            .O(N__14047),
            .I(\this_vram.mem_radregZ0Z_12 ));
    Odrv4 I__3339 (
            .O(N__14042),
            .I(\this_vram.mem_radregZ0Z_12 ));
    Odrv12 I__3338 (
            .O(N__14035),
            .I(\this_vram.mem_radregZ0Z_12 ));
    InMux I__3337 (
            .O(N__14024),
            .I(N__14021));
    LocalMux I__3336 (
            .O(N__14021),
            .I(N__14018));
    Sp12to4 I__3335 (
            .O(N__14018),
            .I(N__14015));
    Span12Mux_v I__3334 (
            .O(N__14015),
            .I(N__14012));
    Odrv12 I__3333 (
            .O(N__14012),
            .I(\this_vram.mem_out_bus5_5 ));
    InMux I__3332 (
            .O(N__14009),
            .I(N__14006));
    LocalMux I__3331 (
            .O(N__14006),
            .I(N__14003));
    Span4Mux_v I__3330 (
            .O(N__14003),
            .I(N__14000));
    Span4Mux_h I__3329 (
            .O(N__14000),
            .I(N__13997));
    Odrv4 I__3328 (
            .O(N__13997),
            .I(\this_vram.mem_mem_5_2_RNI58R11Z0Z_0 ));
    CEMux I__3327 (
            .O(N__13994),
            .I(N__13989));
    CEMux I__3326 (
            .O(N__13993),
            .I(N__13986));
    CEMux I__3325 (
            .O(N__13992),
            .I(N__13983));
    LocalMux I__3324 (
            .O(N__13989),
            .I(N__13978));
    LocalMux I__3323 (
            .O(N__13986),
            .I(N__13978));
    LocalMux I__3322 (
            .O(N__13983),
            .I(N__13975));
    Span4Mux_v I__3321 (
            .O(N__13978),
            .I(N__13972));
    Span4Mux_h I__3320 (
            .O(N__13975),
            .I(N__13969));
    Odrv4 I__3319 (
            .O(N__13972),
            .I(\this_vram.mem_WE_6 ));
    Odrv4 I__3318 (
            .O(N__13969),
            .I(\this_vram.mem_WE_6 ));
    InMux I__3317 (
            .O(N__13964),
            .I(N__13961));
    LocalMux I__3316 (
            .O(N__13961),
            .I(N__13958));
    Span4Mux_v I__3315 (
            .O(N__13958),
            .I(N__13955));
    Odrv4 I__3314 (
            .O(N__13955),
            .I(\this_vram.mem_out_bus9_0 ));
    InMux I__3313 (
            .O(N__13952),
            .I(N__13949));
    LocalMux I__3312 (
            .O(N__13949),
            .I(\this_vram.mem_out_bus8_0 ));
    InMux I__3311 (
            .O(N__13946),
            .I(N__13943));
    LocalMux I__3310 (
            .O(N__13943),
            .I(N__13940));
    Span12Mux_v I__3309 (
            .O(N__13940),
            .I(N__13937));
    Span12Mux_h I__3308 (
            .O(N__13937),
            .I(N__13934));
    Odrv12 I__3307 (
            .O(N__13934),
            .I(\this_vram.mem_mem_8_0_RNI5HZ0Z021 ));
    InMux I__3306 (
            .O(N__13931),
            .I(N__13928));
    LocalMux I__3305 (
            .O(N__13928),
            .I(\this_vram.mem_out_bus8_1 ));
    InMux I__3304 (
            .O(N__13925),
            .I(N__13922));
    LocalMux I__3303 (
            .O(N__13922),
            .I(N__13919));
    Span4Mux_v I__3302 (
            .O(N__13919),
            .I(N__13916));
    Odrv4 I__3301 (
            .O(N__13916),
            .I(\this_vram.mem_out_bus9_1 ));
    InMux I__3300 (
            .O(N__13913),
            .I(N__13910));
    LocalMux I__3299 (
            .O(N__13910),
            .I(N__13907));
    Sp12to4 I__3298 (
            .O(N__13907),
            .I(N__13904));
    Span12Mux_h I__3297 (
            .O(N__13904),
            .I(N__13901));
    Odrv12 I__3296 (
            .O(N__13901),
            .I(\this_vram.mem_mem_8_0_RNI5H021Z0Z_0 ));
    InMux I__3295 (
            .O(N__13898),
            .I(N__13895));
    LocalMux I__3294 (
            .O(N__13895),
            .I(\this_vram.mem_out_bus8_2 ));
    InMux I__3293 (
            .O(N__13892),
            .I(N__13889));
    LocalMux I__3292 (
            .O(N__13889),
            .I(N__13886));
    Span4Mux_v I__3291 (
            .O(N__13886),
            .I(N__13883));
    Odrv4 I__3290 (
            .O(N__13883),
            .I(\this_vram.mem_out_bus9_2 ));
    InMux I__3289 (
            .O(N__13880),
            .I(N__13877));
    LocalMux I__3288 (
            .O(N__13877),
            .I(N__13874));
    Span12Mux_v I__3287 (
            .O(N__13874),
            .I(N__13871));
    Span12Mux_h I__3286 (
            .O(N__13871),
            .I(N__13868));
    Odrv12 I__3285 (
            .O(N__13868),
            .I(\this_vram.mem_mem_8_1_RNI7HZ0Z021 ));
    CascadeMux I__3284 (
            .O(N__13865),
            .I(N__13861));
    InMux I__3283 (
            .O(N__13864),
            .I(N__13855));
    InMux I__3282 (
            .O(N__13861),
            .I(N__13852));
    CascadeMux I__3281 (
            .O(N__13860),
            .I(N__13849));
    CascadeMux I__3280 (
            .O(N__13859),
            .I(N__13846));
    CascadeMux I__3279 (
            .O(N__13858),
            .I(N__13843));
    LocalMux I__3278 (
            .O(N__13855),
            .I(N__13838));
    LocalMux I__3277 (
            .O(N__13852),
            .I(N__13838));
    InMux I__3276 (
            .O(N__13849),
            .I(N__13835));
    InMux I__3275 (
            .O(N__13846),
            .I(N__13832));
    InMux I__3274 (
            .O(N__13843),
            .I(N__13829));
    Span4Mux_v I__3273 (
            .O(N__13838),
            .I(N__13821));
    LocalMux I__3272 (
            .O(N__13835),
            .I(N__13821));
    LocalMux I__3271 (
            .O(N__13832),
            .I(N__13821));
    LocalMux I__3270 (
            .O(N__13829),
            .I(N__13818));
    CascadeMux I__3269 (
            .O(N__13828),
            .I(N__13815));
    Span4Mux_v I__3268 (
            .O(N__13821),
            .I(N__13812));
    Span4Mux_v I__3267 (
            .O(N__13818),
            .I(N__13809));
    InMux I__3266 (
            .O(N__13815),
            .I(N__13806));
    Span4Mux_h I__3265 (
            .O(N__13812),
            .I(N__13801));
    Span4Mux_h I__3264 (
            .O(N__13809),
            .I(N__13798));
    LocalMux I__3263 (
            .O(N__13806),
            .I(N__13795));
    CascadeMux I__3262 (
            .O(N__13805),
            .I(N__13792));
    CascadeMux I__3261 (
            .O(N__13804),
            .I(N__13789));
    Span4Mux_h I__3260 (
            .O(N__13801),
            .I(N__13786));
    Span4Mux_h I__3259 (
            .O(N__13798),
            .I(N__13781));
    Span4Mux_v I__3258 (
            .O(N__13795),
            .I(N__13781));
    InMux I__3257 (
            .O(N__13792),
            .I(N__13776));
    InMux I__3256 (
            .O(N__13789),
            .I(N__13776));
    Span4Mux_h I__3255 (
            .O(N__13786),
            .I(N__13773));
    Span4Mux_h I__3254 (
            .O(N__13781),
            .I(N__13770));
    LocalMux I__3253 (
            .O(N__13776),
            .I(N__13767));
    Odrv4 I__3252 (
            .O(N__13773),
            .I(\this_vram.mem_N_27 ));
    Odrv4 I__3251 (
            .O(N__13770),
            .I(\this_vram.mem_N_27 ));
    Odrv12 I__3250 (
            .O(N__13767),
            .I(\this_vram.mem_N_27 ));
    InMux I__3249 (
            .O(N__13760),
            .I(N__13748));
    InMux I__3248 (
            .O(N__13759),
            .I(N__13748));
    InMux I__3247 (
            .O(N__13758),
            .I(N__13748));
    InMux I__3246 (
            .O(N__13757),
            .I(N__13748));
    LocalMux I__3245 (
            .O(N__13748),
            .I(N__13745));
    Span4Mux_v I__3244 (
            .O(N__13745),
            .I(N__13742));
    Span4Mux_v I__3243 (
            .O(N__13742),
            .I(N__13739));
    Sp12to4 I__3242 (
            .O(N__13739),
            .I(N__13736));
    Odrv12 I__3241 (
            .O(N__13736),
            .I(rst_n_c));
    InMux I__3240 (
            .O(N__13733),
            .I(N__13730));
    LocalMux I__3239 (
            .O(N__13730),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    ClkMux I__3238 (
            .O(N__13727),
            .I(N__13508));
    ClkMux I__3237 (
            .O(N__13726),
            .I(N__13508));
    ClkMux I__3236 (
            .O(N__13725),
            .I(N__13508));
    ClkMux I__3235 (
            .O(N__13724),
            .I(N__13508));
    ClkMux I__3234 (
            .O(N__13723),
            .I(N__13508));
    ClkMux I__3233 (
            .O(N__13722),
            .I(N__13508));
    ClkMux I__3232 (
            .O(N__13721),
            .I(N__13508));
    ClkMux I__3231 (
            .O(N__13720),
            .I(N__13508));
    ClkMux I__3230 (
            .O(N__13719),
            .I(N__13508));
    ClkMux I__3229 (
            .O(N__13718),
            .I(N__13508));
    ClkMux I__3228 (
            .O(N__13717),
            .I(N__13508));
    ClkMux I__3227 (
            .O(N__13716),
            .I(N__13508));
    ClkMux I__3226 (
            .O(N__13715),
            .I(N__13508));
    ClkMux I__3225 (
            .O(N__13714),
            .I(N__13508));
    ClkMux I__3224 (
            .O(N__13713),
            .I(N__13508));
    ClkMux I__3223 (
            .O(N__13712),
            .I(N__13508));
    ClkMux I__3222 (
            .O(N__13711),
            .I(N__13508));
    ClkMux I__3221 (
            .O(N__13710),
            .I(N__13508));
    ClkMux I__3220 (
            .O(N__13709),
            .I(N__13508));
    ClkMux I__3219 (
            .O(N__13708),
            .I(N__13508));
    ClkMux I__3218 (
            .O(N__13707),
            .I(N__13508));
    ClkMux I__3217 (
            .O(N__13706),
            .I(N__13508));
    ClkMux I__3216 (
            .O(N__13705),
            .I(N__13508));
    ClkMux I__3215 (
            .O(N__13704),
            .I(N__13508));
    ClkMux I__3214 (
            .O(N__13703),
            .I(N__13508));
    ClkMux I__3213 (
            .O(N__13702),
            .I(N__13508));
    ClkMux I__3212 (
            .O(N__13701),
            .I(N__13508));
    ClkMux I__3211 (
            .O(N__13700),
            .I(N__13508));
    ClkMux I__3210 (
            .O(N__13699),
            .I(N__13508));
    ClkMux I__3209 (
            .O(N__13698),
            .I(N__13508));
    ClkMux I__3208 (
            .O(N__13697),
            .I(N__13508));
    ClkMux I__3207 (
            .O(N__13696),
            .I(N__13508));
    ClkMux I__3206 (
            .O(N__13695),
            .I(N__13508));
    ClkMux I__3205 (
            .O(N__13694),
            .I(N__13508));
    ClkMux I__3204 (
            .O(N__13693),
            .I(N__13508));
    ClkMux I__3203 (
            .O(N__13692),
            .I(N__13508));
    ClkMux I__3202 (
            .O(N__13691),
            .I(N__13508));
    ClkMux I__3201 (
            .O(N__13690),
            .I(N__13508));
    ClkMux I__3200 (
            .O(N__13689),
            .I(N__13508));
    ClkMux I__3199 (
            .O(N__13688),
            .I(N__13508));
    ClkMux I__3198 (
            .O(N__13687),
            .I(N__13508));
    ClkMux I__3197 (
            .O(N__13686),
            .I(N__13508));
    ClkMux I__3196 (
            .O(N__13685),
            .I(N__13508));
    ClkMux I__3195 (
            .O(N__13684),
            .I(N__13508));
    ClkMux I__3194 (
            .O(N__13683),
            .I(N__13508));
    ClkMux I__3193 (
            .O(N__13682),
            .I(N__13508));
    ClkMux I__3192 (
            .O(N__13681),
            .I(N__13508));
    ClkMux I__3191 (
            .O(N__13680),
            .I(N__13508));
    ClkMux I__3190 (
            .O(N__13679),
            .I(N__13508));
    ClkMux I__3189 (
            .O(N__13678),
            .I(N__13508));
    ClkMux I__3188 (
            .O(N__13677),
            .I(N__13508));
    ClkMux I__3187 (
            .O(N__13676),
            .I(N__13508));
    ClkMux I__3186 (
            .O(N__13675),
            .I(N__13508));
    ClkMux I__3185 (
            .O(N__13674),
            .I(N__13508));
    ClkMux I__3184 (
            .O(N__13673),
            .I(N__13508));
    ClkMux I__3183 (
            .O(N__13672),
            .I(N__13508));
    ClkMux I__3182 (
            .O(N__13671),
            .I(N__13508));
    ClkMux I__3181 (
            .O(N__13670),
            .I(N__13508));
    ClkMux I__3180 (
            .O(N__13669),
            .I(N__13508));
    ClkMux I__3179 (
            .O(N__13668),
            .I(N__13508));
    ClkMux I__3178 (
            .O(N__13667),
            .I(N__13508));
    ClkMux I__3177 (
            .O(N__13666),
            .I(N__13508));
    ClkMux I__3176 (
            .O(N__13665),
            .I(N__13508));
    ClkMux I__3175 (
            .O(N__13664),
            .I(N__13508));
    ClkMux I__3174 (
            .O(N__13663),
            .I(N__13508));
    ClkMux I__3173 (
            .O(N__13662),
            .I(N__13508));
    ClkMux I__3172 (
            .O(N__13661),
            .I(N__13508));
    ClkMux I__3171 (
            .O(N__13660),
            .I(N__13508));
    ClkMux I__3170 (
            .O(N__13659),
            .I(N__13508));
    ClkMux I__3169 (
            .O(N__13658),
            .I(N__13508));
    ClkMux I__3168 (
            .O(N__13657),
            .I(N__13508));
    ClkMux I__3167 (
            .O(N__13656),
            .I(N__13508));
    ClkMux I__3166 (
            .O(N__13655),
            .I(N__13508));
    GlobalMux I__3165 (
            .O(N__13508),
            .I(N__13505));
    gio2CtrlBuf I__3164 (
            .O(N__13505),
            .I(clk_c_g));
    InMux I__3163 (
            .O(N__13502),
            .I(N__13499));
    LocalMux I__3162 (
            .O(N__13499),
            .I(N__13496));
    Span12Mux_v I__3161 (
            .O(N__13496),
            .I(N__13493));
    Odrv12 I__3160 (
            .O(N__13493),
            .I(\this_vram.mem_out_bus6_5 ));
    InMux I__3159 (
            .O(N__13490),
            .I(N__13487));
    LocalMux I__3158 (
            .O(N__13487),
            .I(N__13484));
    Span4Mux_v I__3157 (
            .O(N__13484),
            .I(N__13481));
    Span4Mux_v I__3156 (
            .O(N__13481),
            .I(N__13478));
    Sp12to4 I__3155 (
            .O(N__13478),
            .I(N__13475));
    Span12Mux_h I__3154 (
            .O(N__13475),
            .I(N__13472));
    Odrv12 I__3153 (
            .O(N__13472),
            .I(\this_vram.mem_out_bus4_5 ));
    CascadeMux I__3152 (
            .O(N__13469),
            .I(\this_vram.mem_mem_4_2_RNI34P11Z0Z_0_cascade_ ));
    InMux I__3151 (
            .O(N__13466),
            .I(N__13463));
    LocalMux I__3150 (
            .O(N__13463),
            .I(N__13460));
    Span4Mux_v I__3149 (
            .O(N__13460),
            .I(N__13457));
    Sp12to4 I__3148 (
            .O(N__13457),
            .I(N__13454));
    Odrv12 I__3147 (
            .O(N__13454),
            .I(\this_vram.mem_N_2372 ));
    CEMux I__3146 (
            .O(N__13451),
            .I(N__13448));
    LocalMux I__3145 (
            .O(N__13448),
            .I(N__13443));
    CEMux I__3144 (
            .O(N__13447),
            .I(N__13440));
    CEMux I__3143 (
            .O(N__13446),
            .I(N__13437));
    Span4Mux_s1_v I__3142 (
            .O(N__13443),
            .I(N__13432));
    LocalMux I__3141 (
            .O(N__13440),
            .I(N__13432));
    LocalMux I__3140 (
            .O(N__13437),
            .I(N__13429));
    Span4Mux_v I__3139 (
            .O(N__13432),
            .I(N__13426));
    Span4Mux_s3_v I__3138 (
            .O(N__13429),
            .I(N__13423));
    Sp12to4 I__3137 (
            .O(N__13426),
            .I(N__13420));
    Sp12to4 I__3136 (
            .O(N__13423),
            .I(N__13417));
    Span12Mux_h I__3135 (
            .O(N__13420),
            .I(N__13414));
    Span12Mux_v I__3134 (
            .O(N__13417),
            .I(N__13411));
    Span12Mux_v I__3133 (
            .O(N__13414),
            .I(N__13408));
    Odrv12 I__3132 (
            .O(N__13411),
            .I(\this_vram.mem_WE_12 ));
    Odrv12 I__3131 (
            .O(N__13408),
            .I(\this_vram.mem_WE_12 ));
    SRMux I__3130 (
            .O(N__13403),
            .I(N__13397));
    SRMux I__3129 (
            .O(N__13402),
            .I(N__13393));
    SRMux I__3128 (
            .O(N__13401),
            .I(N__13390));
    SRMux I__3127 (
            .O(N__13400),
            .I(N__13387));
    LocalMux I__3126 (
            .O(N__13397),
            .I(N__13375));
    SRMux I__3125 (
            .O(N__13396),
            .I(N__13372));
    LocalMux I__3124 (
            .O(N__13393),
            .I(N__13367));
    LocalMux I__3123 (
            .O(N__13390),
            .I(N__13367));
    LocalMux I__3122 (
            .O(N__13387),
            .I(N__13364));
    SRMux I__3121 (
            .O(N__13386),
            .I(N__13361));
    SRMux I__3120 (
            .O(N__13385),
            .I(N__13358));
    SRMux I__3119 (
            .O(N__13384),
            .I(N__13355));
    SRMux I__3118 (
            .O(N__13383),
            .I(N__13349));
    SRMux I__3117 (
            .O(N__13382),
            .I(N__13344));
    SRMux I__3116 (
            .O(N__13381),
            .I(N__13341));
    SRMux I__3115 (
            .O(N__13380),
            .I(N__13336));
    SRMux I__3114 (
            .O(N__13379),
            .I(N__13333));
    SRMux I__3113 (
            .O(N__13378),
            .I(N__13329));
    Span4Mux_s3_v I__3112 (
            .O(N__13375),
            .I(N__13326));
    LocalMux I__3111 (
            .O(N__13372),
            .I(N__13323));
    Span4Mux_s3_v I__3110 (
            .O(N__13367),
            .I(N__13314));
    Span4Mux_h I__3109 (
            .O(N__13364),
            .I(N__13314));
    LocalMux I__3108 (
            .O(N__13361),
            .I(N__13314));
    LocalMux I__3107 (
            .O(N__13358),
            .I(N__13314));
    LocalMux I__3106 (
            .O(N__13355),
            .I(N__13311));
    SRMux I__3105 (
            .O(N__13354),
            .I(N__13308));
    SRMux I__3104 (
            .O(N__13353),
            .I(N__13305));
    SRMux I__3103 (
            .O(N__13352),
            .I(N__13302));
    LocalMux I__3102 (
            .O(N__13349),
            .I(N__13297));
    SRMux I__3101 (
            .O(N__13348),
            .I(N__13294));
    SRMux I__3100 (
            .O(N__13347),
            .I(N__13291));
    LocalMux I__3099 (
            .O(N__13344),
            .I(N__13286));
    LocalMux I__3098 (
            .O(N__13341),
            .I(N__13286));
    SRMux I__3097 (
            .O(N__13340),
            .I(N__13283));
    SRMux I__3096 (
            .O(N__13339),
            .I(N__13280));
    LocalMux I__3095 (
            .O(N__13336),
            .I(N__13273));
    LocalMux I__3094 (
            .O(N__13333),
            .I(N__13270));
    SRMux I__3093 (
            .O(N__13332),
            .I(N__13267));
    LocalMux I__3092 (
            .O(N__13329),
            .I(N__13262));
    Span4Mux_v I__3091 (
            .O(N__13326),
            .I(N__13249));
    Span4Mux_v I__3090 (
            .O(N__13323),
            .I(N__13249));
    Span4Mux_v I__3089 (
            .O(N__13314),
            .I(N__13249));
    Span4Mux_h I__3088 (
            .O(N__13311),
            .I(N__13249));
    LocalMux I__3087 (
            .O(N__13308),
            .I(N__13249));
    LocalMux I__3086 (
            .O(N__13305),
            .I(N__13249));
    LocalMux I__3085 (
            .O(N__13302),
            .I(N__13246));
    SRMux I__3084 (
            .O(N__13301),
            .I(N__13243));
    SRMux I__3083 (
            .O(N__13300),
            .I(N__13240));
    Span4Mux_v I__3082 (
            .O(N__13297),
            .I(N__13230));
    LocalMux I__3081 (
            .O(N__13294),
            .I(N__13230));
    LocalMux I__3080 (
            .O(N__13291),
            .I(N__13230));
    Span4Mux_v I__3079 (
            .O(N__13286),
            .I(N__13223));
    LocalMux I__3078 (
            .O(N__13283),
            .I(N__13223));
    LocalMux I__3077 (
            .O(N__13280),
            .I(N__13223));
    SRMux I__3076 (
            .O(N__13279),
            .I(N__13220));
    SRMux I__3075 (
            .O(N__13278),
            .I(N__13217));
    SRMux I__3074 (
            .O(N__13277),
            .I(N__13214));
    SRMux I__3073 (
            .O(N__13276),
            .I(N__13211));
    Span4Mux_v I__3072 (
            .O(N__13273),
            .I(N__13201));
    Span4Mux_h I__3071 (
            .O(N__13270),
            .I(N__13201));
    LocalMux I__3070 (
            .O(N__13267),
            .I(N__13201));
    SRMux I__3069 (
            .O(N__13266),
            .I(N__13198));
    SRMux I__3068 (
            .O(N__13265),
            .I(N__13195));
    Span4Mux_v I__3067 (
            .O(N__13262),
            .I(N__13183));
    Span4Mux_v I__3066 (
            .O(N__13249),
            .I(N__13183));
    Span4Mux_h I__3065 (
            .O(N__13246),
            .I(N__13183));
    LocalMux I__3064 (
            .O(N__13243),
            .I(N__13183));
    LocalMux I__3063 (
            .O(N__13240),
            .I(N__13183));
    SRMux I__3062 (
            .O(N__13239),
            .I(N__13180));
    SRMux I__3061 (
            .O(N__13238),
            .I(N__13177));
    SRMux I__3060 (
            .O(N__13237),
            .I(N__13174));
    Span4Mux_v I__3059 (
            .O(N__13230),
            .I(N__13162));
    Span4Mux_v I__3058 (
            .O(N__13223),
            .I(N__13162));
    LocalMux I__3057 (
            .O(N__13220),
            .I(N__13162));
    LocalMux I__3056 (
            .O(N__13217),
            .I(N__13162));
    LocalMux I__3055 (
            .O(N__13214),
            .I(N__13157));
    LocalMux I__3054 (
            .O(N__13211),
            .I(N__13157));
    SRMux I__3053 (
            .O(N__13210),
            .I(N__13154));
    SRMux I__3052 (
            .O(N__13209),
            .I(N__13151));
    SRMux I__3051 (
            .O(N__13208),
            .I(N__13143));
    Span4Mux_v I__3050 (
            .O(N__13201),
            .I(N__13138));
    LocalMux I__3049 (
            .O(N__13198),
            .I(N__13138));
    LocalMux I__3048 (
            .O(N__13195),
            .I(N__13135));
    SRMux I__3047 (
            .O(N__13194),
            .I(N__13132));
    Span4Mux_v I__3046 (
            .O(N__13183),
            .I(N__13124));
    LocalMux I__3045 (
            .O(N__13180),
            .I(N__13124));
    LocalMux I__3044 (
            .O(N__13177),
            .I(N__13124));
    LocalMux I__3043 (
            .O(N__13174),
            .I(N__13121));
    SRMux I__3042 (
            .O(N__13173),
            .I(N__13118));
    SRMux I__3041 (
            .O(N__13172),
            .I(N__13115));
    SRMux I__3040 (
            .O(N__13171),
            .I(N__13111));
    Span4Mux_v I__3039 (
            .O(N__13162),
            .I(N__13101));
    Span4Mux_v I__3038 (
            .O(N__13157),
            .I(N__13101));
    LocalMux I__3037 (
            .O(N__13154),
            .I(N__13101));
    LocalMux I__3036 (
            .O(N__13151),
            .I(N__13101));
    SRMux I__3035 (
            .O(N__13150),
            .I(N__13098));
    SRMux I__3034 (
            .O(N__13149),
            .I(N__13095));
    SRMux I__3033 (
            .O(N__13148),
            .I(N__13092));
    SRMux I__3032 (
            .O(N__13147),
            .I(N__13089));
    SRMux I__3031 (
            .O(N__13146),
            .I(N__13081));
    LocalMux I__3030 (
            .O(N__13143),
            .I(N__13078));
    Span4Mux_v I__3029 (
            .O(N__13138),
            .I(N__13071));
    Span4Mux_h I__3028 (
            .O(N__13135),
            .I(N__13071));
    LocalMux I__3027 (
            .O(N__13132),
            .I(N__13071));
    SRMux I__3026 (
            .O(N__13131),
            .I(N__13068));
    Span4Mux_v I__3025 (
            .O(N__13124),
            .I(N__13059));
    Span4Mux_h I__3024 (
            .O(N__13121),
            .I(N__13059));
    LocalMux I__3023 (
            .O(N__13118),
            .I(N__13059));
    LocalMux I__3022 (
            .O(N__13115),
            .I(N__13059));
    SRMux I__3021 (
            .O(N__13114),
            .I(N__13056));
    LocalMux I__3020 (
            .O(N__13111),
            .I(N__13053));
    SRMux I__3019 (
            .O(N__13110),
            .I(N__13050));
    Span4Mux_v I__3018 (
            .O(N__13101),
            .I(N__13042));
    LocalMux I__3017 (
            .O(N__13098),
            .I(N__13042));
    LocalMux I__3016 (
            .O(N__13095),
            .I(N__13042));
    LocalMux I__3015 (
            .O(N__13092),
            .I(N__13037));
    LocalMux I__3014 (
            .O(N__13089),
            .I(N__13037));
    SRMux I__3013 (
            .O(N__13088),
            .I(N__13034));
    SRMux I__3012 (
            .O(N__13087),
            .I(N__13031));
    CascadeMux I__3011 (
            .O(N__13086),
            .I(N__13026));
    CascadeMux I__3010 (
            .O(N__13085),
            .I(N__13022));
    CascadeMux I__3009 (
            .O(N__13084),
            .I(N__13018));
    LocalMux I__3008 (
            .O(N__13081),
            .I(N__13007));
    Span4Mux_h I__3007 (
            .O(N__13078),
            .I(N__13007));
    Span4Mux_v I__3006 (
            .O(N__13071),
            .I(N__13007));
    LocalMux I__3005 (
            .O(N__13068),
            .I(N__13007));
    Span4Mux_v I__3004 (
            .O(N__13059),
            .I(N__12998));
    LocalMux I__3003 (
            .O(N__13056),
            .I(N__12998));
    Span4Mux_v I__3002 (
            .O(N__13053),
            .I(N__12998));
    LocalMux I__3001 (
            .O(N__13050),
            .I(N__12998));
    SRMux I__3000 (
            .O(N__13049),
            .I(N__12994));
    Span4Mux_v I__2999 (
            .O(N__13042),
            .I(N__12990));
    Span4Mux_v I__2998 (
            .O(N__13037),
            .I(N__12983));
    LocalMux I__2997 (
            .O(N__13034),
            .I(N__12983));
    LocalMux I__2996 (
            .O(N__13031),
            .I(N__12983));
    SRMux I__2995 (
            .O(N__13030),
            .I(N__12980));
    InMux I__2994 (
            .O(N__13029),
            .I(N__12964));
    InMux I__2993 (
            .O(N__13026),
            .I(N__12964));
    InMux I__2992 (
            .O(N__13025),
            .I(N__12964));
    InMux I__2991 (
            .O(N__13022),
            .I(N__12964));
    InMux I__2990 (
            .O(N__13021),
            .I(N__12964));
    InMux I__2989 (
            .O(N__13018),
            .I(N__12964));
    InMux I__2988 (
            .O(N__13017),
            .I(N__12964));
    SRMux I__2987 (
            .O(N__13016),
            .I(N__12961));
    Span4Mux_v I__2986 (
            .O(N__13007),
            .I(N__12956));
    Span4Mux_v I__2985 (
            .O(N__12998),
            .I(N__12956));
    SRMux I__2984 (
            .O(N__12997),
            .I(N__12951));
    LocalMux I__2983 (
            .O(N__12994),
            .I(N__12948));
    SRMux I__2982 (
            .O(N__12993),
            .I(N__12945));
    Span4Mux_h I__2981 (
            .O(N__12990),
            .I(N__12938));
    Span4Mux_v I__2980 (
            .O(N__12983),
            .I(N__12938));
    LocalMux I__2979 (
            .O(N__12980),
            .I(N__12938));
    SRMux I__2978 (
            .O(N__12979),
            .I(N__12935));
    LocalMux I__2977 (
            .O(N__12964),
            .I(N__12931));
    LocalMux I__2976 (
            .O(N__12961),
            .I(N__12928));
    Span4Mux_h I__2975 (
            .O(N__12956),
            .I(N__12925));
    SRMux I__2974 (
            .O(N__12955),
            .I(N__12922));
    SRMux I__2973 (
            .O(N__12954),
            .I(N__12919));
    LocalMux I__2972 (
            .O(N__12951),
            .I(N__12912));
    Span4Mux_h I__2971 (
            .O(N__12948),
            .I(N__12912));
    LocalMux I__2970 (
            .O(N__12945),
            .I(N__12912));
    Span4Mux_v I__2969 (
            .O(N__12938),
            .I(N__12907));
    LocalMux I__2968 (
            .O(N__12935),
            .I(N__12907));
    SRMux I__2967 (
            .O(N__12934),
            .I(N__12904));
    Span4Mux_v I__2966 (
            .O(N__12931),
            .I(N__12901));
    Span4Mux_h I__2965 (
            .O(N__12928),
            .I(N__12898));
    Span4Mux_h I__2964 (
            .O(N__12925),
            .I(N__12894));
    LocalMux I__2963 (
            .O(N__12922),
            .I(N__12885));
    LocalMux I__2962 (
            .O(N__12919),
            .I(N__12885));
    Span4Mux_v I__2961 (
            .O(N__12912),
            .I(N__12885));
    Span4Mux_v I__2960 (
            .O(N__12907),
            .I(N__12885));
    LocalMux I__2959 (
            .O(N__12904),
            .I(N__12882));
    Sp12to4 I__2958 (
            .O(N__12901),
            .I(N__12879));
    Span4Mux_h I__2957 (
            .O(N__12898),
            .I(N__12876));
    SRMux I__2956 (
            .O(N__12897),
            .I(N__12873));
    Span4Mux_h I__2955 (
            .O(N__12894),
            .I(N__12868));
    Span4Mux_v I__2954 (
            .O(N__12885),
            .I(N__12868));
    Span4Mux_h I__2953 (
            .O(N__12882),
            .I(N__12865));
    Span12Mux_v I__2952 (
            .O(N__12879),
            .I(N__12858));
    Sp12to4 I__2951 (
            .O(N__12876),
            .I(N__12858));
    LocalMux I__2950 (
            .O(N__12873),
            .I(N__12858));
    Odrv4 I__2949 (
            .O(N__12868),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2948 (
            .O(N__12865),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2947 (
            .O(N__12858),
            .I(CONSTANT_ONE_NET));
    InMux I__2946 (
            .O(N__12851),
            .I(N__12848));
    LocalMux I__2945 (
            .O(N__12848),
            .I(N__12845));
    Span4Mux_v I__2944 (
            .O(N__12845),
            .I(N__12842));
    Span4Mux_v I__2943 (
            .O(N__12842),
            .I(N__12839));
    Odrv4 I__2942 (
            .O(N__12839),
            .I(\this_vram.mem_out_bus9_5 ));
    InMux I__2941 (
            .O(N__12836),
            .I(N__12833));
    LocalMux I__2940 (
            .O(N__12833),
            .I(N__12830));
    Odrv4 I__2939 (
            .O(N__12830),
            .I(\this_vram.mem_out_bus8_5 ));
    InMux I__2938 (
            .O(N__12827),
            .I(N__12824));
    LocalMux I__2937 (
            .O(N__12824),
            .I(N__12821));
    Span4Mux_v I__2936 (
            .O(N__12821),
            .I(N__12818));
    Sp12to4 I__2935 (
            .O(N__12818),
            .I(N__12815));
    Span12Mux_h I__2934 (
            .O(N__12815),
            .I(N__12812));
    Odrv12 I__2933 (
            .O(N__12812),
            .I(\this_vram.mem_mem_8_2_RNI9H021Z0Z_0 ));
    InMux I__2932 (
            .O(N__12809),
            .I(N__12806));
    LocalMux I__2931 (
            .O(N__12806),
            .I(N__12803));
    Sp12to4 I__2930 (
            .O(N__12803),
            .I(N__12800));
    Span12Mux_v I__2929 (
            .O(N__12800),
            .I(N__12797));
    Odrv12 I__2928 (
            .O(N__12797),
            .I(\this_vram.mem_out_bus5_2 ));
    InMux I__2927 (
            .O(N__12794),
            .I(N__12791));
    LocalMux I__2926 (
            .O(N__12791),
            .I(\this_vram.mem_out_bus7_2 ));
    InMux I__2925 (
            .O(N__12788),
            .I(N__12785));
    LocalMux I__2924 (
            .O(N__12785),
            .I(N__12782));
    Span4Mux_v I__2923 (
            .O(N__12782),
            .I(N__12779));
    Sp12to4 I__2922 (
            .O(N__12779),
            .I(N__12776));
    Span12Mux_h I__2921 (
            .O(N__12776),
            .I(N__12773));
    Odrv12 I__2920 (
            .O(N__12773),
            .I(\this_vram.mem_mem_5_1_RNI38RZ0Z11 ));
    InMux I__2919 (
            .O(N__12770),
            .I(N__12767));
    LocalMux I__2918 (
            .O(N__12767),
            .I(N__12764));
    Sp12to4 I__2917 (
            .O(N__12764),
            .I(N__12761));
    Span12Mux_v I__2916 (
            .O(N__12761),
            .I(N__12758));
    Odrv12 I__2915 (
            .O(N__12758),
            .I(\this_vram.mem_out_bus5_3 ));
    InMux I__2914 (
            .O(N__12755),
            .I(N__12752));
    LocalMux I__2913 (
            .O(N__12752),
            .I(\this_vram.mem_out_bus7_3 ));
    InMux I__2912 (
            .O(N__12749),
            .I(N__12746));
    LocalMux I__2911 (
            .O(N__12746),
            .I(N__12743));
    Span12Mux_s11_h I__2910 (
            .O(N__12743),
            .I(N__12740));
    Span12Mux_h I__2909 (
            .O(N__12740),
            .I(N__12737));
    Odrv12 I__2908 (
            .O(N__12737),
            .I(\this_vram.mem_mem_5_1_RNI38R11Z0Z_0 ));
    CascadeMux I__2907 (
            .O(N__12734),
            .I(\this_vga_signals.N_37_cascade_ ));
    InMux I__2906 (
            .O(N__12731),
            .I(N__12728));
    LocalMux I__2905 (
            .O(N__12728),
            .I(\this_vga_signals.M_hstate_q_ns_i_i_2_0 ));
    CascadeMux I__2904 (
            .O(N__12725),
            .I(N__12722));
    CascadeBuf I__2903 (
            .O(N__12722),
            .I(N__12719));
    CascadeMux I__2902 (
            .O(N__12719),
            .I(N__12716));
    CascadeBuf I__2901 (
            .O(N__12716),
            .I(N__12713));
    CascadeMux I__2900 (
            .O(N__12713),
            .I(N__12709));
    CascadeMux I__2899 (
            .O(N__12712),
            .I(N__12706));
    CascadeBuf I__2898 (
            .O(N__12709),
            .I(N__12703));
    CascadeBuf I__2897 (
            .O(N__12706),
            .I(N__12700));
    CascadeMux I__2896 (
            .O(N__12703),
            .I(N__12697));
    CascadeMux I__2895 (
            .O(N__12700),
            .I(N__12694));
    CascadeBuf I__2894 (
            .O(N__12697),
            .I(N__12691));
    CascadeBuf I__2893 (
            .O(N__12694),
            .I(N__12688));
    CascadeMux I__2892 (
            .O(N__12691),
            .I(N__12685));
    CascadeMux I__2891 (
            .O(N__12688),
            .I(N__12682));
    CascadeBuf I__2890 (
            .O(N__12685),
            .I(N__12679));
    CascadeBuf I__2889 (
            .O(N__12682),
            .I(N__12676));
    CascadeMux I__2888 (
            .O(N__12679),
            .I(N__12673));
    CascadeMux I__2887 (
            .O(N__12676),
            .I(N__12670));
    CascadeBuf I__2886 (
            .O(N__12673),
            .I(N__12667));
    CascadeBuf I__2885 (
            .O(N__12670),
            .I(N__12664));
    CascadeMux I__2884 (
            .O(N__12667),
            .I(N__12661));
    CascadeMux I__2883 (
            .O(N__12664),
            .I(N__12658));
    CascadeBuf I__2882 (
            .O(N__12661),
            .I(N__12655));
    CascadeBuf I__2881 (
            .O(N__12658),
            .I(N__12652));
    CascadeMux I__2880 (
            .O(N__12655),
            .I(N__12649));
    CascadeMux I__2879 (
            .O(N__12652),
            .I(N__12646));
    CascadeBuf I__2878 (
            .O(N__12649),
            .I(N__12643));
    CascadeBuf I__2877 (
            .O(N__12646),
            .I(N__12640));
    CascadeMux I__2876 (
            .O(N__12643),
            .I(N__12637));
    CascadeMux I__2875 (
            .O(N__12640),
            .I(N__12634));
    CascadeBuf I__2874 (
            .O(N__12637),
            .I(N__12631));
    CascadeBuf I__2873 (
            .O(N__12634),
            .I(N__12628));
    CascadeMux I__2872 (
            .O(N__12631),
            .I(N__12625));
    CascadeMux I__2871 (
            .O(N__12628),
            .I(N__12622));
    CascadeBuf I__2870 (
            .O(N__12625),
            .I(N__12619));
    CascadeBuf I__2869 (
            .O(N__12622),
            .I(N__12616));
    CascadeMux I__2868 (
            .O(N__12619),
            .I(N__12613));
    CascadeMux I__2867 (
            .O(N__12616),
            .I(N__12610));
    CascadeBuf I__2866 (
            .O(N__12613),
            .I(N__12607));
    CascadeBuf I__2865 (
            .O(N__12610),
            .I(N__12604));
    CascadeMux I__2864 (
            .O(N__12607),
            .I(N__12601));
    CascadeMux I__2863 (
            .O(N__12604),
            .I(N__12598));
    CascadeBuf I__2862 (
            .O(N__12601),
            .I(N__12595));
    CascadeBuf I__2861 (
            .O(N__12598),
            .I(N__12592));
    CascadeMux I__2860 (
            .O(N__12595),
            .I(N__12589));
    CascadeMux I__2859 (
            .O(N__12592),
            .I(N__12586));
    CascadeBuf I__2858 (
            .O(N__12589),
            .I(N__12583));
    CascadeBuf I__2857 (
            .O(N__12586),
            .I(N__12580));
    CascadeMux I__2856 (
            .O(N__12583),
            .I(N__12577));
    CascadeMux I__2855 (
            .O(N__12580),
            .I(N__12574));
    CascadeBuf I__2854 (
            .O(N__12577),
            .I(N__12571));
    CascadeBuf I__2853 (
            .O(N__12574),
            .I(N__12568));
    CascadeMux I__2852 (
            .O(N__12571),
            .I(N__12565));
    CascadeMux I__2851 (
            .O(N__12568),
            .I(N__12562));
    CascadeBuf I__2850 (
            .O(N__12565),
            .I(N__12559));
    CascadeBuf I__2849 (
            .O(N__12562),
            .I(N__12556));
    CascadeMux I__2848 (
            .O(N__12559),
            .I(N__12553));
    CascadeMux I__2847 (
            .O(N__12556),
            .I(N__12550));
    InMux I__2846 (
            .O(N__12553),
            .I(N__12547));
    InMux I__2845 (
            .O(N__12550),
            .I(N__12544));
    LocalMux I__2844 (
            .O(N__12547),
            .I(N__12541));
    LocalMux I__2843 (
            .O(N__12544),
            .I(N__12536));
    Span4Mux_h I__2842 (
            .O(N__12541),
            .I(N__12533));
    InMux I__2841 (
            .O(N__12540),
            .I(N__12530));
    InMux I__2840 (
            .O(N__12539),
            .I(N__12527));
    Sp12to4 I__2839 (
            .O(N__12536),
            .I(N__12524));
    Span4Mux_h I__2838 (
            .O(N__12533),
            .I(N__12521));
    LocalMux I__2837 (
            .O(N__12530),
            .I(N__12515));
    LocalMux I__2836 (
            .O(N__12527),
            .I(N__12515));
    Span12Mux_s6_v I__2835 (
            .O(N__12524),
            .I(N__12512));
    Sp12to4 I__2834 (
            .O(N__12521),
            .I(N__12509));
    InMux I__2833 (
            .O(N__12520),
            .I(N__12506));
    Span4Mux_v I__2832 (
            .O(N__12515),
            .I(N__12503));
    Span12Mux_h I__2831 (
            .O(N__12512),
            .I(N__12498));
    Span12Mux_s6_v I__2830 (
            .O(N__12509),
            .I(N__12498));
    LocalMux I__2829 (
            .O(N__12506),
            .I(M_this_vga_signals_address_0));
    Odrv4 I__2828 (
            .O(N__12503),
            .I(M_this_vga_signals_address_0));
    Odrv12 I__2827 (
            .O(N__12498),
            .I(M_this_vga_signals_address_0));
    CascadeMux I__2826 (
            .O(N__12491),
            .I(N__12486));
    CascadeMux I__2825 (
            .O(N__12490),
            .I(N__12482));
    InMux I__2824 (
            .O(N__12489),
            .I(N__12479));
    InMux I__2823 (
            .O(N__12486),
            .I(N__12474));
    InMux I__2822 (
            .O(N__12485),
            .I(N__12474));
    InMux I__2821 (
            .O(N__12482),
            .I(N__12471));
    LocalMux I__2820 (
            .O(N__12479),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    LocalMux I__2819 (
            .O(N__12474),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    LocalMux I__2818 (
            .O(N__12471),
            .I(\this_vga_signals.M_hcounter_qZ0Z_11 ));
    CascadeMux I__2817 (
            .O(N__12464),
            .I(N__12461));
    CascadeBuf I__2816 (
            .O(N__12461),
            .I(N__12458));
    CascadeMux I__2815 (
            .O(N__12458),
            .I(N__12455));
    CascadeBuf I__2814 (
            .O(N__12455),
            .I(N__12451));
    CascadeMux I__2813 (
            .O(N__12454),
            .I(N__12448));
    CascadeMux I__2812 (
            .O(N__12451),
            .I(N__12445));
    CascadeBuf I__2811 (
            .O(N__12448),
            .I(N__12442));
    CascadeBuf I__2810 (
            .O(N__12445),
            .I(N__12439));
    CascadeMux I__2809 (
            .O(N__12442),
            .I(N__12436));
    CascadeMux I__2808 (
            .O(N__12439),
            .I(N__12433));
    CascadeBuf I__2807 (
            .O(N__12436),
            .I(N__12430));
    CascadeBuf I__2806 (
            .O(N__12433),
            .I(N__12427));
    CascadeMux I__2805 (
            .O(N__12430),
            .I(N__12424));
    CascadeMux I__2804 (
            .O(N__12427),
            .I(N__12421));
    CascadeBuf I__2803 (
            .O(N__12424),
            .I(N__12418));
    CascadeBuf I__2802 (
            .O(N__12421),
            .I(N__12415));
    CascadeMux I__2801 (
            .O(N__12418),
            .I(N__12412));
    CascadeMux I__2800 (
            .O(N__12415),
            .I(N__12409));
    CascadeBuf I__2799 (
            .O(N__12412),
            .I(N__12406));
    CascadeBuf I__2798 (
            .O(N__12409),
            .I(N__12403));
    CascadeMux I__2797 (
            .O(N__12406),
            .I(N__12400));
    CascadeMux I__2796 (
            .O(N__12403),
            .I(N__12397));
    CascadeBuf I__2795 (
            .O(N__12400),
            .I(N__12394));
    CascadeBuf I__2794 (
            .O(N__12397),
            .I(N__12391));
    CascadeMux I__2793 (
            .O(N__12394),
            .I(N__12388));
    CascadeMux I__2792 (
            .O(N__12391),
            .I(N__12385));
    CascadeBuf I__2791 (
            .O(N__12388),
            .I(N__12382));
    CascadeBuf I__2790 (
            .O(N__12385),
            .I(N__12379));
    CascadeMux I__2789 (
            .O(N__12382),
            .I(N__12376));
    CascadeMux I__2788 (
            .O(N__12379),
            .I(N__12373));
    CascadeBuf I__2787 (
            .O(N__12376),
            .I(N__12370));
    CascadeBuf I__2786 (
            .O(N__12373),
            .I(N__12367));
    CascadeMux I__2785 (
            .O(N__12370),
            .I(N__12364));
    CascadeMux I__2784 (
            .O(N__12367),
            .I(N__12361));
    CascadeBuf I__2783 (
            .O(N__12364),
            .I(N__12358));
    CascadeBuf I__2782 (
            .O(N__12361),
            .I(N__12355));
    CascadeMux I__2781 (
            .O(N__12358),
            .I(N__12352));
    CascadeMux I__2780 (
            .O(N__12355),
            .I(N__12349));
    CascadeBuf I__2779 (
            .O(N__12352),
            .I(N__12346));
    CascadeBuf I__2778 (
            .O(N__12349),
            .I(N__12343));
    CascadeMux I__2777 (
            .O(N__12346),
            .I(N__12340));
    CascadeMux I__2776 (
            .O(N__12343),
            .I(N__12337));
    CascadeBuf I__2775 (
            .O(N__12340),
            .I(N__12334));
    CascadeBuf I__2774 (
            .O(N__12337),
            .I(N__12331));
    CascadeMux I__2773 (
            .O(N__12334),
            .I(N__12328));
    CascadeMux I__2772 (
            .O(N__12331),
            .I(N__12325));
    CascadeBuf I__2771 (
            .O(N__12328),
            .I(N__12322));
    CascadeBuf I__2770 (
            .O(N__12325),
            .I(N__12319));
    CascadeMux I__2769 (
            .O(N__12322),
            .I(N__12316));
    CascadeMux I__2768 (
            .O(N__12319),
            .I(N__12313));
    CascadeBuf I__2767 (
            .O(N__12316),
            .I(N__12310));
    CascadeBuf I__2766 (
            .O(N__12313),
            .I(N__12307));
    CascadeMux I__2765 (
            .O(N__12310),
            .I(N__12304));
    CascadeMux I__2764 (
            .O(N__12307),
            .I(N__12301));
    CascadeBuf I__2763 (
            .O(N__12304),
            .I(N__12298));
    CascadeBuf I__2762 (
            .O(N__12301),
            .I(N__12295));
    CascadeMux I__2761 (
            .O(N__12298),
            .I(N__12292));
    CascadeMux I__2760 (
            .O(N__12295),
            .I(N__12289));
    InMux I__2759 (
            .O(N__12292),
            .I(N__12285));
    InMux I__2758 (
            .O(N__12289),
            .I(N__12282));
    CascadeMux I__2757 (
            .O(N__12288),
            .I(N__12279));
    LocalMux I__2756 (
            .O(N__12285),
            .I(N__12275));
    LocalMux I__2755 (
            .O(N__12282),
            .I(N__12272));
    InMux I__2754 (
            .O(N__12279),
            .I(N__12266));
    InMux I__2753 (
            .O(N__12278),
            .I(N__12266));
    Span12Mux_h I__2752 (
            .O(N__12275),
            .I(N__12263));
    Span12Mux_h I__2751 (
            .O(N__12272),
            .I(N__12260));
    InMux I__2750 (
            .O(N__12271),
            .I(N__12257));
    LocalMux I__2749 (
            .O(N__12266),
            .I(N__12254));
    Span12Mux_v I__2748 (
            .O(N__12263),
            .I(N__12251));
    Span12Mux_v I__2747 (
            .O(N__12260),
            .I(N__12248));
    LocalMux I__2746 (
            .O(N__12257),
            .I(M_this_vga_signals_address_1));
    Odrv4 I__2745 (
            .O(N__12254),
            .I(M_this_vga_signals_address_1));
    Odrv12 I__2744 (
            .O(N__12251),
            .I(M_this_vga_signals_address_1));
    Odrv12 I__2743 (
            .O(N__12248),
            .I(M_this_vga_signals_address_1));
    CascadeMux I__2742 (
            .O(N__12239),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa_0_a2_0_a2_0_cascade_ ));
    InMux I__2741 (
            .O(N__12236),
            .I(N__12230));
    InMux I__2740 (
            .O(N__12235),
            .I(N__12230));
    LocalMux I__2739 (
            .O(N__12230),
            .I(\this_vga_signals.N_169_4 ));
    InMux I__2738 (
            .O(N__12227),
            .I(N__12220));
    CascadeMux I__2737 (
            .O(N__12226),
            .I(N__12217));
    InMux I__2736 (
            .O(N__12225),
            .I(N__12214));
    InMux I__2735 (
            .O(N__12224),
            .I(N__12211));
    InMux I__2734 (
            .O(N__12223),
            .I(N__12208));
    LocalMux I__2733 (
            .O(N__12220),
            .I(N__12205));
    InMux I__2732 (
            .O(N__12217),
            .I(N__12202));
    LocalMux I__2731 (
            .O(N__12214),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    LocalMux I__2730 (
            .O(N__12211),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    LocalMux I__2729 (
            .O(N__12208),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    Odrv4 I__2728 (
            .O(N__12205),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    LocalMux I__2727 (
            .O(N__12202),
            .I(\this_vga_signals.M_hstate_d_0_sqmuxa ));
    InMux I__2726 (
            .O(N__12191),
            .I(N__12188));
    LocalMux I__2725 (
            .O(N__12188),
            .I(N__12184));
    InMux I__2724 (
            .O(N__12187),
            .I(N__12181));
    Odrv4 I__2723 (
            .O(N__12184),
            .I(\this_vga_signals.N_169 ));
    LocalMux I__2722 (
            .O(N__12181),
            .I(\this_vga_signals.N_169 ));
    InMux I__2721 (
            .O(N__12176),
            .I(N__12172));
    InMux I__2720 (
            .O(N__12175),
            .I(N__12169));
    LocalMux I__2719 (
            .O(N__12172),
            .I(\this_vga_signals.N_42 ));
    LocalMux I__2718 (
            .O(N__12169),
            .I(\this_vga_signals.N_42 ));
    InMux I__2717 (
            .O(N__12164),
            .I(N__12158));
    InMux I__2716 (
            .O(N__12163),
            .I(N__12158));
    LocalMux I__2715 (
            .O(N__12158),
            .I(\this_vga_signals.N_46 ));
    CascadeMux I__2714 (
            .O(N__12155),
            .I(N__12152));
    InMux I__2713 (
            .O(N__12152),
            .I(N__12143));
    InMux I__2712 (
            .O(N__12151),
            .I(N__12143));
    InMux I__2711 (
            .O(N__12150),
            .I(N__12143));
    LocalMux I__2710 (
            .O(N__12143),
            .I(\this_vga_signals.N_83 ));
    InMux I__2709 (
            .O(N__12140),
            .I(N__12136));
    InMux I__2708 (
            .O(N__12139),
            .I(N__12133));
    LocalMux I__2707 (
            .O(N__12136),
            .I(N__12130));
    LocalMux I__2706 (
            .O(N__12133),
            .I(N__12127));
    Span4Mux_v I__2705 (
            .O(N__12130),
            .I(N__12121));
    Span4Mux_v I__2704 (
            .O(N__12127),
            .I(N__12121));
    InMux I__2703 (
            .O(N__12126),
            .I(N__12118));
    Span4Mux_h I__2702 (
            .O(N__12121),
            .I(N__12115));
    LocalMux I__2701 (
            .O(N__12118),
            .I(N__12112));
    Sp12to4 I__2700 (
            .O(N__12115),
            .I(N__12102));
    Span12Mux_s5_h I__2699 (
            .O(N__12112),
            .I(N__12102));
    InMux I__2698 (
            .O(N__12111),
            .I(N__12099));
    InMux I__2697 (
            .O(N__12110),
            .I(N__12090));
    InMux I__2696 (
            .O(N__12109),
            .I(N__12090));
    InMux I__2695 (
            .O(N__12108),
            .I(N__12090));
    InMux I__2694 (
            .O(N__12107),
            .I(N__12090));
    Odrv12 I__2693 (
            .O(N__12102),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    LocalMux I__2692 (
            .O(N__12099),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    LocalMux I__2691 (
            .O(N__12090),
            .I(\this_vga_signals.M_hstate_qZ0Z_1 ));
    InMux I__2690 (
            .O(N__12083),
            .I(N__12080));
    LocalMux I__2689 (
            .O(N__12080),
            .I(\this_vga_signals.N_27 ));
    InMux I__2688 (
            .O(N__12077),
            .I(N__12071));
    InMux I__2687 (
            .O(N__12076),
            .I(N__12071));
    LocalMux I__2686 (
            .O(N__12071),
            .I(N__12067));
    IoInMux I__2685 (
            .O(N__12070),
            .I(N__12062));
    Span4Mux_v I__2684 (
            .O(N__12067),
            .I(N__12059));
    InMux I__2683 (
            .O(N__12066),
            .I(N__12056));
    CascadeMux I__2682 (
            .O(N__12065),
            .I(N__12053));
    LocalMux I__2681 (
            .O(N__12062),
            .I(N__12050));
    Span4Mux_h I__2680 (
            .O(N__12059),
            .I(N__12047));
    LocalMux I__2679 (
            .O(N__12056),
            .I(N__12044));
    InMux I__2678 (
            .O(N__12053),
            .I(N__12041));
    Span12Mux_s11_v I__2677 (
            .O(N__12050),
            .I(N__12038));
    Odrv4 I__2676 (
            .O(N__12047),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__2675 (
            .O(N__12044),
            .I(M_this_reset_cond_out_0));
    LocalMux I__2674 (
            .O(N__12041),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__2673 (
            .O(N__12038),
            .I(M_this_reset_cond_out_0));
    InMux I__2672 (
            .O(N__12029),
            .I(N__12026));
    LocalMux I__2671 (
            .O(N__12026),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__2670 (
            .O(N__12023),
            .I(N__12020));
    LocalMux I__2669 (
            .O(N__12020),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__2668 (
            .O(N__12017),
            .I(N__12012));
    InMux I__2667 (
            .O(N__12016),
            .I(N__12006));
    InMux I__2666 (
            .O(N__12015),
            .I(N__12006));
    LocalMux I__2665 (
            .O(N__12012),
            .I(N__12003));
    InMux I__2664 (
            .O(N__12011),
            .I(N__12000));
    LocalMux I__2663 (
            .O(N__12006),
            .I(N__11997));
    Odrv4 I__2662 (
            .O(N__12003),
            .I(\this_vga_signals.N_68 ));
    LocalMux I__2661 (
            .O(N__12000),
            .I(\this_vga_signals.N_68 ));
    Odrv4 I__2660 (
            .O(N__11997),
            .I(\this_vga_signals.N_68 ));
    InMux I__2659 (
            .O(N__11990),
            .I(bfn_14_20_0_));
    InMux I__2658 (
            .O(N__11987),
            .I(N__11981));
    InMux I__2657 (
            .O(N__11986),
            .I(N__11978));
    CascadeMux I__2656 (
            .O(N__11985),
            .I(N__11975));
    InMux I__2655 (
            .O(N__11984),
            .I(N__11972));
    LocalMux I__2654 (
            .O(N__11981),
            .I(N__11968));
    LocalMux I__2653 (
            .O(N__11978),
            .I(N__11965));
    InMux I__2652 (
            .O(N__11975),
            .I(N__11962));
    LocalMux I__2651 (
            .O(N__11972),
            .I(N__11959));
    InMux I__2650 (
            .O(N__11971),
            .I(N__11956));
    Span4Mux_v I__2649 (
            .O(N__11968),
            .I(N__11951));
    Span4Mux_h I__2648 (
            .O(N__11965),
            .I(N__11951));
    LocalMux I__2647 (
            .O(N__11962),
            .I(N__11948));
    Span4Mux_h I__2646 (
            .O(N__11959),
            .I(N__11945));
    LocalMux I__2645 (
            .O(N__11956),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2644 (
            .O(N__11951),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2643 (
            .O(N__11948),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__2642 (
            .O(N__11945),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    CascadeMux I__2641 (
            .O(N__11936),
            .I(N__11930));
    CascadeMux I__2640 (
            .O(N__11935),
            .I(N__11926));
    CascadeMux I__2639 (
            .O(N__11934),
            .I(N__11923));
    InMux I__2638 (
            .O(N__11933),
            .I(N__11918));
    InMux I__2637 (
            .O(N__11930),
            .I(N__11918));
    InMux I__2636 (
            .O(N__11929),
            .I(N__11915));
    InMux I__2635 (
            .O(N__11926),
            .I(N__11912));
    InMux I__2634 (
            .O(N__11923),
            .I(N__11909));
    LocalMux I__2633 (
            .O(N__11918),
            .I(N__11901));
    LocalMux I__2632 (
            .O(N__11915),
            .I(N__11898));
    LocalMux I__2631 (
            .O(N__11912),
            .I(N__11895));
    LocalMux I__2630 (
            .O(N__11909),
            .I(N__11892));
    SRMux I__2629 (
            .O(N__11908),
            .I(N__11873));
    SRMux I__2628 (
            .O(N__11907),
            .I(N__11873));
    SRMux I__2627 (
            .O(N__11906),
            .I(N__11873));
    SRMux I__2626 (
            .O(N__11905),
            .I(N__11873));
    SRMux I__2625 (
            .O(N__11904),
            .I(N__11873));
    Glb2LocalMux I__2624 (
            .O(N__11901),
            .I(N__11873));
    Glb2LocalMux I__2623 (
            .O(N__11898),
            .I(N__11873));
    Glb2LocalMux I__2622 (
            .O(N__11895),
            .I(N__11873));
    Glb2LocalMux I__2621 (
            .O(N__11892),
            .I(N__11873));
    GlobalMux I__2620 (
            .O(N__11873),
            .I(N__11870));
    gio2CtrlBuf I__2619 (
            .O(N__11870),
            .I(N_112_g));
    InMux I__2618 (
            .O(N__11867),
            .I(N__11859));
    InMux I__2617 (
            .O(N__11866),
            .I(N__11859));
    InMux I__2616 (
            .O(N__11865),
            .I(N__11856));
    InMux I__2615 (
            .O(N__11864),
            .I(N__11853));
    LocalMux I__2614 (
            .O(N__11859),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2613 (
            .O(N__11856),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2612 (
            .O(N__11853),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    InMux I__2611 (
            .O(N__11846),
            .I(N__11842));
    InMux I__2610 (
            .O(N__11845),
            .I(N__11839));
    LocalMux I__2609 (
            .O(N__11842),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2608 (
            .O(N__11839),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    CascadeMux I__2607 (
            .O(N__11834),
            .I(N__11829));
    CascadeMux I__2606 (
            .O(N__11833),
            .I(N__11826));
    InMux I__2605 (
            .O(N__11832),
            .I(N__11823));
    InMux I__2604 (
            .O(N__11829),
            .I(N__11820));
    InMux I__2603 (
            .O(N__11826),
            .I(N__11817));
    LocalMux I__2602 (
            .O(N__11823),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2601 (
            .O(N__11820),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2600 (
            .O(N__11817),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__2599 (
            .O(N__11810),
            .I(N__11806));
    InMux I__2598 (
            .O(N__11809),
            .I(N__11803));
    LocalMux I__2597 (
            .O(N__11806),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2596 (
            .O(N__11803),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__2595 (
            .O(N__11798),
            .I(N__11794));
    InMux I__2594 (
            .O(N__11797),
            .I(N__11791));
    LocalMux I__2593 (
            .O(N__11794),
            .I(N__11788));
    LocalMux I__2592 (
            .O(N__11791),
            .I(N__11785));
    Span4Mux_v I__2591 (
            .O(N__11788),
            .I(N__11779));
    Span4Mux_v I__2590 (
            .O(N__11785),
            .I(N__11779));
    InMux I__2589 (
            .O(N__11784),
            .I(N__11776));
    Sp12to4 I__2588 (
            .O(N__11779),
            .I(N__11771));
    LocalMux I__2587 (
            .O(N__11776),
            .I(N__11771));
    Span12Mux_s10_h I__2586 (
            .O(N__11771),
            .I(N__11764));
    InMux I__2585 (
            .O(N__11770),
            .I(N__11757));
    InMux I__2584 (
            .O(N__11769),
            .I(N__11757));
    InMux I__2583 (
            .O(N__11768),
            .I(N__11757));
    InMux I__2582 (
            .O(N__11767),
            .I(N__11754));
    Odrv12 I__2581 (
            .O(N__11764),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    LocalMux I__2580 (
            .O(N__11757),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    LocalMux I__2579 (
            .O(N__11754),
            .I(\this_vga_signals.M_hstate_qZ0Z_0 ));
    CascadeMux I__2578 (
            .O(N__11747),
            .I(N__11741));
    CascadeMux I__2577 (
            .O(N__11746),
            .I(N__11737));
    InMux I__2576 (
            .O(N__11745),
            .I(N__11734));
    InMux I__2575 (
            .O(N__11744),
            .I(N__11731));
    InMux I__2574 (
            .O(N__11741),
            .I(N__11728));
    InMux I__2573 (
            .O(N__11740),
            .I(N__11723));
    InMux I__2572 (
            .O(N__11737),
            .I(N__11723));
    LocalMux I__2571 (
            .O(N__11734),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2570 (
            .O(N__11731),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2569 (
            .O(N__11728),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2568 (
            .O(N__11723),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    CascadeMux I__2567 (
            .O(N__11714),
            .I(N__11708));
    CascadeMux I__2566 (
            .O(N__11713),
            .I(N__11705));
    CascadeMux I__2565 (
            .O(N__11712),
            .I(N__11701));
    InMux I__2564 (
            .O(N__11711),
            .I(N__11698));
    InMux I__2563 (
            .O(N__11708),
            .I(N__11695));
    InMux I__2562 (
            .O(N__11705),
            .I(N__11690));
    InMux I__2561 (
            .O(N__11704),
            .I(N__11690));
    InMux I__2560 (
            .O(N__11701),
            .I(N__11687));
    LocalMux I__2559 (
            .O(N__11698),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    LocalMux I__2558 (
            .O(N__11695),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    LocalMux I__2557 (
            .O(N__11690),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    LocalMux I__2556 (
            .O(N__11687),
            .I(\this_vga_signals.M_hcounter_qZ0Z_10 ));
    CascadeMux I__2555 (
            .O(N__11678),
            .I(N__11675));
    CascadeBuf I__2554 (
            .O(N__11675),
            .I(N__11672));
    CascadeMux I__2553 (
            .O(N__11672),
            .I(N__11669));
    CascadeBuf I__2552 (
            .O(N__11669),
            .I(N__11666));
    CascadeMux I__2551 (
            .O(N__11666),
            .I(N__11663));
    CascadeBuf I__2550 (
            .O(N__11663),
            .I(N__11660));
    CascadeMux I__2549 (
            .O(N__11660),
            .I(N__11656));
    CascadeMux I__2548 (
            .O(N__11659),
            .I(N__11653));
    CascadeBuf I__2547 (
            .O(N__11656),
            .I(N__11650));
    CascadeBuf I__2546 (
            .O(N__11653),
            .I(N__11647));
    CascadeMux I__2545 (
            .O(N__11650),
            .I(N__11644));
    CascadeMux I__2544 (
            .O(N__11647),
            .I(N__11641));
    CascadeBuf I__2543 (
            .O(N__11644),
            .I(N__11638));
    CascadeBuf I__2542 (
            .O(N__11641),
            .I(N__11635));
    CascadeMux I__2541 (
            .O(N__11638),
            .I(N__11632));
    CascadeMux I__2540 (
            .O(N__11635),
            .I(N__11629));
    CascadeBuf I__2539 (
            .O(N__11632),
            .I(N__11626));
    CascadeBuf I__2538 (
            .O(N__11629),
            .I(N__11623));
    CascadeMux I__2537 (
            .O(N__11626),
            .I(N__11620));
    CascadeMux I__2536 (
            .O(N__11623),
            .I(N__11617));
    CascadeBuf I__2535 (
            .O(N__11620),
            .I(N__11614));
    CascadeBuf I__2534 (
            .O(N__11617),
            .I(N__11611));
    CascadeMux I__2533 (
            .O(N__11614),
            .I(N__11608));
    CascadeMux I__2532 (
            .O(N__11611),
            .I(N__11605));
    CascadeBuf I__2531 (
            .O(N__11608),
            .I(N__11602));
    CascadeBuf I__2530 (
            .O(N__11605),
            .I(N__11599));
    CascadeMux I__2529 (
            .O(N__11602),
            .I(N__11596));
    CascadeMux I__2528 (
            .O(N__11599),
            .I(N__11593));
    CascadeBuf I__2527 (
            .O(N__11596),
            .I(N__11590));
    CascadeBuf I__2526 (
            .O(N__11593),
            .I(N__11587));
    CascadeMux I__2525 (
            .O(N__11590),
            .I(N__11584));
    CascadeMux I__2524 (
            .O(N__11587),
            .I(N__11581));
    CascadeBuf I__2523 (
            .O(N__11584),
            .I(N__11578));
    CascadeBuf I__2522 (
            .O(N__11581),
            .I(N__11575));
    CascadeMux I__2521 (
            .O(N__11578),
            .I(N__11572));
    CascadeMux I__2520 (
            .O(N__11575),
            .I(N__11569));
    CascadeBuf I__2519 (
            .O(N__11572),
            .I(N__11566));
    CascadeBuf I__2518 (
            .O(N__11569),
            .I(N__11563));
    CascadeMux I__2517 (
            .O(N__11566),
            .I(N__11560));
    CascadeMux I__2516 (
            .O(N__11563),
            .I(N__11557));
    CascadeBuf I__2515 (
            .O(N__11560),
            .I(N__11554));
    CascadeBuf I__2514 (
            .O(N__11557),
            .I(N__11551));
    CascadeMux I__2513 (
            .O(N__11554),
            .I(N__11548));
    CascadeMux I__2512 (
            .O(N__11551),
            .I(N__11545));
    CascadeBuf I__2511 (
            .O(N__11548),
            .I(N__11542));
    CascadeBuf I__2510 (
            .O(N__11545),
            .I(N__11539));
    CascadeMux I__2509 (
            .O(N__11542),
            .I(N__11536));
    CascadeMux I__2508 (
            .O(N__11539),
            .I(N__11533));
    CascadeBuf I__2507 (
            .O(N__11536),
            .I(N__11530));
    CascadeBuf I__2506 (
            .O(N__11533),
            .I(N__11527));
    CascadeMux I__2505 (
            .O(N__11530),
            .I(N__11524));
    CascadeMux I__2504 (
            .O(N__11527),
            .I(N__11521));
    CascadeBuf I__2503 (
            .O(N__11524),
            .I(N__11518));
    CascadeBuf I__2502 (
            .O(N__11521),
            .I(N__11515));
    CascadeMux I__2501 (
            .O(N__11518),
            .I(N__11512));
    CascadeMux I__2500 (
            .O(N__11515),
            .I(N__11509));
    InMux I__2499 (
            .O(N__11512),
            .I(N__11506));
    CascadeBuf I__2498 (
            .O(N__11509),
            .I(N__11503));
    LocalMux I__2497 (
            .O(N__11506),
            .I(N__11500));
    CascadeMux I__2496 (
            .O(N__11503),
            .I(N__11497));
    Span4Mux_h I__2495 (
            .O(N__11500),
            .I(N__11494));
    InMux I__2494 (
            .O(N__11497),
            .I(N__11490));
    Span4Mux_h I__2493 (
            .O(N__11494),
            .I(N__11487));
    InMux I__2492 (
            .O(N__11493),
            .I(N__11482));
    LocalMux I__2491 (
            .O(N__11490),
            .I(N__11478));
    Sp12to4 I__2490 (
            .O(N__11487),
            .I(N__11475));
    InMux I__2489 (
            .O(N__11486),
            .I(N__11470));
    InMux I__2488 (
            .O(N__11485),
            .I(N__11470));
    LocalMux I__2487 (
            .O(N__11482),
            .I(N__11467));
    InMux I__2486 (
            .O(N__11481),
            .I(N__11464));
    Span12Mux_v I__2485 (
            .O(N__11478),
            .I(N__11461));
    Span12Mux_v I__2484 (
            .O(N__11475),
            .I(N__11458));
    LocalMux I__2483 (
            .O(N__11470),
            .I(M_this_vga_signals_address_2));
    Odrv4 I__2482 (
            .O(N__11467),
            .I(M_this_vga_signals_address_2));
    LocalMux I__2481 (
            .O(N__11464),
            .I(M_this_vga_signals_address_2));
    Odrv12 I__2480 (
            .O(N__11461),
            .I(M_this_vga_signals_address_2));
    Odrv12 I__2479 (
            .O(N__11458),
            .I(M_this_vga_signals_address_2));
    CascadeMux I__2478 (
            .O(N__11447),
            .I(N__11444));
    CascadeBuf I__2477 (
            .O(N__11444),
            .I(N__11441));
    CascadeMux I__2476 (
            .O(N__11441),
            .I(N__11438));
    CascadeBuf I__2475 (
            .O(N__11438),
            .I(N__11435));
    CascadeMux I__2474 (
            .O(N__11435),
            .I(N__11432));
    CascadeBuf I__2473 (
            .O(N__11432),
            .I(N__11428));
    CascadeMux I__2472 (
            .O(N__11431),
            .I(N__11425));
    CascadeMux I__2471 (
            .O(N__11428),
            .I(N__11422));
    CascadeBuf I__2470 (
            .O(N__11425),
            .I(N__11419));
    CascadeBuf I__2469 (
            .O(N__11422),
            .I(N__11416));
    CascadeMux I__2468 (
            .O(N__11419),
            .I(N__11413));
    CascadeMux I__2467 (
            .O(N__11416),
            .I(N__11410));
    CascadeBuf I__2466 (
            .O(N__11413),
            .I(N__11407));
    CascadeBuf I__2465 (
            .O(N__11410),
            .I(N__11404));
    CascadeMux I__2464 (
            .O(N__11407),
            .I(N__11401));
    CascadeMux I__2463 (
            .O(N__11404),
            .I(N__11398));
    CascadeBuf I__2462 (
            .O(N__11401),
            .I(N__11395));
    CascadeBuf I__2461 (
            .O(N__11398),
            .I(N__11392));
    CascadeMux I__2460 (
            .O(N__11395),
            .I(N__11389));
    CascadeMux I__2459 (
            .O(N__11392),
            .I(N__11386));
    CascadeBuf I__2458 (
            .O(N__11389),
            .I(N__11383));
    CascadeBuf I__2457 (
            .O(N__11386),
            .I(N__11380));
    CascadeMux I__2456 (
            .O(N__11383),
            .I(N__11377));
    CascadeMux I__2455 (
            .O(N__11380),
            .I(N__11374));
    CascadeBuf I__2454 (
            .O(N__11377),
            .I(N__11371));
    CascadeBuf I__2453 (
            .O(N__11374),
            .I(N__11368));
    CascadeMux I__2452 (
            .O(N__11371),
            .I(N__11365));
    CascadeMux I__2451 (
            .O(N__11368),
            .I(N__11362));
    CascadeBuf I__2450 (
            .O(N__11365),
            .I(N__11359));
    CascadeBuf I__2449 (
            .O(N__11362),
            .I(N__11356));
    CascadeMux I__2448 (
            .O(N__11359),
            .I(N__11353));
    CascadeMux I__2447 (
            .O(N__11356),
            .I(N__11350));
    CascadeBuf I__2446 (
            .O(N__11353),
            .I(N__11347));
    CascadeBuf I__2445 (
            .O(N__11350),
            .I(N__11344));
    CascadeMux I__2444 (
            .O(N__11347),
            .I(N__11341));
    CascadeMux I__2443 (
            .O(N__11344),
            .I(N__11338));
    CascadeBuf I__2442 (
            .O(N__11341),
            .I(N__11335));
    CascadeBuf I__2441 (
            .O(N__11338),
            .I(N__11332));
    CascadeMux I__2440 (
            .O(N__11335),
            .I(N__11329));
    CascadeMux I__2439 (
            .O(N__11332),
            .I(N__11326));
    CascadeBuf I__2438 (
            .O(N__11329),
            .I(N__11323));
    CascadeBuf I__2437 (
            .O(N__11326),
            .I(N__11320));
    CascadeMux I__2436 (
            .O(N__11323),
            .I(N__11317));
    CascadeMux I__2435 (
            .O(N__11320),
            .I(N__11314));
    CascadeBuf I__2434 (
            .O(N__11317),
            .I(N__11311));
    CascadeBuf I__2433 (
            .O(N__11314),
            .I(N__11308));
    CascadeMux I__2432 (
            .O(N__11311),
            .I(N__11305));
    CascadeMux I__2431 (
            .O(N__11308),
            .I(N__11302));
    CascadeBuf I__2430 (
            .O(N__11305),
            .I(N__11299));
    CascadeBuf I__2429 (
            .O(N__11302),
            .I(N__11296));
    CascadeMux I__2428 (
            .O(N__11299),
            .I(N__11293));
    CascadeMux I__2427 (
            .O(N__11296),
            .I(N__11290));
    CascadeBuf I__2426 (
            .O(N__11293),
            .I(N__11287));
    CascadeBuf I__2425 (
            .O(N__11290),
            .I(N__11284));
    CascadeMux I__2424 (
            .O(N__11287),
            .I(N__11281));
    CascadeMux I__2423 (
            .O(N__11284),
            .I(N__11278));
    CascadeBuf I__2422 (
            .O(N__11281),
            .I(N__11275));
    InMux I__2421 (
            .O(N__11278),
            .I(N__11272));
    CascadeMux I__2420 (
            .O(N__11275),
            .I(N__11269));
    LocalMux I__2419 (
            .O(N__11272),
            .I(N__11266));
    InMux I__2418 (
            .O(N__11269),
            .I(N__11263));
    Span4Mux_h I__2417 (
            .O(N__11266),
            .I(N__11260));
    LocalMux I__2416 (
            .O(N__11263),
            .I(N__11256));
    Span4Mux_h I__2415 (
            .O(N__11260),
            .I(N__11252));
    InMux I__2414 (
            .O(N__11259),
            .I(N__11247));
    Span12Mux_s8_h I__2413 (
            .O(N__11256),
            .I(N__11244));
    InMux I__2412 (
            .O(N__11255),
            .I(N__11241));
    Sp12to4 I__2411 (
            .O(N__11252),
            .I(N__11238));
    InMux I__2410 (
            .O(N__11251),
            .I(N__11235));
    InMux I__2409 (
            .O(N__11250),
            .I(N__11232));
    LocalMux I__2408 (
            .O(N__11247),
            .I(N__11229));
    Span12Mux_v I__2407 (
            .O(N__11244),
            .I(N__11226));
    LocalMux I__2406 (
            .O(N__11241),
            .I(N__11221));
    Span12Mux_s11_v I__2405 (
            .O(N__11238),
            .I(N__11221));
    LocalMux I__2404 (
            .O(N__11235),
            .I(M_this_vga_signals_address_3));
    LocalMux I__2403 (
            .O(N__11232),
            .I(M_this_vga_signals_address_3));
    Odrv4 I__2402 (
            .O(N__11229),
            .I(M_this_vga_signals_address_3));
    Odrv12 I__2401 (
            .O(N__11226),
            .I(M_this_vga_signals_address_3));
    Odrv12 I__2400 (
            .O(N__11221),
            .I(M_this_vga_signals_address_3));
    CascadeMux I__2399 (
            .O(N__11210),
            .I(N__11207));
    CascadeBuf I__2398 (
            .O(N__11207),
            .I(N__11204));
    CascadeMux I__2397 (
            .O(N__11204),
            .I(N__11201));
    CascadeBuf I__2396 (
            .O(N__11201),
            .I(N__11198));
    CascadeMux I__2395 (
            .O(N__11198),
            .I(N__11195));
    CascadeBuf I__2394 (
            .O(N__11195),
            .I(N__11191));
    CascadeMux I__2393 (
            .O(N__11194),
            .I(N__11188));
    CascadeMux I__2392 (
            .O(N__11191),
            .I(N__11185));
    CascadeBuf I__2391 (
            .O(N__11188),
            .I(N__11182));
    CascadeBuf I__2390 (
            .O(N__11185),
            .I(N__11179));
    CascadeMux I__2389 (
            .O(N__11182),
            .I(N__11176));
    CascadeMux I__2388 (
            .O(N__11179),
            .I(N__11173));
    CascadeBuf I__2387 (
            .O(N__11176),
            .I(N__11170));
    CascadeBuf I__2386 (
            .O(N__11173),
            .I(N__11167));
    CascadeMux I__2385 (
            .O(N__11170),
            .I(N__11164));
    CascadeMux I__2384 (
            .O(N__11167),
            .I(N__11161));
    CascadeBuf I__2383 (
            .O(N__11164),
            .I(N__11158));
    CascadeBuf I__2382 (
            .O(N__11161),
            .I(N__11155));
    CascadeMux I__2381 (
            .O(N__11158),
            .I(N__11152));
    CascadeMux I__2380 (
            .O(N__11155),
            .I(N__11149));
    CascadeBuf I__2379 (
            .O(N__11152),
            .I(N__11146));
    CascadeBuf I__2378 (
            .O(N__11149),
            .I(N__11143));
    CascadeMux I__2377 (
            .O(N__11146),
            .I(N__11140));
    CascadeMux I__2376 (
            .O(N__11143),
            .I(N__11137));
    CascadeBuf I__2375 (
            .O(N__11140),
            .I(N__11134));
    CascadeBuf I__2374 (
            .O(N__11137),
            .I(N__11131));
    CascadeMux I__2373 (
            .O(N__11134),
            .I(N__11128));
    CascadeMux I__2372 (
            .O(N__11131),
            .I(N__11125));
    CascadeBuf I__2371 (
            .O(N__11128),
            .I(N__11122));
    CascadeBuf I__2370 (
            .O(N__11125),
            .I(N__11119));
    CascadeMux I__2369 (
            .O(N__11122),
            .I(N__11116));
    CascadeMux I__2368 (
            .O(N__11119),
            .I(N__11113));
    CascadeBuf I__2367 (
            .O(N__11116),
            .I(N__11110));
    CascadeBuf I__2366 (
            .O(N__11113),
            .I(N__11107));
    CascadeMux I__2365 (
            .O(N__11110),
            .I(N__11104));
    CascadeMux I__2364 (
            .O(N__11107),
            .I(N__11101));
    CascadeBuf I__2363 (
            .O(N__11104),
            .I(N__11098));
    CascadeBuf I__2362 (
            .O(N__11101),
            .I(N__11095));
    CascadeMux I__2361 (
            .O(N__11098),
            .I(N__11092));
    CascadeMux I__2360 (
            .O(N__11095),
            .I(N__11089));
    CascadeBuf I__2359 (
            .O(N__11092),
            .I(N__11086));
    CascadeBuf I__2358 (
            .O(N__11089),
            .I(N__11083));
    CascadeMux I__2357 (
            .O(N__11086),
            .I(N__11080));
    CascadeMux I__2356 (
            .O(N__11083),
            .I(N__11077));
    CascadeBuf I__2355 (
            .O(N__11080),
            .I(N__11074));
    CascadeBuf I__2354 (
            .O(N__11077),
            .I(N__11071));
    CascadeMux I__2353 (
            .O(N__11074),
            .I(N__11068));
    CascadeMux I__2352 (
            .O(N__11071),
            .I(N__11065));
    CascadeBuf I__2351 (
            .O(N__11068),
            .I(N__11062));
    CascadeBuf I__2350 (
            .O(N__11065),
            .I(N__11059));
    CascadeMux I__2349 (
            .O(N__11062),
            .I(N__11056));
    CascadeMux I__2348 (
            .O(N__11059),
            .I(N__11053));
    CascadeBuf I__2347 (
            .O(N__11056),
            .I(N__11050));
    CascadeBuf I__2346 (
            .O(N__11053),
            .I(N__11047));
    CascadeMux I__2345 (
            .O(N__11050),
            .I(N__11044));
    CascadeMux I__2344 (
            .O(N__11047),
            .I(N__11041));
    CascadeBuf I__2343 (
            .O(N__11044),
            .I(N__11038));
    InMux I__2342 (
            .O(N__11041),
            .I(N__11035));
    CascadeMux I__2341 (
            .O(N__11038),
            .I(N__11032));
    LocalMux I__2340 (
            .O(N__11035),
            .I(N__11029));
    InMux I__2339 (
            .O(N__11032),
            .I(N__11026));
    Span4Mux_h I__2338 (
            .O(N__11029),
            .I(N__11023));
    LocalMux I__2337 (
            .O(N__11026),
            .I(N__11019));
    Span4Mux_h I__2336 (
            .O(N__11023),
            .I(N__11015));
    InMux I__2335 (
            .O(N__11022),
            .I(N__11011));
    Span12Mux_s9_h I__2334 (
            .O(N__11019),
            .I(N__11007));
    InMux I__2333 (
            .O(N__11018),
            .I(N__11004));
    Sp12to4 I__2332 (
            .O(N__11015),
            .I(N__11001));
    InMux I__2331 (
            .O(N__11014),
            .I(N__10998));
    LocalMux I__2330 (
            .O(N__11011),
            .I(N__10995));
    InMux I__2329 (
            .O(N__11010),
            .I(N__10992));
    Span12Mux_v I__2328 (
            .O(N__11007),
            .I(N__10989));
    LocalMux I__2327 (
            .O(N__11004),
            .I(N__10984));
    Span12Mux_s10_v I__2326 (
            .O(N__11001),
            .I(N__10984));
    LocalMux I__2325 (
            .O(N__10998),
            .I(M_this_vga_signals_address_4));
    Odrv4 I__2324 (
            .O(N__10995),
            .I(M_this_vga_signals_address_4));
    LocalMux I__2323 (
            .O(N__10992),
            .I(M_this_vga_signals_address_4));
    Odrv12 I__2322 (
            .O(N__10989),
            .I(M_this_vga_signals_address_4));
    Odrv12 I__2321 (
            .O(N__10984),
            .I(M_this_vga_signals_address_4));
    CascadeMux I__2320 (
            .O(N__10973),
            .I(N__10970));
    InMux I__2319 (
            .O(N__10970),
            .I(N__10967));
    LocalMux I__2318 (
            .O(N__10967),
            .I(N__10964));
    Span4Mux_h I__2317 (
            .O(N__10964),
            .I(N__10957));
    InMux I__2316 (
            .O(N__10963),
            .I(N__10954));
    InMux I__2315 (
            .O(N__10962),
            .I(N__10949));
    InMux I__2314 (
            .O(N__10961),
            .I(N__10949));
    InMux I__2313 (
            .O(N__10960),
            .I(N__10946));
    Odrv4 I__2312 (
            .O(N__10957),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2311 (
            .O(N__10954),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2310 (
            .O(N__10949),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    LocalMux I__2309 (
            .O(N__10946),
            .I(\this_vga_signals.M_vcounter_qZ0Z_7 ));
    InMux I__2308 (
            .O(N__10937),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_6 ));
    CascadeMux I__2307 (
            .O(N__10934),
            .I(N__10930));
    InMux I__2306 (
            .O(N__10933),
            .I(N__10927));
    InMux I__2305 (
            .O(N__10930),
            .I(N__10924));
    LocalMux I__2304 (
            .O(N__10927),
            .I(N__10919));
    LocalMux I__2303 (
            .O(N__10924),
            .I(N__10915));
    InMux I__2302 (
            .O(N__10923),
            .I(N__10912));
    InMux I__2301 (
            .O(N__10922),
            .I(N__10909));
    Span4Mux_v I__2300 (
            .O(N__10919),
            .I(N__10906));
    InMux I__2299 (
            .O(N__10918),
            .I(N__10903));
    Span4Mux_v I__2298 (
            .O(N__10915),
            .I(N__10898));
    LocalMux I__2297 (
            .O(N__10912),
            .I(N__10898));
    LocalMux I__2296 (
            .O(N__10909),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2295 (
            .O(N__10906),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    LocalMux I__2294 (
            .O(N__10903),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    Odrv4 I__2293 (
            .O(N__10898),
            .I(\this_vga_signals.M_vcounter_qZ0Z_8 ));
    InMux I__2292 (
            .O(N__10889),
            .I(bfn_14_19_0_));
    InMux I__2291 (
            .O(N__10886),
            .I(N__10883));
    LocalMux I__2290 (
            .O(N__10883),
            .I(N__10880));
    Odrv4 I__2289 (
            .O(N__10880),
            .I(\this_vga_signals.M_hstate_q_ns_i_i_1_0 ));
    CascadeMux I__2288 (
            .O(N__10877),
            .I(\this_vga_signals.N_76_cascade_ ));
    CascadeMux I__2287 (
            .O(N__10874),
            .I(\this_vga_signals.N_29_cascade_ ));
    InMux I__2286 (
            .O(N__10871),
            .I(N__10866));
    InMux I__2285 (
            .O(N__10870),
            .I(N__10863));
    CascadeMux I__2284 (
            .O(N__10869),
            .I(N__10859));
    LocalMux I__2283 (
            .O(N__10866),
            .I(N__10854));
    LocalMux I__2282 (
            .O(N__10863),
            .I(N__10854));
    InMux I__2281 (
            .O(N__10862),
            .I(N__10849));
    InMux I__2280 (
            .O(N__10859),
            .I(N__10849));
    Odrv4 I__2279 (
            .O(N__10854),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__2278 (
            .O(N__10849),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__2277 (
            .O(N__10844),
            .I(N__10839));
    CascadeMux I__2276 (
            .O(N__10843),
            .I(N__10835));
    InMux I__2275 (
            .O(N__10842),
            .I(N__10831));
    InMux I__2274 (
            .O(N__10839),
            .I(N__10828));
    InMux I__2273 (
            .O(N__10838),
            .I(N__10823));
    InMux I__2272 (
            .O(N__10835),
            .I(N__10823));
    InMux I__2271 (
            .O(N__10834),
            .I(N__10820));
    LocalMux I__2270 (
            .O(N__10831),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2269 (
            .O(N__10828),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2268 (
            .O(N__10823),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__2267 (
            .O(N__10820),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    InMux I__2266 (
            .O(N__10811),
            .I(N__10808));
    LocalMux I__2265 (
            .O(N__10808),
            .I(N__10805));
    Odrv4 I__2264 (
            .O(N__10805),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_CO ));
    InMux I__2263 (
            .O(N__10802),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_0 ));
    InMux I__2262 (
            .O(N__10799),
            .I(N__10794));
    InMux I__2261 (
            .O(N__10798),
            .I(N__10789));
    InMux I__2260 (
            .O(N__10797),
            .I(N__10784));
    LocalMux I__2259 (
            .O(N__10794),
            .I(N__10781));
    InMux I__2258 (
            .O(N__10793),
            .I(N__10778));
    InMux I__2257 (
            .O(N__10792),
            .I(N__10775));
    LocalMux I__2256 (
            .O(N__10789),
            .I(N__10772));
    InMux I__2255 (
            .O(N__10788),
            .I(N__10769));
    InMux I__2254 (
            .O(N__10787),
            .I(N__10766));
    LocalMux I__2253 (
            .O(N__10784),
            .I(\this_vga_signals.address_1_0 ));
    Odrv4 I__2252 (
            .O(N__10781),
            .I(\this_vga_signals.address_1_0 ));
    LocalMux I__2251 (
            .O(N__10778),
            .I(\this_vga_signals.address_1_0 ));
    LocalMux I__2250 (
            .O(N__10775),
            .I(\this_vga_signals.address_1_0 ));
    Odrv4 I__2249 (
            .O(N__10772),
            .I(\this_vga_signals.address_1_0 ));
    LocalMux I__2248 (
            .O(N__10769),
            .I(\this_vga_signals.address_1_0 ));
    LocalMux I__2247 (
            .O(N__10766),
            .I(\this_vga_signals.address_1_0 ));
    InMux I__2246 (
            .O(N__10751),
            .I(N__10748));
    LocalMux I__2245 (
            .O(N__10748),
            .I(N__10745));
    Odrv4 I__2244 (
            .O(N__10745),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_CO ));
    InMux I__2243 (
            .O(N__10742),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_1 ));
    InMux I__2242 (
            .O(N__10739),
            .I(N__10734));
    InMux I__2241 (
            .O(N__10738),
            .I(N__10731));
    InMux I__2240 (
            .O(N__10737),
            .I(N__10724));
    LocalMux I__2239 (
            .O(N__10734),
            .I(N__10719));
    LocalMux I__2238 (
            .O(N__10731),
            .I(N__10719));
    InMux I__2237 (
            .O(N__10730),
            .I(N__10714));
    InMux I__2236 (
            .O(N__10729),
            .I(N__10714));
    InMux I__2235 (
            .O(N__10728),
            .I(N__10711));
    InMux I__2234 (
            .O(N__10727),
            .I(N__10708));
    LocalMux I__2233 (
            .O(N__10724),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__2232 (
            .O(N__10719),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2231 (
            .O(N__10714),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2230 (
            .O(N__10711),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__2229 (
            .O(N__10708),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    CascadeMux I__2228 (
            .O(N__10697),
            .I(N__10694));
    InMux I__2227 (
            .O(N__10694),
            .I(N__10691));
    LocalMux I__2226 (
            .O(N__10691),
            .I(N__10688));
    Odrv4 I__2225 (
            .O(N__10688),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_CO ));
    InMux I__2224 (
            .O(N__10685),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_2 ));
    InMux I__2223 (
            .O(N__10682),
            .I(N__10677));
    InMux I__2222 (
            .O(N__10681),
            .I(N__10672));
    InMux I__2221 (
            .O(N__10680),
            .I(N__10672));
    LocalMux I__2220 (
            .O(N__10677),
            .I(N__10667));
    LocalMux I__2219 (
            .O(N__10672),
            .I(N__10663));
    InMux I__2218 (
            .O(N__10671),
            .I(N__10660));
    InMux I__2217 (
            .O(N__10670),
            .I(N__10657));
    Span4Mux_v I__2216 (
            .O(N__10667),
            .I(N__10654));
    InMux I__2215 (
            .O(N__10666),
            .I(N__10651));
    Odrv4 I__2214 (
            .O(N__10663),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2213 (
            .O(N__10660),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2212 (
            .O(N__10657),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2211 (
            .O(N__10654),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2210 (
            .O(N__10651),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    InMux I__2209 (
            .O(N__10640),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_3 ));
    InMux I__2208 (
            .O(N__10637),
            .I(N__10633));
    CascadeMux I__2207 (
            .O(N__10636),
            .I(N__10627));
    LocalMux I__2206 (
            .O(N__10633),
            .I(N__10624));
    InMux I__2205 (
            .O(N__10632),
            .I(N__10621));
    InMux I__2204 (
            .O(N__10631),
            .I(N__10616));
    InMux I__2203 (
            .O(N__10630),
            .I(N__10616));
    InMux I__2202 (
            .O(N__10627),
            .I(N__10613));
    Odrv4 I__2201 (
            .O(N__10624),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2200 (
            .O(N__10621),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2199 (
            .O(N__10616),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2198 (
            .O(N__10613),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__2197 (
            .O(N__10604),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_4 ));
    CascadeMux I__2196 (
            .O(N__10601),
            .I(N__10598));
    InMux I__2195 (
            .O(N__10598),
            .I(N__10595));
    LocalMux I__2194 (
            .O(N__10595),
            .I(N__10592));
    Span4Mux_h I__2193 (
            .O(N__10592),
            .I(N__10585));
    InMux I__2192 (
            .O(N__10591),
            .I(N__10582));
    InMux I__2191 (
            .O(N__10590),
            .I(N__10577));
    InMux I__2190 (
            .O(N__10589),
            .I(N__10577));
    InMux I__2189 (
            .O(N__10588),
            .I(N__10574));
    Odrv4 I__2188 (
            .O(N__10585),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2187 (
            .O(N__10582),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2186 (
            .O(N__10577),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2185 (
            .O(N__10574),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    InMux I__2184 (
            .O(N__10565),
            .I(\this_vga_signals.un1_M_vcounter_q_6_cry_5 ));
    InMux I__2183 (
            .O(N__10562),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__2182 (
            .O(N__10559),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__2181 (
            .O(N__10556),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__2180 (
            .O(N__10553),
            .I(bfn_14_16_0_));
    InMux I__2179 (
            .O(N__10550),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_9 ));
    InMux I__2178 (
            .O(N__10547),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_10 ));
    CascadeMux I__2177 (
            .O(N__10544),
            .I(\this_vga_signals.N_68_cascade_ ));
    InMux I__2176 (
            .O(N__10541),
            .I(N__10536));
    InMux I__2175 (
            .O(N__10540),
            .I(N__10531));
    InMux I__2174 (
            .O(N__10539),
            .I(N__10531));
    LocalMux I__2173 (
            .O(N__10536),
            .I(\this_vga_signals.m27_0_a2_1_4 ));
    LocalMux I__2172 (
            .O(N__10531),
            .I(\this_vga_signals.m27_0_a2_1_4 ));
    InMux I__2171 (
            .O(N__10526),
            .I(N__10523));
    LocalMux I__2170 (
            .O(N__10523),
            .I(\this_vga_signals.M_vcounter_q_0_i_a2_0_0 ));
    CascadeMux I__2169 (
            .O(N__10520),
            .I(N__10516));
    InMux I__2168 (
            .O(N__10519),
            .I(N__10510));
    InMux I__2167 (
            .O(N__10516),
            .I(N__10510));
    InMux I__2166 (
            .O(N__10515),
            .I(N__10507));
    LocalMux I__2165 (
            .O(N__10510),
            .I(N__10502));
    LocalMux I__2164 (
            .O(N__10507),
            .I(N__10502));
    Span12Mux_s5_h I__2163 (
            .O(N__10502),
            .I(N__10493));
    InMux I__2162 (
            .O(N__10501),
            .I(N__10484));
    InMux I__2161 (
            .O(N__10500),
            .I(N__10484));
    InMux I__2160 (
            .O(N__10499),
            .I(N__10484));
    InMux I__2159 (
            .O(N__10498),
            .I(N__10484));
    InMux I__2158 (
            .O(N__10497),
            .I(N__10479));
    InMux I__2157 (
            .O(N__10496),
            .I(N__10479));
    Odrv12 I__2156 (
            .O(N__10493),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    LocalMux I__2155 (
            .O(N__10484),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    LocalMux I__2154 (
            .O(N__10479),
            .I(\this_vga_signals.M_vstate_qZ0Z_0 ));
    InMux I__2153 (
            .O(N__10472),
            .I(N__10466));
    InMux I__2152 (
            .O(N__10471),
            .I(N__10466));
    LocalMux I__2151 (
            .O(N__10466),
            .I(N__10458));
    InMux I__2150 (
            .O(N__10465),
            .I(N__10455));
    CascadeMux I__2149 (
            .O(N__10464),
            .I(N__10450));
    CascadeMux I__2148 (
            .O(N__10463),
            .I(N__10447));
    CascadeMux I__2147 (
            .O(N__10462),
            .I(N__10444));
    CascadeMux I__2146 (
            .O(N__10461),
            .I(N__10440));
    Sp12to4 I__2145 (
            .O(N__10458),
            .I(N__10435));
    LocalMux I__2144 (
            .O(N__10455),
            .I(N__10435));
    InMux I__2143 (
            .O(N__10454),
            .I(N__10428));
    InMux I__2142 (
            .O(N__10453),
            .I(N__10428));
    InMux I__2141 (
            .O(N__10450),
            .I(N__10428));
    InMux I__2140 (
            .O(N__10447),
            .I(N__10423));
    InMux I__2139 (
            .O(N__10444),
            .I(N__10423));
    InMux I__2138 (
            .O(N__10443),
            .I(N__10418));
    InMux I__2137 (
            .O(N__10440),
            .I(N__10418));
    Odrv12 I__2136 (
            .O(N__10435),
            .I(\this_vga_signals.M_vstate_qZ0Z_1 ));
    LocalMux I__2135 (
            .O(N__10428),
            .I(\this_vga_signals.M_vstate_qZ0Z_1 ));
    LocalMux I__2134 (
            .O(N__10423),
            .I(\this_vga_signals.M_vstate_qZ0Z_1 ));
    LocalMux I__2133 (
            .O(N__10418),
            .I(\this_vga_signals.M_vstate_qZ0Z_1 ));
    InMux I__2132 (
            .O(N__10409),
            .I(N__10406));
    LocalMux I__2131 (
            .O(N__10406),
            .I(\this_vga_signals.m24_0_0 ));
    InMux I__2130 (
            .O(N__10403),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__2129 (
            .O(N__10400),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__2128 (
            .O(N__10397),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__2127 (
            .O(N__10394),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__2126 (
            .O(N__10391),
            .I(\this_vga_signals.address_1_0_cry_2 ));
    CascadeMux I__2125 (
            .O(N__10388),
            .I(N__10385));
    InMux I__2124 (
            .O(N__10385),
            .I(N__10382));
    LocalMux I__2123 (
            .O(N__10382),
            .I(N__10379));
    Odrv4 I__2122 (
            .O(N__10379),
            .I(\this_vga_signals.address_1_0_4 ));
    InMux I__2121 (
            .O(N__10376),
            .I(\this_vga_signals.address_1_0_cry_3 ));
    CascadeMux I__2120 (
            .O(N__10373),
            .I(N__10370));
    InMux I__2119 (
            .O(N__10370),
            .I(N__10367));
    LocalMux I__2118 (
            .O(N__10367),
            .I(N__10364));
    Odrv4 I__2117 (
            .O(N__10364),
            .I(\this_vga_signals.address_1_0_5 ));
    InMux I__2116 (
            .O(N__10361),
            .I(\this_vga_signals.address_1_0_cry_4 ));
    InMux I__2115 (
            .O(N__10358),
            .I(N__10355));
    LocalMux I__2114 (
            .O(N__10355),
            .I(N__10352));
    Odrv4 I__2113 (
            .O(N__10352),
            .I(\this_vga_signals.address_1_0_6 ));
    InMux I__2112 (
            .O(N__10349),
            .I(\this_vga_signals.address_1_0_cry_5 ));
    InMux I__2111 (
            .O(N__10346),
            .I(N__10343));
    LocalMux I__2110 (
            .O(N__10343),
            .I(N__10340));
    Odrv4 I__2109 (
            .O(N__10340),
            .I(\this_vga_signals.address_1_0_7 ));
    InMux I__2108 (
            .O(N__10337),
            .I(\this_vga_signals.address_1_0_cry_6 ));
    InMux I__2107 (
            .O(N__10334),
            .I(bfn_13_18_0_));
    InMux I__2106 (
            .O(N__10331),
            .I(N__10328));
    LocalMux I__2105 (
            .O(N__10328),
            .I(N__10325));
    Odrv4 I__2104 (
            .O(N__10325),
            .I(\this_vga_signals.address_1_0_8_THRU_CO ));
    InMux I__2103 (
            .O(N__10322),
            .I(N__10319));
    LocalMux I__2102 (
            .O(N__10319),
            .I(\this_vga_signals.m27_0_o2_0_3 ));
    InMux I__2101 (
            .O(N__10316),
            .I(N__10313));
    LocalMux I__2100 (
            .O(N__10313),
            .I(\this_vga_signals.N_36 ));
    InMux I__2099 (
            .O(N__10310),
            .I(N__10304));
    InMux I__2098 (
            .O(N__10309),
            .I(N__10304));
    LocalMux I__2097 (
            .O(N__10304),
            .I(\this_vga_signals.m27_0_a2_1_5 ));
    CascadeMux I__2096 (
            .O(N__10301),
            .I(\this_vga_signals.m27_0_a2_1_5_cascade_ ));
    InMux I__2095 (
            .O(N__10298),
            .I(\this_vga_signals.address_1_cry_4 ));
    InMux I__2094 (
            .O(N__10295),
            .I(N__10290));
    InMux I__2093 (
            .O(N__10294),
            .I(N__10287));
    InMux I__2092 (
            .O(N__10293),
            .I(N__10284));
    LocalMux I__2091 (
            .O(N__10290),
            .I(N__10274));
    LocalMux I__2090 (
            .O(N__10287),
            .I(N__10274));
    LocalMux I__2089 (
            .O(N__10284),
            .I(N__10274));
    InMux I__2088 (
            .O(N__10283),
            .I(N__10270));
    InMux I__2087 (
            .O(N__10282),
            .I(N__10267));
    InMux I__2086 (
            .O(N__10281),
            .I(N__10264));
    Span4Mux_v I__2085 (
            .O(N__10274),
            .I(N__10261));
    InMux I__2084 (
            .O(N__10273),
            .I(N__10258));
    LocalMux I__2083 (
            .O(N__10270),
            .I(N__10251));
    LocalMux I__2082 (
            .O(N__10267),
            .I(N__10251));
    LocalMux I__2081 (
            .O(N__10264),
            .I(N__10251));
    Sp12to4 I__2080 (
            .O(N__10261),
            .I(N__10246));
    LocalMux I__2079 (
            .O(N__10258),
            .I(N__10246));
    Span4Mux_v I__2078 (
            .O(N__10251),
            .I(N__10243));
    Odrv12 I__2077 (
            .O(N__10246),
            .I(\this_vram.mem_radregZ0Z_13 ));
    Odrv4 I__2076 (
            .O(N__10243),
            .I(\this_vram.mem_radregZ0Z_13 ));
    InMux I__2075 (
            .O(N__10238),
            .I(\this_vga_signals.address_1_cry_5 ));
    InMux I__2074 (
            .O(N__10235),
            .I(\this_vga_signals.address_1_cry_6 ));
    InMux I__2073 (
            .O(N__10232),
            .I(N__10225));
    InMux I__2072 (
            .O(N__10231),
            .I(N__10225));
    InMux I__2071 (
            .O(N__10230),
            .I(N__10222));
    LocalMux I__2070 (
            .O(N__10225),
            .I(N__10217));
    LocalMux I__2069 (
            .O(N__10222),
            .I(N__10217));
    Span4Mux_v I__2068 (
            .O(N__10217),
            .I(N__10211));
    InMux I__2067 (
            .O(N__10216),
            .I(N__10208));
    InMux I__2066 (
            .O(N__10215),
            .I(N__10203));
    InMux I__2065 (
            .O(N__10214),
            .I(N__10203));
    Span4Mux_h I__2064 (
            .O(N__10211),
            .I(N__10199));
    LocalMux I__2063 (
            .O(N__10208),
            .I(N__10194));
    LocalMux I__2062 (
            .O(N__10203),
            .I(N__10194));
    InMux I__2061 (
            .O(N__10202),
            .I(N__10191));
    Span4Mux_v I__2060 (
            .O(N__10199),
            .I(N__10188));
    Span4Mux_v I__2059 (
            .O(N__10194),
            .I(N__10185));
    LocalMux I__2058 (
            .O(N__10191),
            .I(N__10182));
    Odrv4 I__2057 (
            .O(N__10188),
            .I(\this_vram.mem_radregZ0Z_14 ));
    Odrv4 I__2056 (
            .O(N__10185),
            .I(\this_vram.mem_radregZ0Z_14 ));
    Odrv12 I__2055 (
            .O(N__10182),
            .I(\this_vram.mem_radregZ0Z_14 ));
    CascadeMux I__2054 (
            .O(N__10175),
            .I(N__10172));
    CascadeBuf I__2053 (
            .O(N__10172),
            .I(N__10169));
    CascadeMux I__2052 (
            .O(N__10169),
            .I(N__10166));
    CascadeBuf I__2051 (
            .O(N__10166),
            .I(N__10163));
    CascadeMux I__2050 (
            .O(N__10163),
            .I(N__10159));
    CascadeMux I__2049 (
            .O(N__10162),
            .I(N__10156));
    CascadeBuf I__2048 (
            .O(N__10159),
            .I(N__10153));
    CascadeBuf I__2047 (
            .O(N__10156),
            .I(N__10150));
    CascadeMux I__2046 (
            .O(N__10153),
            .I(N__10147));
    CascadeMux I__2045 (
            .O(N__10150),
            .I(N__10144));
    CascadeBuf I__2044 (
            .O(N__10147),
            .I(N__10141));
    CascadeBuf I__2043 (
            .O(N__10144),
            .I(N__10138));
    CascadeMux I__2042 (
            .O(N__10141),
            .I(N__10135));
    CascadeMux I__2041 (
            .O(N__10138),
            .I(N__10132));
    CascadeBuf I__2040 (
            .O(N__10135),
            .I(N__10129));
    CascadeBuf I__2039 (
            .O(N__10132),
            .I(N__10126));
    CascadeMux I__2038 (
            .O(N__10129),
            .I(N__10123));
    CascadeMux I__2037 (
            .O(N__10126),
            .I(N__10120));
    CascadeBuf I__2036 (
            .O(N__10123),
            .I(N__10117));
    CascadeBuf I__2035 (
            .O(N__10120),
            .I(N__10114));
    CascadeMux I__2034 (
            .O(N__10117),
            .I(N__10111));
    CascadeMux I__2033 (
            .O(N__10114),
            .I(N__10108));
    CascadeBuf I__2032 (
            .O(N__10111),
            .I(N__10105));
    CascadeBuf I__2031 (
            .O(N__10108),
            .I(N__10102));
    CascadeMux I__2030 (
            .O(N__10105),
            .I(N__10099));
    CascadeMux I__2029 (
            .O(N__10102),
            .I(N__10096));
    CascadeBuf I__2028 (
            .O(N__10099),
            .I(N__10093));
    CascadeBuf I__2027 (
            .O(N__10096),
            .I(N__10090));
    CascadeMux I__2026 (
            .O(N__10093),
            .I(N__10087));
    CascadeMux I__2025 (
            .O(N__10090),
            .I(N__10084));
    CascadeBuf I__2024 (
            .O(N__10087),
            .I(N__10081));
    CascadeBuf I__2023 (
            .O(N__10084),
            .I(N__10078));
    CascadeMux I__2022 (
            .O(N__10081),
            .I(N__10075));
    CascadeMux I__2021 (
            .O(N__10078),
            .I(N__10072));
    CascadeBuf I__2020 (
            .O(N__10075),
            .I(N__10069));
    CascadeBuf I__2019 (
            .O(N__10072),
            .I(N__10066));
    CascadeMux I__2018 (
            .O(N__10069),
            .I(N__10063));
    CascadeMux I__2017 (
            .O(N__10066),
            .I(N__10060));
    CascadeBuf I__2016 (
            .O(N__10063),
            .I(N__10057));
    CascadeBuf I__2015 (
            .O(N__10060),
            .I(N__10054));
    CascadeMux I__2014 (
            .O(N__10057),
            .I(N__10051));
    CascadeMux I__2013 (
            .O(N__10054),
            .I(N__10048));
    CascadeBuf I__2012 (
            .O(N__10051),
            .I(N__10045));
    CascadeBuf I__2011 (
            .O(N__10048),
            .I(N__10042));
    CascadeMux I__2010 (
            .O(N__10045),
            .I(N__10039));
    CascadeMux I__2009 (
            .O(N__10042),
            .I(N__10036));
    CascadeBuf I__2008 (
            .O(N__10039),
            .I(N__10033));
    CascadeBuf I__2007 (
            .O(N__10036),
            .I(N__10030));
    CascadeMux I__2006 (
            .O(N__10033),
            .I(N__10027));
    CascadeMux I__2005 (
            .O(N__10030),
            .I(N__10024));
    CascadeBuf I__2004 (
            .O(N__10027),
            .I(N__10021));
    CascadeBuf I__2003 (
            .O(N__10024),
            .I(N__10018));
    CascadeMux I__2002 (
            .O(N__10021),
            .I(N__10015));
    CascadeMux I__2001 (
            .O(N__10018),
            .I(N__10012));
    CascadeBuf I__2000 (
            .O(N__10015),
            .I(N__10009));
    CascadeBuf I__1999 (
            .O(N__10012),
            .I(N__10006));
    CascadeMux I__1998 (
            .O(N__10009),
            .I(N__10003));
    CascadeMux I__1997 (
            .O(N__10006),
            .I(N__10000));
    InMux I__1996 (
            .O(N__10003),
            .I(N__9997));
    InMux I__1995 (
            .O(N__10000),
            .I(N__9994));
    LocalMux I__1994 (
            .O(N__9997),
            .I(N__9991));
    LocalMux I__1993 (
            .O(N__9994),
            .I(N__9988));
    Sp12to4 I__1992 (
            .O(N__9991),
            .I(N__9985));
    Span12Mux_v I__1991 (
            .O(N__9988),
            .I(N__9982));
    Span12Mux_s3_v I__1990 (
            .O(N__9985),
            .I(N__9979));
    Span12Mux_h I__1989 (
            .O(N__9982),
            .I(N__9976));
    Span12Mux_v I__1988 (
            .O(N__9979),
            .I(N__9973));
    Odrv12 I__1987 (
            .O(N__9976),
            .I(M_this_vga_signals_address_5));
    Odrv12 I__1986 (
            .O(N__9973),
            .I(M_this_vga_signals_address_5));
    CascadeMux I__1985 (
            .O(N__9968),
            .I(N__9965));
    CascadeBuf I__1984 (
            .O(N__9965),
            .I(N__9962));
    CascadeMux I__1983 (
            .O(N__9962),
            .I(N__9959));
    CascadeBuf I__1982 (
            .O(N__9959),
            .I(N__9956));
    CascadeMux I__1981 (
            .O(N__9956),
            .I(N__9952));
    CascadeMux I__1980 (
            .O(N__9955),
            .I(N__9949));
    CascadeBuf I__1979 (
            .O(N__9952),
            .I(N__9946));
    CascadeBuf I__1978 (
            .O(N__9949),
            .I(N__9943));
    CascadeMux I__1977 (
            .O(N__9946),
            .I(N__9940));
    CascadeMux I__1976 (
            .O(N__9943),
            .I(N__9937));
    CascadeBuf I__1975 (
            .O(N__9940),
            .I(N__9934));
    CascadeBuf I__1974 (
            .O(N__9937),
            .I(N__9931));
    CascadeMux I__1973 (
            .O(N__9934),
            .I(N__9928));
    CascadeMux I__1972 (
            .O(N__9931),
            .I(N__9925));
    CascadeBuf I__1971 (
            .O(N__9928),
            .I(N__9922));
    CascadeBuf I__1970 (
            .O(N__9925),
            .I(N__9919));
    CascadeMux I__1969 (
            .O(N__9922),
            .I(N__9916));
    CascadeMux I__1968 (
            .O(N__9919),
            .I(N__9913));
    CascadeBuf I__1967 (
            .O(N__9916),
            .I(N__9910));
    CascadeBuf I__1966 (
            .O(N__9913),
            .I(N__9907));
    CascadeMux I__1965 (
            .O(N__9910),
            .I(N__9904));
    CascadeMux I__1964 (
            .O(N__9907),
            .I(N__9901));
    CascadeBuf I__1963 (
            .O(N__9904),
            .I(N__9898));
    CascadeBuf I__1962 (
            .O(N__9901),
            .I(N__9895));
    CascadeMux I__1961 (
            .O(N__9898),
            .I(N__9892));
    CascadeMux I__1960 (
            .O(N__9895),
            .I(N__9889));
    CascadeBuf I__1959 (
            .O(N__9892),
            .I(N__9886));
    CascadeBuf I__1958 (
            .O(N__9889),
            .I(N__9883));
    CascadeMux I__1957 (
            .O(N__9886),
            .I(N__9880));
    CascadeMux I__1956 (
            .O(N__9883),
            .I(N__9877));
    CascadeBuf I__1955 (
            .O(N__9880),
            .I(N__9874));
    CascadeBuf I__1954 (
            .O(N__9877),
            .I(N__9871));
    CascadeMux I__1953 (
            .O(N__9874),
            .I(N__9868));
    CascadeMux I__1952 (
            .O(N__9871),
            .I(N__9865));
    CascadeBuf I__1951 (
            .O(N__9868),
            .I(N__9862));
    CascadeBuf I__1950 (
            .O(N__9865),
            .I(N__9859));
    CascadeMux I__1949 (
            .O(N__9862),
            .I(N__9856));
    CascadeMux I__1948 (
            .O(N__9859),
            .I(N__9853));
    CascadeBuf I__1947 (
            .O(N__9856),
            .I(N__9850));
    CascadeBuf I__1946 (
            .O(N__9853),
            .I(N__9847));
    CascadeMux I__1945 (
            .O(N__9850),
            .I(N__9844));
    CascadeMux I__1944 (
            .O(N__9847),
            .I(N__9841));
    CascadeBuf I__1943 (
            .O(N__9844),
            .I(N__9838));
    CascadeBuf I__1942 (
            .O(N__9841),
            .I(N__9835));
    CascadeMux I__1941 (
            .O(N__9838),
            .I(N__9832));
    CascadeMux I__1940 (
            .O(N__9835),
            .I(N__9829));
    CascadeBuf I__1939 (
            .O(N__9832),
            .I(N__9826));
    CascadeBuf I__1938 (
            .O(N__9829),
            .I(N__9823));
    CascadeMux I__1937 (
            .O(N__9826),
            .I(N__9820));
    CascadeMux I__1936 (
            .O(N__9823),
            .I(N__9817));
    CascadeBuf I__1935 (
            .O(N__9820),
            .I(N__9814));
    CascadeBuf I__1934 (
            .O(N__9817),
            .I(N__9811));
    CascadeMux I__1933 (
            .O(N__9814),
            .I(N__9808));
    CascadeMux I__1932 (
            .O(N__9811),
            .I(N__9805));
    CascadeBuf I__1931 (
            .O(N__9808),
            .I(N__9802));
    CascadeBuf I__1930 (
            .O(N__9805),
            .I(N__9799));
    CascadeMux I__1929 (
            .O(N__9802),
            .I(N__9796));
    CascadeMux I__1928 (
            .O(N__9799),
            .I(N__9793));
    InMux I__1927 (
            .O(N__9796),
            .I(N__9790));
    InMux I__1926 (
            .O(N__9793),
            .I(N__9787));
    LocalMux I__1925 (
            .O(N__9790),
            .I(N__9784));
    LocalMux I__1924 (
            .O(N__9787),
            .I(N__9781));
    Span4Mux_s2_v I__1923 (
            .O(N__9784),
            .I(N__9778));
    Span12Mux_v I__1922 (
            .O(N__9781),
            .I(N__9775));
    Sp12to4 I__1921 (
            .O(N__9778),
            .I(N__9772));
    Span12Mux_h I__1920 (
            .O(N__9775),
            .I(N__9769));
    Span12Mux_v I__1919 (
            .O(N__9772),
            .I(N__9766));
    Odrv12 I__1918 (
            .O(N__9769),
            .I(M_this_vga_signals_address_6));
    Odrv12 I__1917 (
            .O(N__9766),
            .I(M_this_vga_signals_address_6));
    InMux I__1916 (
            .O(N__9761),
            .I(\this_vga_signals.address_1_0_cry_0 ));
    CascadeMux I__1915 (
            .O(N__9758),
            .I(N__9755));
    InMux I__1914 (
            .O(N__9755),
            .I(N__9752));
    LocalMux I__1913 (
            .O(N__9752),
            .I(N__9749));
    Odrv4 I__1912 (
            .O(N__9749),
            .I(\this_vga_signals.address_1 ));
    InMux I__1911 (
            .O(N__9746),
            .I(\this_vga_signals.address_1_0_cry_1 ));
    CascadeMux I__1910 (
            .O(N__9743),
            .I(N__9740));
    InMux I__1909 (
            .O(N__9740),
            .I(N__9737));
    LocalMux I__1908 (
            .O(N__9737),
            .I(N__9734));
    Odrv4 I__1907 (
            .O(N__9734),
            .I(\this_vga_signals.address_1_0_3 ));
    InMux I__1906 (
            .O(N__9731),
            .I(N__9725));
    InMux I__1905 (
            .O(N__9730),
            .I(N__9725));
    LocalMux I__1904 (
            .O(N__9725),
            .I(\this_vga_signals.m27_0_o2_1 ));
    CascadeMux I__1903 (
            .O(N__9722),
            .I(\this_vga_signals.m27_0_0_cascade_ ));
    CascadeMux I__1902 (
            .O(N__9719),
            .I(\this_vga_signals.i9_mux_cascade_ ));
    InMux I__1901 (
            .O(N__9716),
            .I(N__9710));
    InMux I__1900 (
            .O(N__9715),
            .I(N__9710));
    LocalMux I__1899 (
            .O(N__9710),
            .I(\this_vga_signals.N_40 ));
    CascadeMux I__1898 (
            .O(N__9707),
            .I(N__9704));
    CascadeBuf I__1897 (
            .O(N__9704),
            .I(N__9701));
    CascadeMux I__1896 (
            .O(N__9701),
            .I(N__9698));
    CascadeBuf I__1895 (
            .O(N__9698),
            .I(N__9695));
    CascadeMux I__1894 (
            .O(N__9695),
            .I(N__9691));
    CascadeMux I__1893 (
            .O(N__9694),
            .I(N__9688));
    CascadeBuf I__1892 (
            .O(N__9691),
            .I(N__9685));
    CascadeBuf I__1891 (
            .O(N__9688),
            .I(N__9682));
    CascadeMux I__1890 (
            .O(N__9685),
            .I(N__9679));
    CascadeMux I__1889 (
            .O(N__9682),
            .I(N__9676));
    CascadeBuf I__1888 (
            .O(N__9679),
            .I(N__9673));
    CascadeBuf I__1887 (
            .O(N__9676),
            .I(N__9670));
    CascadeMux I__1886 (
            .O(N__9673),
            .I(N__9667));
    CascadeMux I__1885 (
            .O(N__9670),
            .I(N__9664));
    CascadeBuf I__1884 (
            .O(N__9667),
            .I(N__9661));
    CascadeBuf I__1883 (
            .O(N__9664),
            .I(N__9658));
    CascadeMux I__1882 (
            .O(N__9661),
            .I(N__9655));
    CascadeMux I__1881 (
            .O(N__9658),
            .I(N__9652));
    CascadeBuf I__1880 (
            .O(N__9655),
            .I(N__9649));
    CascadeBuf I__1879 (
            .O(N__9652),
            .I(N__9646));
    CascadeMux I__1878 (
            .O(N__9649),
            .I(N__9643));
    CascadeMux I__1877 (
            .O(N__9646),
            .I(N__9640));
    CascadeBuf I__1876 (
            .O(N__9643),
            .I(N__9637));
    CascadeBuf I__1875 (
            .O(N__9640),
            .I(N__9634));
    CascadeMux I__1874 (
            .O(N__9637),
            .I(N__9631));
    CascadeMux I__1873 (
            .O(N__9634),
            .I(N__9628));
    CascadeBuf I__1872 (
            .O(N__9631),
            .I(N__9625));
    CascadeBuf I__1871 (
            .O(N__9628),
            .I(N__9622));
    CascadeMux I__1870 (
            .O(N__9625),
            .I(N__9619));
    CascadeMux I__1869 (
            .O(N__9622),
            .I(N__9616));
    CascadeBuf I__1868 (
            .O(N__9619),
            .I(N__9613));
    CascadeBuf I__1867 (
            .O(N__9616),
            .I(N__9610));
    CascadeMux I__1866 (
            .O(N__9613),
            .I(N__9607));
    CascadeMux I__1865 (
            .O(N__9610),
            .I(N__9604));
    CascadeBuf I__1864 (
            .O(N__9607),
            .I(N__9601));
    CascadeBuf I__1863 (
            .O(N__9604),
            .I(N__9598));
    CascadeMux I__1862 (
            .O(N__9601),
            .I(N__9595));
    CascadeMux I__1861 (
            .O(N__9598),
            .I(N__9592));
    CascadeBuf I__1860 (
            .O(N__9595),
            .I(N__9589));
    CascadeBuf I__1859 (
            .O(N__9592),
            .I(N__9586));
    CascadeMux I__1858 (
            .O(N__9589),
            .I(N__9583));
    CascadeMux I__1857 (
            .O(N__9586),
            .I(N__9580));
    CascadeBuf I__1856 (
            .O(N__9583),
            .I(N__9577));
    CascadeBuf I__1855 (
            .O(N__9580),
            .I(N__9574));
    CascadeMux I__1854 (
            .O(N__9577),
            .I(N__9571));
    CascadeMux I__1853 (
            .O(N__9574),
            .I(N__9568));
    CascadeBuf I__1852 (
            .O(N__9571),
            .I(N__9565));
    CascadeBuf I__1851 (
            .O(N__9568),
            .I(N__9562));
    CascadeMux I__1850 (
            .O(N__9565),
            .I(N__9559));
    CascadeMux I__1849 (
            .O(N__9562),
            .I(N__9556));
    CascadeBuf I__1848 (
            .O(N__9559),
            .I(N__9553));
    CascadeBuf I__1847 (
            .O(N__9556),
            .I(N__9550));
    CascadeMux I__1846 (
            .O(N__9553),
            .I(N__9547));
    CascadeMux I__1845 (
            .O(N__9550),
            .I(N__9544));
    CascadeBuf I__1844 (
            .O(N__9547),
            .I(N__9541));
    CascadeBuf I__1843 (
            .O(N__9544),
            .I(N__9538));
    CascadeMux I__1842 (
            .O(N__9541),
            .I(N__9535));
    CascadeMux I__1841 (
            .O(N__9538),
            .I(N__9532));
    InMux I__1840 (
            .O(N__9535),
            .I(N__9529));
    InMux I__1839 (
            .O(N__9532),
            .I(N__9526));
    LocalMux I__1838 (
            .O(N__9529),
            .I(N__9523));
    LocalMux I__1837 (
            .O(N__9526),
            .I(N__9520));
    Sp12to4 I__1836 (
            .O(N__9523),
            .I(N__9517));
    Span12Mux_s9_v I__1835 (
            .O(N__9520),
            .I(N__9514));
    Span12Mux_s5_v I__1834 (
            .O(N__9517),
            .I(N__9511));
    Span12Mux_h I__1833 (
            .O(N__9514),
            .I(N__9508));
    Span12Mux_v I__1832 (
            .O(N__9511),
            .I(N__9505));
    Odrv12 I__1831 (
            .O(N__9508),
            .I(M_this_vga_signals_address_7));
    Odrv12 I__1830 (
            .O(N__9505),
            .I(M_this_vga_signals_address_7));
    CascadeMux I__1829 (
            .O(N__9500),
            .I(N__9497));
    CascadeBuf I__1828 (
            .O(N__9497),
            .I(N__9494));
    CascadeMux I__1827 (
            .O(N__9494),
            .I(N__9491));
    CascadeBuf I__1826 (
            .O(N__9491),
            .I(N__9488));
    CascadeMux I__1825 (
            .O(N__9488),
            .I(N__9484));
    CascadeMux I__1824 (
            .O(N__9487),
            .I(N__9481));
    CascadeBuf I__1823 (
            .O(N__9484),
            .I(N__9478));
    CascadeBuf I__1822 (
            .O(N__9481),
            .I(N__9475));
    CascadeMux I__1821 (
            .O(N__9478),
            .I(N__9472));
    CascadeMux I__1820 (
            .O(N__9475),
            .I(N__9469));
    CascadeBuf I__1819 (
            .O(N__9472),
            .I(N__9466));
    CascadeBuf I__1818 (
            .O(N__9469),
            .I(N__9463));
    CascadeMux I__1817 (
            .O(N__9466),
            .I(N__9460));
    CascadeMux I__1816 (
            .O(N__9463),
            .I(N__9457));
    CascadeBuf I__1815 (
            .O(N__9460),
            .I(N__9454));
    CascadeBuf I__1814 (
            .O(N__9457),
            .I(N__9451));
    CascadeMux I__1813 (
            .O(N__9454),
            .I(N__9448));
    CascadeMux I__1812 (
            .O(N__9451),
            .I(N__9445));
    CascadeBuf I__1811 (
            .O(N__9448),
            .I(N__9442));
    CascadeBuf I__1810 (
            .O(N__9445),
            .I(N__9439));
    CascadeMux I__1809 (
            .O(N__9442),
            .I(N__9436));
    CascadeMux I__1808 (
            .O(N__9439),
            .I(N__9433));
    CascadeBuf I__1807 (
            .O(N__9436),
            .I(N__9430));
    CascadeBuf I__1806 (
            .O(N__9433),
            .I(N__9427));
    CascadeMux I__1805 (
            .O(N__9430),
            .I(N__9424));
    CascadeMux I__1804 (
            .O(N__9427),
            .I(N__9421));
    CascadeBuf I__1803 (
            .O(N__9424),
            .I(N__9418));
    CascadeBuf I__1802 (
            .O(N__9421),
            .I(N__9415));
    CascadeMux I__1801 (
            .O(N__9418),
            .I(N__9412));
    CascadeMux I__1800 (
            .O(N__9415),
            .I(N__9409));
    CascadeBuf I__1799 (
            .O(N__9412),
            .I(N__9406));
    CascadeBuf I__1798 (
            .O(N__9409),
            .I(N__9403));
    CascadeMux I__1797 (
            .O(N__9406),
            .I(N__9400));
    CascadeMux I__1796 (
            .O(N__9403),
            .I(N__9397));
    CascadeBuf I__1795 (
            .O(N__9400),
            .I(N__9394));
    CascadeBuf I__1794 (
            .O(N__9397),
            .I(N__9391));
    CascadeMux I__1793 (
            .O(N__9394),
            .I(N__9388));
    CascadeMux I__1792 (
            .O(N__9391),
            .I(N__9385));
    CascadeBuf I__1791 (
            .O(N__9388),
            .I(N__9382));
    CascadeBuf I__1790 (
            .O(N__9385),
            .I(N__9379));
    CascadeMux I__1789 (
            .O(N__9382),
            .I(N__9376));
    CascadeMux I__1788 (
            .O(N__9379),
            .I(N__9373));
    CascadeBuf I__1787 (
            .O(N__9376),
            .I(N__9370));
    CascadeBuf I__1786 (
            .O(N__9373),
            .I(N__9367));
    CascadeMux I__1785 (
            .O(N__9370),
            .I(N__9364));
    CascadeMux I__1784 (
            .O(N__9367),
            .I(N__9361));
    CascadeBuf I__1783 (
            .O(N__9364),
            .I(N__9358));
    CascadeBuf I__1782 (
            .O(N__9361),
            .I(N__9355));
    CascadeMux I__1781 (
            .O(N__9358),
            .I(N__9352));
    CascadeMux I__1780 (
            .O(N__9355),
            .I(N__9349));
    CascadeBuf I__1779 (
            .O(N__9352),
            .I(N__9346));
    CascadeBuf I__1778 (
            .O(N__9349),
            .I(N__9343));
    CascadeMux I__1777 (
            .O(N__9346),
            .I(N__9340));
    CascadeMux I__1776 (
            .O(N__9343),
            .I(N__9337));
    CascadeBuf I__1775 (
            .O(N__9340),
            .I(N__9334));
    CascadeBuf I__1774 (
            .O(N__9337),
            .I(N__9331));
    CascadeMux I__1773 (
            .O(N__9334),
            .I(N__9328));
    CascadeMux I__1772 (
            .O(N__9331),
            .I(N__9325));
    InMux I__1771 (
            .O(N__9328),
            .I(N__9322));
    InMux I__1770 (
            .O(N__9325),
            .I(N__9319));
    LocalMux I__1769 (
            .O(N__9322),
            .I(N__9316));
    LocalMux I__1768 (
            .O(N__9319),
            .I(N__9313));
    Sp12to4 I__1767 (
            .O(N__9316),
            .I(N__9310));
    Span12Mux_s8_v I__1766 (
            .O(N__9313),
            .I(N__9307));
    Span12Mux_s5_v I__1765 (
            .O(N__9310),
            .I(N__9304));
    Span12Mux_h I__1764 (
            .O(N__9307),
            .I(N__9301));
    Span12Mux_v I__1763 (
            .O(N__9304),
            .I(N__9298));
    Odrv12 I__1762 (
            .O(N__9301),
            .I(M_this_vga_signals_address_8));
    Odrv12 I__1761 (
            .O(N__9298),
            .I(M_this_vga_signals_address_8));
    InMux I__1760 (
            .O(N__9293),
            .I(\this_vga_signals.address_1_cry_0 ));
    CascadeMux I__1759 (
            .O(N__9290),
            .I(N__9287));
    CascadeBuf I__1758 (
            .O(N__9287),
            .I(N__9283));
    CascadeMux I__1757 (
            .O(N__9286),
            .I(N__9280));
    CascadeMux I__1756 (
            .O(N__9283),
            .I(N__9277));
    CascadeBuf I__1755 (
            .O(N__9280),
            .I(N__9274));
    CascadeBuf I__1754 (
            .O(N__9277),
            .I(N__9271));
    CascadeMux I__1753 (
            .O(N__9274),
            .I(N__9268));
    CascadeMux I__1752 (
            .O(N__9271),
            .I(N__9265));
    CascadeBuf I__1751 (
            .O(N__9268),
            .I(N__9262));
    CascadeBuf I__1750 (
            .O(N__9265),
            .I(N__9259));
    CascadeMux I__1749 (
            .O(N__9262),
            .I(N__9256));
    CascadeMux I__1748 (
            .O(N__9259),
            .I(N__9253));
    CascadeBuf I__1747 (
            .O(N__9256),
            .I(N__9250));
    CascadeBuf I__1746 (
            .O(N__9253),
            .I(N__9247));
    CascadeMux I__1745 (
            .O(N__9250),
            .I(N__9244));
    CascadeMux I__1744 (
            .O(N__9247),
            .I(N__9241));
    CascadeBuf I__1743 (
            .O(N__9244),
            .I(N__9238));
    CascadeBuf I__1742 (
            .O(N__9241),
            .I(N__9235));
    CascadeMux I__1741 (
            .O(N__9238),
            .I(N__9232));
    CascadeMux I__1740 (
            .O(N__9235),
            .I(N__9229));
    CascadeBuf I__1739 (
            .O(N__9232),
            .I(N__9226));
    CascadeBuf I__1738 (
            .O(N__9229),
            .I(N__9223));
    CascadeMux I__1737 (
            .O(N__9226),
            .I(N__9220));
    CascadeMux I__1736 (
            .O(N__9223),
            .I(N__9217));
    CascadeBuf I__1735 (
            .O(N__9220),
            .I(N__9214));
    CascadeBuf I__1734 (
            .O(N__9217),
            .I(N__9211));
    CascadeMux I__1733 (
            .O(N__9214),
            .I(N__9208));
    CascadeMux I__1732 (
            .O(N__9211),
            .I(N__9205));
    CascadeBuf I__1731 (
            .O(N__9208),
            .I(N__9202));
    CascadeBuf I__1730 (
            .O(N__9205),
            .I(N__9199));
    CascadeMux I__1729 (
            .O(N__9202),
            .I(N__9196));
    CascadeMux I__1728 (
            .O(N__9199),
            .I(N__9193));
    CascadeBuf I__1727 (
            .O(N__9196),
            .I(N__9190));
    CascadeBuf I__1726 (
            .O(N__9193),
            .I(N__9187));
    CascadeMux I__1725 (
            .O(N__9190),
            .I(N__9184));
    CascadeMux I__1724 (
            .O(N__9187),
            .I(N__9181));
    CascadeBuf I__1723 (
            .O(N__9184),
            .I(N__9178));
    CascadeBuf I__1722 (
            .O(N__9181),
            .I(N__9175));
    CascadeMux I__1721 (
            .O(N__9178),
            .I(N__9172));
    CascadeMux I__1720 (
            .O(N__9175),
            .I(N__9169));
    CascadeBuf I__1719 (
            .O(N__9172),
            .I(N__9166));
    CascadeBuf I__1718 (
            .O(N__9169),
            .I(N__9163));
    CascadeMux I__1717 (
            .O(N__9166),
            .I(N__9160));
    CascadeMux I__1716 (
            .O(N__9163),
            .I(N__9157));
    CascadeBuf I__1715 (
            .O(N__9160),
            .I(N__9154));
    CascadeBuf I__1714 (
            .O(N__9157),
            .I(N__9151));
    CascadeMux I__1713 (
            .O(N__9154),
            .I(N__9148));
    CascadeMux I__1712 (
            .O(N__9151),
            .I(N__9145));
    CascadeBuf I__1711 (
            .O(N__9148),
            .I(N__9142));
    CascadeBuf I__1710 (
            .O(N__9145),
            .I(N__9139));
    CascadeMux I__1709 (
            .O(N__9142),
            .I(N__9136));
    CascadeMux I__1708 (
            .O(N__9139),
            .I(N__9133));
    CascadeBuf I__1707 (
            .O(N__9136),
            .I(N__9130));
    CascadeBuf I__1706 (
            .O(N__9133),
            .I(N__9127));
    CascadeMux I__1705 (
            .O(N__9130),
            .I(N__9124));
    CascadeMux I__1704 (
            .O(N__9127),
            .I(N__9121));
    InMux I__1703 (
            .O(N__9124),
            .I(N__9118));
    CascadeBuf I__1702 (
            .O(N__9121),
            .I(N__9115));
    LocalMux I__1701 (
            .O(N__9118),
            .I(N__9112));
    CascadeMux I__1700 (
            .O(N__9115),
            .I(N__9109));
    Span4Mux_v I__1699 (
            .O(N__9112),
            .I(N__9106));
    InMux I__1698 (
            .O(N__9109),
            .I(N__9103));
    Span4Mux_v I__1697 (
            .O(N__9106),
            .I(N__9100));
    LocalMux I__1696 (
            .O(N__9103),
            .I(N__9097));
    Span4Mux_h I__1695 (
            .O(N__9100),
            .I(N__9094));
    Span4Mux_v I__1694 (
            .O(N__9097),
            .I(N__9091));
    Span4Mux_h I__1693 (
            .O(N__9094),
            .I(N__9088));
    Span4Mux_v I__1692 (
            .O(N__9091),
            .I(N__9085));
    Span4Mux_h I__1691 (
            .O(N__9088),
            .I(N__9080));
    Span4Mux_h I__1690 (
            .O(N__9085),
            .I(N__9080));
    Sp12to4 I__1689 (
            .O(N__9080),
            .I(N__9077));
    Odrv12 I__1688 (
            .O(N__9077),
            .I(M_this_vga_signals_address_9));
    InMux I__1687 (
            .O(N__9074),
            .I(\this_vga_signals.address_1_cry_1 ));
    CascadeMux I__1686 (
            .O(N__9071),
            .I(N__9068));
    CascadeBuf I__1685 (
            .O(N__9068),
            .I(N__9064));
    CascadeMux I__1684 (
            .O(N__9067),
            .I(N__9061));
    CascadeMux I__1683 (
            .O(N__9064),
            .I(N__9058));
    CascadeBuf I__1682 (
            .O(N__9061),
            .I(N__9055));
    CascadeBuf I__1681 (
            .O(N__9058),
            .I(N__9052));
    CascadeMux I__1680 (
            .O(N__9055),
            .I(N__9049));
    CascadeMux I__1679 (
            .O(N__9052),
            .I(N__9046));
    CascadeBuf I__1678 (
            .O(N__9049),
            .I(N__9043));
    CascadeBuf I__1677 (
            .O(N__9046),
            .I(N__9040));
    CascadeMux I__1676 (
            .O(N__9043),
            .I(N__9037));
    CascadeMux I__1675 (
            .O(N__9040),
            .I(N__9034));
    CascadeBuf I__1674 (
            .O(N__9037),
            .I(N__9031));
    CascadeBuf I__1673 (
            .O(N__9034),
            .I(N__9028));
    CascadeMux I__1672 (
            .O(N__9031),
            .I(N__9025));
    CascadeMux I__1671 (
            .O(N__9028),
            .I(N__9022));
    CascadeBuf I__1670 (
            .O(N__9025),
            .I(N__9019));
    CascadeBuf I__1669 (
            .O(N__9022),
            .I(N__9016));
    CascadeMux I__1668 (
            .O(N__9019),
            .I(N__9013));
    CascadeMux I__1667 (
            .O(N__9016),
            .I(N__9010));
    CascadeBuf I__1666 (
            .O(N__9013),
            .I(N__9007));
    CascadeBuf I__1665 (
            .O(N__9010),
            .I(N__9004));
    CascadeMux I__1664 (
            .O(N__9007),
            .I(N__9001));
    CascadeMux I__1663 (
            .O(N__9004),
            .I(N__8998));
    CascadeBuf I__1662 (
            .O(N__9001),
            .I(N__8995));
    CascadeBuf I__1661 (
            .O(N__8998),
            .I(N__8992));
    CascadeMux I__1660 (
            .O(N__8995),
            .I(N__8989));
    CascadeMux I__1659 (
            .O(N__8992),
            .I(N__8986));
    CascadeBuf I__1658 (
            .O(N__8989),
            .I(N__8983));
    CascadeBuf I__1657 (
            .O(N__8986),
            .I(N__8980));
    CascadeMux I__1656 (
            .O(N__8983),
            .I(N__8977));
    CascadeMux I__1655 (
            .O(N__8980),
            .I(N__8974));
    CascadeBuf I__1654 (
            .O(N__8977),
            .I(N__8971));
    CascadeBuf I__1653 (
            .O(N__8974),
            .I(N__8968));
    CascadeMux I__1652 (
            .O(N__8971),
            .I(N__8965));
    CascadeMux I__1651 (
            .O(N__8968),
            .I(N__8962));
    CascadeBuf I__1650 (
            .O(N__8965),
            .I(N__8959));
    CascadeBuf I__1649 (
            .O(N__8962),
            .I(N__8956));
    CascadeMux I__1648 (
            .O(N__8959),
            .I(N__8953));
    CascadeMux I__1647 (
            .O(N__8956),
            .I(N__8950));
    CascadeBuf I__1646 (
            .O(N__8953),
            .I(N__8947));
    CascadeBuf I__1645 (
            .O(N__8950),
            .I(N__8944));
    CascadeMux I__1644 (
            .O(N__8947),
            .I(N__8941));
    CascadeMux I__1643 (
            .O(N__8944),
            .I(N__8938));
    CascadeBuf I__1642 (
            .O(N__8941),
            .I(N__8935));
    CascadeBuf I__1641 (
            .O(N__8938),
            .I(N__8932));
    CascadeMux I__1640 (
            .O(N__8935),
            .I(N__8929));
    CascadeMux I__1639 (
            .O(N__8932),
            .I(N__8926));
    CascadeBuf I__1638 (
            .O(N__8929),
            .I(N__8923));
    CascadeBuf I__1637 (
            .O(N__8926),
            .I(N__8920));
    CascadeMux I__1636 (
            .O(N__8923),
            .I(N__8917));
    CascadeMux I__1635 (
            .O(N__8920),
            .I(N__8914));
    CascadeBuf I__1634 (
            .O(N__8917),
            .I(N__8911));
    CascadeBuf I__1633 (
            .O(N__8914),
            .I(N__8908));
    CascadeMux I__1632 (
            .O(N__8911),
            .I(N__8905));
    CascadeMux I__1631 (
            .O(N__8908),
            .I(N__8902));
    InMux I__1630 (
            .O(N__8905),
            .I(N__8899));
    CascadeBuf I__1629 (
            .O(N__8902),
            .I(N__8896));
    LocalMux I__1628 (
            .O(N__8899),
            .I(N__8893));
    CascadeMux I__1627 (
            .O(N__8896),
            .I(N__8890));
    Span4Mux_v I__1626 (
            .O(N__8893),
            .I(N__8887));
    InMux I__1625 (
            .O(N__8890),
            .I(N__8884));
    Span4Mux_h I__1624 (
            .O(N__8887),
            .I(N__8881));
    LocalMux I__1623 (
            .O(N__8884),
            .I(N__8878));
    Span4Mux_h I__1622 (
            .O(N__8881),
            .I(N__8875));
    Span4Mux_v I__1621 (
            .O(N__8878),
            .I(N__8872));
    Span4Mux_h I__1620 (
            .O(N__8875),
            .I(N__8869));
    Span4Mux_h I__1619 (
            .O(N__8872),
            .I(N__8866));
    Sp12to4 I__1618 (
            .O(N__8869),
            .I(N__8861));
    Sp12to4 I__1617 (
            .O(N__8866),
            .I(N__8861));
    Odrv12 I__1616 (
            .O(N__8861),
            .I(M_this_vga_signals_address_10));
    InMux I__1615 (
            .O(N__8858),
            .I(\this_vga_signals.address_1_cry_2 ));
    InMux I__1614 (
            .O(N__8855),
            .I(\this_vga_signals.address_1_cry_3 ));
    InMux I__1613 (
            .O(N__8852),
            .I(N__8849));
    LocalMux I__1612 (
            .O(N__8849),
            .I(N__8846));
    Span12Mux_s11_h I__1611 (
            .O(N__8846),
            .I(N__8843));
    Span12Mux_v I__1610 (
            .O(N__8843),
            .I(N__8840));
    Odrv12 I__1609 (
            .O(N__8840),
            .I(\this_vram.mem_out_bus4_2 ));
    InMux I__1608 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__1607 (
            .O(N__8834),
            .I(N__8831));
    Span4Mux_h I__1606 (
            .O(N__8831),
            .I(N__8828));
    Sp12to4 I__1605 (
            .O(N__8828),
            .I(N__8825));
    Span12Mux_v I__1604 (
            .O(N__8825),
            .I(N__8822));
    Span12Mux_h I__1603 (
            .O(N__8822),
            .I(N__8819));
    Odrv12 I__1602 (
            .O(N__8819),
            .I(\this_vram.mem_out_bus6_2 ));
    CascadeMux I__1601 (
            .O(N__8816),
            .I(\this_vram.mem_mem_4_1_RNI14PZ0Z11_cascade_ ));
    InMux I__1600 (
            .O(N__8813),
            .I(N__8810));
    LocalMux I__1599 (
            .O(N__8810),
            .I(\this_vram.mem_N_2345 ));
    CEMux I__1598 (
            .O(N__8807),
            .I(N__8804));
    LocalMux I__1597 (
            .O(N__8804),
            .I(N__8799));
    CEMux I__1596 (
            .O(N__8803),
            .I(N__8796));
    CEMux I__1595 (
            .O(N__8802),
            .I(N__8793));
    Span4Mux_s3_v I__1594 (
            .O(N__8799),
            .I(N__8786));
    LocalMux I__1593 (
            .O(N__8796),
            .I(N__8786));
    LocalMux I__1592 (
            .O(N__8793),
            .I(N__8786));
    Span4Mux_v I__1591 (
            .O(N__8786),
            .I(N__8783));
    Span4Mux_v I__1590 (
            .O(N__8783),
            .I(N__8780));
    Odrv4 I__1589 (
            .O(N__8780),
            .I(\this_vram.mem_WE_15 ));
    CascadeMux I__1588 (
            .O(N__8777),
            .I(\this_vga_signals.m24_0_1_cascade_ ));
    CascadeMux I__1587 (
            .O(N__8774),
            .I(\this_vga_signals.N_25_cascade_ ));
    InMux I__1586 (
            .O(N__8771),
            .I(N__8768));
    LocalMux I__1585 (
            .O(N__8768),
            .I(\this_vga_signals.m24_0_1_0 ));
    InMux I__1584 (
            .O(N__8765),
            .I(N__8762));
    LocalMux I__1583 (
            .O(N__8762),
            .I(N__8759));
    Odrv4 I__1582 (
            .O(N__8759),
            .I(\this_vram.mem_N_2327 ));
    InMux I__1581 (
            .O(N__8756),
            .I(N__8753));
    LocalMux I__1580 (
            .O(N__8753),
            .I(N__8750));
    Span12Mux_v I__1579 (
            .O(N__8750),
            .I(N__8747));
    Odrv12 I__1578 (
            .O(N__8747),
            .I(\this_vram.mem_N_2353 ));
    CascadeMux I__1577 (
            .O(N__8744),
            .I(\this_vram.mem_N_2355_cascade_ ));
    CascadeMux I__1576 (
            .O(N__8741),
            .I(N__8737));
    CascadeMux I__1575 (
            .O(N__8740),
            .I(N__8734));
    InMux I__1574 (
            .O(N__8737),
            .I(N__8727));
    InMux I__1573 (
            .O(N__8734),
            .I(N__8727));
    InMux I__1572 (
            .O(N__8733),
            .I(N__8724));
    InMux I__1571 (
            .O(N__8732),
            .I(N__8721));
    LocalMux I__1570 (
            .O(N__8727),
            .I(N__8716));
    LocalMux I__1569 (
            .O(N__8724),
            .I(N__8716));
    LocalMux I__1568 (
            .O(N__8721),
            .I(N__8713));
    Span4Mux_v I__1567 (
            .O(N__8716),
            .I(N__8707));
    Span4Mux_v I__1566 (
            .O(N__8713),
            .I(N__8707));
    InMux I__1565 (
            .O(N__8712),
            .I(N__8704));
    Odrv4 I__1564 (
            .O(N__8707),
            .I(\this_vram.mem_G_25_0 ));
    LocalMux I__1563 (
            .O(N__8704),
            .I(\this_vram.mem_G_25_0 ));
    IoInMux I__1562 (
            .O(N__8699),
            .I(N__8696));
    LocalMux I__1561 (
            .O(N__8696),
            .I(N__8693));
    Odrv12 I__1560 (
            .O(N__8693),
            .I(M_this_vram_read_data_1));
    InMux I__1559 (
            .O(N__8690),
            .I(N__8687));
    LocalMux I__1558 (
            .O(N__8687),
            .I(N__8684));
    Span4Mux_v I__1557 (
            .O(N__8684),
            .I(N__8681));
    Span4Mux_v I__1556 (
            .O(N__8681),
            .I(N__8678));
    Odrv4 I__1555 (
            .O(N__8678),
            .I(\this_vram.mem_out_bus4_4 ));
    InMux I__1554 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__1553 (
            .O(N__8672),
            .I(N__8669));
    Span4Mux_v I__1552 (
            .O(N__8669),
            .I(N__8666));
    Sp12to4 I__1551 (
            .O(N__8666),
            .I(N__8663));
    Span12Mux_h I__1550 (
            .O(N__8663),
            .I(N__8660));
    Span12Mux_v I__1549 (
            .O(N__8660),
            .I(N__8657));
    Odrv12 I__1548 (
            .O(N__8657),
            .I(\this_vram.mem_out_bus6_4 ));
    InMux I__1547 (
            .O(N__8654),
            .I(N__8651));
    LocalMux I__1546 (
            .O(N__8651),
            .I(\this_vram.mem_mem_4_2_RNI34PZ0Z11 ));
    CEMux I__1545 (
            .O(N__8648),
            .I(N__8645));
    LocalMux I__1544 (
            .O(N__8645),
            .I(N__8640));
    CEMux I__1543 (
            .O(N__8644),
            .I(N__8637));
    CEMux I__1542 (
            .O(N__8643),
            .I(N__8634));
    Span4Mux_v I__1541 (
            .O(N__8640),
            .I(N__8627));
    LocalMux I__1540 (
            .O(N__8637),
            .I(N__8627));
    LocalMux I__1539 (
            .O(N__8634),
            .I(N__8627));
    Span4Mux_v I__1538 (
            .O(N__8627),
            .I(N__8624));
    Odrv4 I__1537 (
            .O(N__8624),
            .I(\this_vram.mem_WE_18 ));
    InMux I__1536 (
            .O(N__8621),
            .I(N__8618));
    LocalMux I__1535 (
            .O(N__8618),
            .I(N__8615));
    Span4Mux_v I__1534 (
            .O(N__8615),
            .I(N__8612));
    Sp12to4 I__1533 (
            .O(N__8612),
            .I(N__8609));
    Span12Mux_h I__1532 (
            .O(N__8609),
            .I(N__8606));
    Span12Mux_v I__1531 (
            .O(N__8606),
            .I(N__8603));
    Odrv12 I__1530 (
            .O(N__8603),
            .I(\this_vram.mem_out_bus6_1 ));
    InMux I__1529 (
            .O(N__8600),
            .I(N__8597));
    LocalMux I__1528 (
            .O(N__8597),
            .I(N__8594));
    Span4Mux_v I__1527 (
            .O(N__8594),
            .I(N__8591));
    Odrv4 I__1526 (
            .O(N__8591),
            .I(\this_vram.mem_out_bus4_1 ));
    InMux I__1525 (
            .O(N__8588),
            .I(N__8585));
    LocalMux I__1524 (
            .O(N__8585),
            .I(N__8582));
    Span4Mux_v I__1523 (
            .O(N__8582),
            .I(N__8579));
    Span4Mux_v I__1522 (
            .O(N__8579),
            .I(N__8576));
    Odrv4 I__1521 (
            .O(N__8576),
            .I(\this_vram.mem_out_bus5_1 ));
    InMux I__1520 (
            .O(N__8573),
            .I(N__8570));
    LocalMux I__1519 (
            .O(N__8570),
            .I(N__8567));
    Span4Mux_v I__1518 (
            .O(N__8567),
            .I(N__8564));
    Sp12to4 I__1517 (
            .O(N__8564),
            .I(N__8561));
    Span12Mux_h I__1516 (
            .O(N__8561),
            .I(N__8558));
    Span12Mux_v I__1515 (
            .O(N__8558),
            .I(N__8555));
    Odrv12 I__1514 (
            .O(N__8555),
            .I(\this_vram.mem_out_bus7_1 ));
    InMux I__1513 (
            .O(N__8552),
            .I(N__8549));
    LocalMux I__1512 (
            .O(N__8549),
            .I(\this_vram.mem_mem_4_0_RNIV3P11Z0Z_0 ));
    CascadeMux I__1511 (
            .O(N__8546),
            .I(\this_vram.mem_mem_5_0_RNI18R11Z0Z_0_cascade_ ));
    InMux I__1510 (
            .O(N__8543),
            .I(N__8540));
    LocalMux I__1509 (
            .O(N__8540),
            .I(N__8537));
    Odrv12 I__1508 (
            .O(N__8537),
            .I(\this_vram.mem_N_2354 ));
    CEMux I__1507 (
            .O(N__8534),
            .I(N__8530));
    CEMux I__1506 (
            .O(N__8533),
            .I(N__8527));
    LocalMux I__1505 (
            .O(N__8530),
            .I(N__8521));
    LocalMux I__1504 (
            .O(N__8527),
            .I(N__8521));
    CEMux I__1503 (
            .O(N__8526),
            .I(N__8518));
    Span4Mux_v I__1502 (
            .O(N__8521),
            .I(N__8513));
    LocalMux I__1501 (
            .O(N__8518),
            .I(N__8513));
    Span4Mux_v I__1500 (
            .O(N__8513),
            .I(N__8510));
    Odrv4 I__1499 (
            .O(N__8510),
            .I(\this_vram.mem_WE_24 ));
    InMux I__1498 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__1497 (
            .O(N__8504),
            .I(N__8501));
    Odrv12 I__1496 (
            .O(N__8501),
            .I(\this_vram.mem_mem_0_0_RNILGF11Z0Z_0 ));
    CascadeMux I__1495 (
            .O(N__8498),
            .I(\this_vram.mem_mem_2_0_RNIPOJ11Z0Z_0_cascade_ ));
    InMux I__1494 (
            .O(N__8495),
            .I(N__8492));
    LocalMux I__1493 (
            .O(N__8492),
            .I(N__8489));
    Span4Mux_v I__1492 (
            .O(N__8489),
            .I(N__8486));
    Sp12to4 I__1491 (
            .O(N__8486),
            .I(N__8483));
    Span12Mux_h I__1490 (
            .O(N__8483),
            .I(N__8480));
    Span12Mux_v I__1489 (
            .O(N__8480),
            .I(N__8477));
    Odrv12 I__1488 (
            .O(N__8477),
            .I(\this_vram.mem_out_bus6_0 ));
    InMux I__1487 (
            .O(N__8474),
            .I(N__8471));
    LocalMux I__1486 (
            .O(N__8471),
            .I(N__8468));
    Span4Mux_v I__1485 (
            .O(N__8468),
            .I(N__8465));
    Span4Mux_v I__1484 (
            .O(N__8465),
            .I(N__8462));
    Odrv4 I__1483 (
            .O(N__8462),
            .I(\this_vram.mem_out_bus4_0 ));
    CEMux I__1482 (
            .O(N__8459),
            .I(N__8455));
    CEMux I__1481 (
            .O(N__8458),
            .I(N__8452));
    LocalMux I__1480 (
            .O(N__8455),
            .I(N__8446));
    LocalMux I__1479 (
            .O(N__8452),
            .I(N__8446));
    CEMux I__1478 (
            .O(N__8451),
            .I(N__8443));
    Span4Mux_v I__1477 (
            .O(N__8446),
            .I(N__8438));
    LocalMux I__1476 (
            .O(N__8443),
            .I(N__8438));
    Span4Mux_v I__1475 (
            .O(N__8438),
            .I(N__8435));
    Span4Mux_v I__1474 (
            .O(N__8435),
            .I(N__8432));
    Odrv4 I__1473 (
            .O(N__8432),
            .I(\this_vram.mem_WE_27 ));
    InMux I__1472 (
            .O(N__8429),
            .I(N__8426));
    LocalMux I__1471 (
            .O(N__8426),
            .I(N__8423));
    Span4Mux_v I__1470 (
            .O(N__8423),
            .I(N__8420));
    Span4Mux_v I__1469 (
            .O(N__8420),
            .I(N__8417));
    Span4Mux_v I__1468 (
            .O(N__8417),
            .I(N__8414));
    Span4Mux_v I__1467 (
            .O(N__8414),
            .I(N__8411));
    Odrv4 I__1466 (
            .O(N__8411),
            .I(\this_vram.mem_out_bus5_0 ));
    InMux I__1465 (
            .O(N__8408),
            .I(N__8405));
    LocalMux I__1464 (
            .O(N__8405),
            .I(N__8402));
    Span4Mux_v I__1463 (
            .O(N__8402),
            .I(N__8399));
    Sp12to4 I__1462 (
            .O(N__8399),
            .I(N__8396));
    Span12Mux_h I__1461 (
            .O(N__8396),
            .I(N__8393));
    Odrv12 I__1460 (
            .O(N__8393),
            .I(\this_vram.mem_out_bus7_0 ));
    CascadeMux I__1459 (
            .O(N__8390),
            .I(\this_vram.mem_mem_5_0_RNI18RZ0Z11_cascade_ ));
    InMux I__1458 (
            .O(N__8387),
            .I(N__8384));
    LocalMux I__1457 (
            .O(N__8384),
            .I(\this_vram.mem_mem_4_0_RNIV3PZ0Z11 ));
    InMux I__1456 (
            .O(N__8381),
            .I(N__8378));
    LocalMux I__1455 (
            .O(N__8378),
            .I(N__8375));
    Span4Mux_h I__1454 (
            .O(N__8375),
            .I(N__8372));
    Odrv4 I__1453 (
            .O(N__8372),
            .I(\this_vram.mem_N_2363 ));
    InMux I__1452 (
            .O(N__8369),
            .I(N__8366));
    LocalMux I__1451 (
            .O(N__8366),
            .I(N__8363));
    Odrv4 I__1450 (
            .O(N__8363),
            .I(\this_vram.mem_N_2344 ));
    InMux I__1449 (
            .O(N__8360),
            .I(N__8357));
    LocalMux I__1448 (
            .O(N__8357),
            .I(\this_vram.mem_N_2346 ));
    CascadeMux I__1447 (
            .O(N__8354),
            .I(\this_vram.mem_G_25_0_cascade_ ));
    IoInMux I__1446 (
            .O(N__8351),
            .I(N__8348));
    LocalMux I__1445 (
            .O(N__8348),
            .I(N__8345));
    Odrv12 I__1444 (
            .O(N__8345),
            .I(M_this_vram_read_data_2));
    CEMux I__1443 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1442 (
            .O(N__8339),
            .I(N__8334));
    CEMux I__1441 (
            .O(N__8338),
            .I(N__8331));
    CEMux I__1440 (
            .O(N__8337),
            .I(N__8328));
    Span4Mux_v I__1439 (
            .O(N__8334),
            .I(N__8321));
    LocalMux I__1438 (
            .O(N__8331),
            .I(N__8321));
    LocalMux I__1437 (
            .O(N__8328),
            .I(N__8321));
    Odrv4 I__1436 (
            .O(N__8321),
            .I(\this_vram.mem_WE_21 ));
    InMux I__1435 (
            .O(N__8318),
            .I(N__8315));
    LocalMux I__1434 (
            .O(N__8315),
            .I(\this_vram.mem_out_bus2_4 ));
    InMux I__1433 (
            .O(N__8312),
            .I(N__8309));
    LocalMux I__1432 (
            .O(N__8309),
            .I(N__8306));
    Span4Mux_v I__1431 (
            .O(N__8306),
            .I(N__8303));
    Odrv4 I__1430 (
            .O(N__8303),
            .I(\this_vram.mem_out_bus3_4 ));
    InMux I__1429 (
            .O(N__8300),
            .I(N__8297));
    LocalMux I__1428 (
            .O(N__8297),
            .I(N__8294));
    Span4Mux_v I__1427 (
            .O(N__8294),
            .I(N__8291));
    Odrv4 I__1426 (
            .O(N__8291),
            .I(\this_vram.mem_mem_0_2_RNIPGFZ0Z11 ));
    CascadeMux I__1425 (
            .O(N__8288),
            .I(\this_vram.mem_mem_2_2_RNITOJZ0Z11_cascade_ ));
    CascadeMux I__1424 (
            .O(N__8285),
            .I(\this_vram.mem_N_2326_cascade_ ));
    CascadeMux I__1423 (
            .O(N__8282),
            .I(N__8279));
    InMux I__1422 (
            .O(N__8279),
            .I(N__8276));
    LocalMux I__1421 (
            .O(N__8276),
            .I(N__8273));
    Odrv4 I__1420 (
            .O(N__8273),
            .I(\this_vram.mem_N_2373 ));
    IoInMux I__1419 (
            .O(N__8270),
            .I(N__8267));
    LocalMux I__1418 (
            .O(N__8267),
            .I(N__8264));
    Span4Mux_s1_h I__1417 (
            .O(N__8264),
            .I(N__8261));
    Sp12to4 I__1416 (
            .O(N__8261),
            .I(N__8258));
    Span12Mux_v I__1415 (
            .O(N__8258),
            .I(N__8255));
    Odrv12 I__1414 (
            .O(N__8255),
            .I(M_this_vram_read_data_5));
    InMux I__1413 (
            .O(N__8252),
            .I(N__8249));
    LocalMux I__1412 (
            .O(N__8249),
            .I(N__8246));
    Odrv4 I__1411 (
            .O(N__8246),
            .I(\this_vram.mem_N_2328 ));
    IoInMux I__1410 (
            .O(N__8243),
            .I(N__8240));
    LocalMux I__1409 (
            .O(N__8240),
            .I(N__8237));
    IoSpan4Mux I__1408 (
            .O(N__8237),
            .I(N__8234));
    Sp12to4 I__1407 (
            .O(N__8234),
            .I(N__8231));
    Span12Mux_s6_h I__1406 (
            .O(N__8231),
            .I(N__8228));
    Odrv12 I__1405 (
            .O(N__8228),
            .I(M_this_vram_read_data_4));
    InMux I__1404 (
            .O(N__8225),
            .I(N__8222));
    LocalMux I__1403 (
            .O(N__8222),
            .I(N__8219));
    Odrv12 I__1402 (
            .O(N__8219),
            .I(\this_vram.mem_N_2337 ));
    IoInMux I__1401 (
            .O(N__8216),
            .I(N__8213));
    LocalMux I__1400 (
            .O(N__8213),
            .I(N__8210));
    Span4Mux_s3_h I__1399 (
            .O(N__8210),
            .I(N__8207));
    Span4Mux_v I__1398 (
            .O(N__8207),
            .I(N__8204));
    Odrv4 I__1397 (
            .O(N__8204),
            .I(M_this_vram_read_data_3));
    InMux I__1396 (
            .O(N__8201),
            .I(N__8198));
    LocalMux I__1395 (
            .O(N__8198),
            .I(N__8195));
    Span4Mux_v I__1394 (
            .O(N__8195),
            .I(N__8192));
    Odrv4 I__1393 (
            .O(N__8192),
            .I(\this_vram.mem_out_bus0_1 ));
    InMux I__1392 (
            .O(N__8189),
            .I(N__8186));
    LocalMux I__1391 (
            .O(N__8186),
            .I(\this_vram.mem_out_bus1_1 ));
    InMux I__1390 (
            .O(N__8183),
            .I(N__8180));
    LocalMux I__1389 (
            .O(N__8180),
            .I(N__8177));
    Span4Mux_v I__1388 (
            .O(N__8177),
            .I(N__8174));
    Odrv4 I__1387 (
            .O(N__8174),
            .I(\this_vram.mem_out_bus3_1 ));
    InMux I__1386 (
            .O(N__8171),
            .I(N__8168));
    LocalMux I__1385 (
            .O(N__8168),
            .I(\this_vram.mem_out_bus2_1 ));
    InMux I__1384 (
            .O(N__8165),
            .I(N__8162));
    LocalMux I__1383 (
            .O(N__8162),
            .I(N__8159));
    Odrv12 I__1382 (
            .O(N__8159),
            .I(\this_vram.mem_mem_0_1_RNINGF11Z0Z_0 ));
    CascadeMux I__1381 (
            .O(N__8156),
            .I(\this_vram.mem_mem_2_1_RNIROJ11Z0Z_0_cascade_ ));
    InMux I__1380 (
            .O(N__8153),
            .I(N__8150));
    LocalMux I__1379 (
            .O(N__8150),
            .I(N__8147));
    Sp12to4 I__1378 (
            .O(N__8147),
            .I(N__8144));
    Span12Mux_v I__1377 (
            .O(N__8144),
            .I(N__8141));
    Odrv12 I__1376 (
            .O(N__8141),
            .I(\this_vram.mem_out_bus4_3 ));
    InMux I__1375 (
            .O(N__8138),
            .I(N__8135));
    LocalMux I__1374 (
            .O(N__8135),
            .I(N__8132));
    Span4Mux_v I__1373 (
            .O(N__8132),
            .I(N__8129));
    Sp12to4 I__1372 (
            .O(N__8129),
            .I(N__8126));
    Span12Mux_h I__1371 (
            .O(N__8126),
            .I(N__8123));
    Span12Mux_v I__1370 (
            .O(N__8123),
            .I(N__8120));
    Odrv12 I__1369 (
            .O(N__8120),
            .I(\this_vram.mem_out_bus6_3 ));
    CascadeMux I__1368 (
            .O(N__8117),
            .I(\this_vram.mem_mem_4_1_RNI14P11Z0Z_0_cascade_ ));
    CascadeMux I__1367 (
            .O(N__8114),
            .I(\this_vram.mem_N_2336_cascade_ ));
    InMux I__1366 (
            .O(N__8111),
            .I(N__8108));
    LocalMux I__1365 (
            .O(N__8108),
            .I(\this_vram.mem_N_2335 ));
    InMux I__1364 (
            .O(N__8105),
            .I(N__8102));
    LocalMux I__1363 (
            .O(N__8102),
            .I(N__8099));
    Span4Mux_v I__1362 (
            .O(N__8099),
            .I(N__8096));
    Odrv4 I__1361 (
            .O(N__8096),
            .I(\this_vram.mem_out_bus3_2 ));
    InMux I__1360 (
            .O(N__8093),
            .I(N__8090));
    LocalMux I__1359 (
            .O(N__8090),
            .I(\this_vram.mem_out_bus2_2 ));
    CascadeMux I__1358 (
            .O(N__8087),
            .I(\this_vram.mem_mem_2_1_RNIROJZ0Z11_cascade_ ));
    InMux I__1357 (
            .O(N__8084),
            .I(N__8081));
    LocalMux I__1356 (
            .O(N__8081),
            .I(N__8078));
    Span4Mux_v I__1355 (
            .O(N__8078),
            .I(N__8075));
    Odrv4 I__1354 (
            .O(N__8075),
            .I(\this_vram.mem_mem_0_1_RNINGFZ0Z11 ));
    InMux I__1353 (
            .O(N__8072),
            .I(N__8069));
    LocalMux I__1352 (
            .O(N__8069),
            .I(N__8066));
    Span4Mux_v I__1351 (
            .O(N__8066),
            .I(N__8063));
    Odrv4 I__1350 (
            .O(N__8063),
            .I(\this_vram.mem_out_bus3_5 ));
    InMux I__1349 (
            .O(N__8060),
            .I(N__8057));
    LocalMux I__1348 (
            .O(N__8057),
            .I(\this_vram.mem_out_bus2_5 ));
    InMux I__1347 (
            .O(N__8054),
            .I(N__8051));
    LocalMux I__1346 (
            .O(N__8051),
            .I(N__8048));
    Span4Mux_v I__1345 (
            .O(N__8048),
            .I(N__8045));
    Odrv4 I__1344 (
            .O(N__8045),
            .I(\this_vram.mem_mem_0_2_RNIPGF11Z0Z_0 ));
    CascadeMux I__1343 (
            .O(N__8042),
            .I(\this_vram.mem_mem_2_2_RNITOJ11Z0Z_0_cascade_ ));
    CascadeMux I__1342 (
            .O(N__8039),
            .I(\this_vram.mem_N_2371_cascade_ ));
    InMux I__1341 (
            .O(N__8036),
            .I(N__8033));
    LocalMux I__1340 (
            .O(N__8033),
            .I(N__8030));
    Span4Mux_v I__1339 (
            .O(N__8030),
            .I(N__8027));
    Odrv4 I__1338 (
            .O(N__8027),
            .I(\this_vram.mem_out_bus0_3 ));
    InMux I__1337 (
            .O(N__8024),
            .I(N__8021));
    LocalMux I__1336 (
            .O(N__8021),
            .I(\this_vram.mem_out_bus1_3 ));
    InMux I__1335 (
            .O(N__8018),
            .I(N__8015));
    LocalMux I__1334 (
            .O(N__8015),
            .I(N__8012));
    Span4Mux_v I__1333 (
            .O(N__8012),
            .I(N__8009));
    Odrv4 I__1332 (
            .O(N__8009),
            .I(\this_vram.mem_out_bus0_4 ));
    InMux I__1331 (
            .O(N__8006),
            .I(N__8003));
    LocalMux I__1330 (
            .O(N__8003),
            .I(\this_vram.mem_out_bus1_4 ));
    InMux I__1329 (
            .O(N__8000),
            .I(N__7997));
    LocalMux I__1328 (
            .O(N__7997),
            .I(\this_vram.mem_out_bus1_5 ));
    InMux I__1327 (
            .O(N__7994),
            .I(N__7991));
    LocalMux I__1326 (
            .O(N__7991),
            .I(N__7988));
    Span4Mux_v I__1325 (
            .O(N__7988),
            .I(N__7985));
    Odrv4 I__1324 (
            .O(N__7985),
            .I(\this_vram.mem_out_bus0_5 ));
    InMux I__1323 (
            .O(N__7982),
            .I(N__7979));
    LocalMux I__1322 (
            .O(N__7979),
            .I(N__7976));
    Span4Mux_v I__1321 (
            .O(N__7976),
            .I(N__7973));
    Odrv4 I__1320 (
            .O(N__7973),
            .I(\this_vram.mem_out_bus3_0 ));
    InMux I__1319 (
            .O(N__7970),
            .I(N__7967));
    LocalMux I__1318 (
            .O(N__7967),
            .I(\this_vram.mem_out_bus2_0 ));
    InMux I__1317 (
            .O(N__7964),
            .I(N__7961));
    LocalMux I__1316 (
            .O(N__7961),
            .I(N__7958));
    Odrv12 I__1315 (
            .O(N__7958),
            .I(\this_vram.mem_mem_0_0_RNILGFZ0Z11 ));
    CascadeMux I__1314 (
            .O(N__7955),
            .I(\this_vram.mem_mem_2_0_RNIPOJZ0Z11_cascade_ ));
    InMux I__1313 (
            .O(N__7952),
            .I(N__7949));
    LocalMux I__1312 (
            .O(N__7949),
            .I(N__7946));
    Odrv4 I__1311 (
            .O(N__7946),
            .I(\this_vram.mem_N_2362 ));
    CascadeMux I__1310 (
            .O(N__7943),
            .I(\this_vram.mem_N_2364_cascade_ ));
    IoInMux I__1309 (
            .O(N__7940),
            .I(N__7937));
    LocalMux I__1308 (
            .O(N__7937),
            .I(N__7934));
    Span12Mux_s6_h I__1307 (
            .O(N__7934),
            .I(N__7931));
    Odrv12 I__1306 (
            .O(N__7931),
            .I(M_this_vram_read_data_0));
    InMux I__1305 (
            .O(N__7928),
            .I(N__7925));
    LocalMux I__1304 (
            .O(N__7925),
            .I(N__7922));
    Span4Mux_v I__1303 (
            .O(N__7922),
            .I(N__7919));
    Odrv4 I__1302 (
            .O(N__7919),
            .I(\this_vram.mem_out_bus3_3 ));
    InMux I__1301 (
            .O(N__7916),
            .I(N__7913));
    LocalMux I__1300 (
            .O(N__7913),
            .I(\this_vram.mem_out_bus2_3 ));
    IoInMux I__1299 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__1298 (
            .O(N__7907),
            .I(N__7904));
    Span12Mux_s0_h I__1297 (
            .O(N__7904),
            .I(N__7901));
    Odrv12 I__1296 (
            .O(N__7901),
            .I(this_vga_signals_N_170_i));
    IoInMux I__1295 (
            .O(N__7898),
            .I(N__7895));
    LocalMux I__1294 (
            .O(N__7895),
            .I(this_vga_signals_N_171_i));
    IoInMux I__1293 (
            .O(N__7892),
            .I(N__7889));
    LocalMux I__1292 (
            .O(N__7889),
            .I(N__7884));
    IoInMux I__1291 (
            .O(N__7888),
            .I(N__7881));
    IoInMux I__1290 (
            .O(N__7887),
            .I(N__7878));
    Span4Mux_s0_h I__1289 (
            .O(N__7884),
            .I(N__7874));
    LocalMux I__1288 (
            .O(N__7881),
            .I(N__7869));
    LocalMux I__1287 (
            .O(N__7878),
            .I(N__7869));
    IoInMux I__1286 (
            .O(N__7877),
            .I(N__7866));
    Span4Mux_v I__1285 (
            .O(N__7874),
            .I(N__7863));
    IoSpan4Mux I__1284 (
            .O(N__7869),
            .I(N__7858));
    LocalMux I__1283 (
            .O(N__7866),
            .I(N__7858));
    Span4Mux_v I__1282 (
            .O(N__7863),
            .I(N__7855));
    IoSpan4Mux I__1281 (
            .O(N__7858),
            .I(N__7852));
    Span4Mux_v I__1280 (
            .O(N__7855),
            .I(N__7847));
    Span4Mux_s0_h I__1279 (
            .O(N__7852),
            .I(N__7847));
    Span4Mux_v I__1278 (
            .O(N__7847),
            .I(N__7842));
    IoInMux I__1277 (
            .O(N__7846),
            .I(N__7839));
    IoInMux I__1276 (
            .O(N__7845),
            .I(N__7836));
    Odrv4 I__1275 (
            .O(N__7842),
            .I(rgb5_i));
    LocalMux I__1274 (
            .O(N__7839),
            .I(rgb5_i));
    LocalMux I__1273 (
            .O(N__7836),
            .I(rgb5_i));
    IoInMux I__1272 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__1271 (
            .O(N__7826),
            .I(vsync_c));
    IoInMux I__1270 (
            .O(N__7823),
            .I(N__7820));
    LocalMux I__1269 (
            .O(N__7820),
            .I(N__7817));
    Span4Mux_s1_h I__1268 (
            .O(N__7817),
            .I(N__7814));
    Span4Mux_v I__1267 (
            .O(N__7814),
            .I(N__7811));
    Odrv4 I__1266 (
            .O(N__7811),
            .I(this_vga_signals_N_94_i));
    InMux I__1265 (
            .O(N__7808),
            .I(N__7805));
    LocalMux I__1264 (
            .O(N__7805),
            .I(N__7802));
    Span4Mux_v I__1263 (
            .O(N__7802),
            .I(N__7799));
    Odrv4 I__1262 (
            .O(N__7799),
            .I(\this_vram.mem_out_bus0_0 ));
    InMux I__1261 (
            .O(N__7796),
            .I(N__7793));
    LocalMux I__1260 (
            .O(N__7793),
            .I(\this_vram.mem_out_bus1_0 ));
    InMux I__1259 (
            .O(N__7790),
            .I(N__7787));
    LocalMux I__1258 (
            .O(N__7787),
            .I(N__7784));
    Span4Mux_v I__1257 (
            .O(N__7784),
            .I(N__7781));
    Odrv4 I__1256 (
            .O(N__7781),
            .I(\this_vram.mem_out_bus0_2 ));
    InMux I__1255 (
            .O(N__7778),
            .I(N__7775));
    LocalMux I__1254 (
            .O(N__7775),
            .I(\this_vram.mem_out_bus1_2 ));
    InMux I__1253 (
            .O(N__7772),
            .I(N__7767));
    InMux I__1252 (
            .O(N__7771),
            .I(N__7762));
    InMux I__1251 (
            .O(N__7770),
            .I(N__7759));
    LocalMux I__1250 (
            .O(N__7767),
            .I(N__7755));
    InMux I__1249 (
            .O(N__7766),
            .I(N__7752));
    InMux I__1248 (
            .O(N__7765),
            .I(N__7749));
    LocalMux I__1247 (
            .O(N__7762),
            .I(N__7745));
    LocalMux I__1246 (
            .O(N__7759),
            .I(N__7742));
    InMux I__1245 (
            .O(N__7758),
            .I(N__7739));
    Span12Mux_s9_h I__1244 (
            .O(N__7755),
            .I(N__7735));
    LocalMux I__1243 (
            .O(N__7752),
            .I(N__7732));
    LocalMux I__1242 (
            .O(N__7749),
            .I(N__7729));
    InMux I__1241 (
            .O(N__7748),
            .I(N__7726));
    Span4Mux_h I__1240 (
            .O(N__7745),
            .I(N__7723));
    Span4Mux_v I__1239 (
            .O(N__7742),
            .I(N__7720));
    LocalMux I__1238 (
            .O(N__7739),
            .I(N__7717));
    InMux I__1237 (
            .O(N__7738),
            .I(N__7714));
    Span12Mux_h I__1236 (
            .O(N__7735),
            .I(N__7709));
    Span12Mux_s9_h I__1235 (
            .O(N__7732),
            .I(N__7706));
    Span4Mux_h I__1234 (
            .O(N__7729),
            .I(N__7703));
    LocalMux I__1233 (
            .O(N__7726),
            .I(N__7700));
    Sp12to4 I__1232 (
            .O(N__7723),
            .I(N__7697));
    Span4Mux_h I__1231 (
            .O(N__7720),
            .I(N__7694));
    Span12Mux_s10_h I__1230 (
            .O(N__7717),
            .I(N__7691));
    LocalMux I__1229 (
            .O(N__7714),
            .I(N__7688));
    InMux I__1228 (
            .O(N__7713),
            .I(N__7685));
    InMux I__1227 (
            .O(N__7712),
            .I(N__7682));
    Span12Mux_v I__1226 (
            .O(N__7709),
            .I(N__7677));
    Span12Mux_h I__1225 (
            .O(N__7706),
            .I(N__7677));
    Sp12to4 I__1224 (
            .O(N__7703),
            .I(N__7674));
    Span4Mux_h I__1223 (
            .O(N__7700),
            .I(N__7671));
    Span12Mux_v I__1222 (
            .O(N__7697),
            .I(N__7666));
    Sp12to4 I__1221 (
            .O(N__7694),
            .I(N__7666));
    Span12Mux_v I__1220 (
            .O(N__7691),
            .I(N__7661));
    Span12Mux_s10_h I__1219 (
            .O(N__7688),
            .I(N__7661));
    LocalMux I__1218 (
            .O(N__7685),
            .I(N__7658));
    LocalMux I__1217 (
            .O(N__7682),
            .I(N__7655));
    Span12Mux_v I__1216 (
            .O(N__7677),
            .I(N__7652));
    Span12Mux_v I__1215 (
            .O(N__7674),
            .I(N__7647));
    Sp12to4 I__1214 (
            .O(N__7671),
            .I(N__7647));
    Span12Mux_h I__1213 (
            .O(N__7666),
            .I(N__7640));
    Span12Mux_v I__1212 (
            .O(N__7661),
            .I(N__7640));
    Span12Mux_s10_h I__1211 (
            .O(N__7658),
            .I(N__7640));
    Span4Mux_h I__1210 (
            .O(N__7655),
            .I(N__7637));
    Odrv12 I__1209 (
            .O(N__7652),
            .I(write_data_c_1));
    Odrv12 I__1208 (
            .O(N__7647),
            .I(write_data_c_1));
    Odrv12 I__1207 (
            .O(N__7640),
            .I(write_data_c_1));
    Odrv4 I__1206 (
            .O(N__7637),
            .I(write_data_c_1));
    InMux I__1205 (
            .O(N__7628),
            .I(N__7625));
    LocalMux I__1204 (
            .O(N__7625),
            .I(N__7621));
    InMux I__1203 (
            .O(N__7624),
            .I(N__7618));
    Span4Mux_h I__1202 (
            .O(N__7621),
            .I(N__7615));
    LocalMux I__1201 (
            .O(N__7618),
            .I(N__7611));
    Span4Mux_v I__1200 (
            .O(N__7615),
            .I(N__7607));
    InMux I__1199 (
            .O(N__7614),
            .I(N__7604));
    Span4Mux_h I__1198 (
            .O(N__7611),
            .I(N__7601));
    InMux I__1197 (
            .O(N__7610),
            .I(N__7597));
    Span4Mux_v I__1196 (
            .O(N__7607),
            .I(N__7594));
    LocalMux I__1195 (
            .O(N__7604),
            .I(N__7591));
    Span4Mux_v I__1194 (
            .O(N__7601),
            .I(N__7587));
    InMux I__1193 (
            .O(N__7600),
            .I(N__7584));
    LocalMux I__1192 (
            .O(N__7597),
            .I(N__7581));
    Span4Mux_v I__1191 (
            .O(N__7594),
            .I(N__7575));
    Span4Mux_h I__1190 (
            .O(N__7591),
            .I(N__7575));
    InMux I__1189 (
            .O(N__7590),
            .I(N__7572));
    Span4Mux_v I__1188 (
            .O(N__7587),
            .I(N__7569));
    LocalMux I__1187 (
            .O(N__7584),
            .I(N__7566));
    Span4Mux_s2_v I__1186 (
            .O(N__7581),
            .I(N__7562));
    InMux I__1185 (
            .O(N__7580),
            .I(N__7559));
    Span4Mux_h I__1184 (
            .O(N__7575),
            .I(N__7556));
    LocalMux I__1183 (
            .O(N__7572),
            .I(N__7553));
    Span4Mux_v I__1182 (
            .O(N__7569),
            .I(N__7548));
    Span4Mux_h I__1181 (
            .O(N__7566),
            .I(N__7548));
    InMux I__1180 (
            .O(N__7565),
            .I(N__7545));
    Span4Mux_v I__1179 (
            .O(N__7562),
            .I(N__7540));
    LocalMux I__1178 (
            .O(N__7559),
            .I(N__7540));
    Span4Mux_h I__1177 (
            .O(N__7556),
            .I(N__7537));
    Span4Mux_h I__1176 (
            .O(N__7553),
            .I(N__7534));
    Span4Mux_h I__1175 (
            .O(N__7548),
            .I(N__7530));
    LocalMux I__1174 (
            .O(N__7545),
            .I(N__7527));
    Span4Mux_v I__1173 (
            .O(N__7540),
            .I(N__7524));
    Span4Mux_h I__1172 (
            .O(N__7537),
            .I(N__7519));
    Span4Mux_v I__1171 (
            .O(N__7534),
            .I(N__7519));
    InMux I__1170 (
            .O(N__7533),
            .I(N__7516));
    Span4Mux_h I__1169 (
            .O(N__7530),
            .I(N__7513));
    Span4Mux_h I__1168 (
            .O(N__7527),
            .I(N__7510));
    Sp12to4 I__1167 (
            .O(N__7524),
            .I(N__7506));
    Span4Mux_v I__1166 (
            .O(N__7519),
            .I(N__7503));
    LocalMux I__1165 (
            .O(N__7516),
            .I(N__7500));
    Span4Mux_h I__1164 (
            .O(N__7513),
            .I(N__7495));
    Span4Mux_v I__1163 (
            .O(N__7510),
            .I(N__7495));
    InMux I__1162 (
            .O(N__7509),
            .I(N__7492));
    Span12Mux_s10_h I__1161 (
            .O(N__7506),
            .I(N__7489));
    Span4Mux_v I__1160 (
            .O(N__7503),
            .I(N__7484));
    Span4Mux_h I__1159 (
            .O(N__7500),
            .I(N__7484));
    Span4Mux_v I__1158 (
            .O(N__7495),
            .I(N__7481));
    LocalMux I__1157 (
            .O(N__7492),
            .I(N__7478));
    Span12Mux_v I__1156 (
            .O(N__7489),
            .I(N__7475));
    Span4Mux_v I__1155 (
            .O(N__7484),
            .I(N__7472));
    Span4Mux_v I__1154 (
            .O(N__7481),
            .I(N__7467));
    Span4Mux_h I__1153 (
            .O(N__7478),
            .I(N__7467));
    Odrv12 I__1152 (
            .O(N__7475),
            .I(write_data_c_0));
    Odrv4 I__1151 (
            .O(N__7472),
            .I(write_data_c_0));
    Odrv4 I__1150 (
            .O(N__7467),
            .I(write_data_c_0));
    CascadeMux I__1149 (
            .O(N__7460),
            .I(N__7457));
    CascadeBuf I__1148 (
            .O(N__7457),
            .I(N__7454));
    CascadeMux I__1147 (
            .O(N__7454),
            .I(N__7451));
    CascadeBuf I__1146 (
            .O(N__7451),
            .I(N__7448));
    CascadeMux I__1145 (
            .O(N__7448),
            .I(N__7445));
    CascadeBuf I__1144 (
            .O(N__7445),
            .I(N__7442));
    CascadeMux I__1143 (
            .O(N__7442),
            .I(N__7438));
    CascadeMux I__1142 (
            .O(N__7441),
            .I(N__7435));
    CascadeBuf I__1141 (
            .O(N__7438),
            .I(N__7432));
    CascadeBuf I__1140 (
            .O(N__7435),
            .I(N__7429));
    CascadeMux I__1139 (
            .O(N__7432),
            .I(N__7426));
    CascadeMux I__1138 (
            .O(N__7429),
            .I(N__7423));
    CascadeBuf I__1137 (
            .O(N__7426),
            .I(N__7420));
    CascadeBuf I__1136 (
            .O(N__7423),
            .I(N__7417));
    CascadeMux I__1135 (
            .O(N__7420),
            .I(N__7414));
    CascadeMux I__1134 (
            .O(N__7417),
            .I(N__7411));
    CascadeBuf I__1133 (
            .O(N__7414),
            .I(N__7408));
    CascadeBuf I__1132 (
            .O(N__7411),
            .I(N__7405));
    CascadeMux I__1131 (
            .O(N__7408),
            .I(N__7402));
    CascadeMux I__1130 (
            .O(N__7405),
            .I(N__7399));
    CascadeBuf I__1129 (
            .O(N__7402),
            .I(N__7396));
    CascadeBuf I__1128 (
            .O(N__7399),
            .I(N__7393));
    CascadeMux I__1127 (
            .O(N__7396),
            .I(N__7390));
    CascadeMux I__1126 (
            .O(N__7393),
            .I(N__7387));
    CascadeBuf I__1125 (
            .O(N__7390),
            .I(N__7384));
    CascadeBuf I__1124 (
            .O(N__7387),
            .I(N__7381));
    CascadeMux I__1123 (
            .O(N__7384),
            .I(N__7378));
    CascadeMux I__1122 (
            .O(N__7381),
            .I(N__7375));
    CascadeBuf I__1121 (
            .O(N__7378),
            .I(N__7372));
    CascadeBuf I__1120 (
            .O(N__7375),
            .I(N__7369));
    CascadeMux I__1119 (
            .O(N__7372),
            .I(N__7366));
    CascadeMux I__1118 (
            .O(N__7369),
            .I(N__7363));
    CascadeBuf I__1117 (
            .O(N__7366),
            .I(N__7360));
    CascadeBuf I__1116 (
            .O(N__7363),
            .I(N__7357));
    CascadeMux I__1115 (
            .O(N__7360),
            .I(N__7354));
    CascadeMux I__1114 (
            .O(N__7357),
            .I(N__7351));
    CascadeBuf I__1113 (
            .O(N__7354),
            .I(N__7348));
    CascadeBuf I__1112 (
            .O(N__7351),
            .I(N__7345));
    CascadeMux I__1111 (
            .O(N__7348),
            .I(N__7342));
    CascadeMux I__1110 (
            .O(N__7345),
            .I(N__7339));
    CascadeBuf I__1109 (
            .O(N__7342),
            .I(N__7336));
    CascadeBuf I__1108 (
            .O(N__7339),
            .I(N__7333));
    CascadeMux I__1107 (
            .O(N__7336),
            .I(N__7330));
    CascadeMux I__1106 (
            .O(N__7333),
            .I(N__7327));
    CascadeBuf I__1105 (
            .O(N__7330),
            .I(N__7324));
    CascadeBuf I__1104 (
            .O(N__7327),
            .I(N__7321));
    CascadeMux I__1103 (
            .O(N__7324),
            .I(N__7318));
    CascadeMux I__1102 (
            .O(N__7321),
            .I(N__7315));
    CascadeBuf I__1101 (
            .O(N__7318),
            .I(N__7312));
    CascadeBuf I__1100 (
            .O(N__7315),
            .I(N__7309));
    CascadeMux I__1099 (
            .O(N__7312),
            .I(N__7306));
    CascadeMux I__1098 (
            .O(N__7309),
            .I(N__7303));
    CascadeBuf I__1097 (
            .O(N__7306),
            .I(N__7300));
    CascadeBuf I__1096 (
            .O(N__7303),
            .I(N__7297));
    CascadeMux I__1095 (
            .O(N__7300),
            .I(N__7294));
    CascadeMux I__1094 (
            .O(N__7297),
            .I(N__7291));
    InMux I__1093 (
            .O(N__7294),
            .I(N__7288));
    CascadeBuf I__1092 (
            .O(N__7291),
            .I(N__7285));
    LocalMux I__1091 (
            .O(N__7288),
            .I(N__7282));
    CascadeMux I__1090 (
            .O(N__7285),
            .I(N__7279));
    Span4Mux_s3_v I__1089 (
            .O(N__7282),
            .I(N__7276));
    InMux I__1088 (
            .O(N__7279),
            .I(N__7273));
    Span4Mux_h I__1087 (
            .O(N__7276),
            .I(N__7270));
    LocalMux I__1086 (
            .O(N__7273),
            .I(N__7267));
    Sp12to4 I__1085 (
            .O(N__7270),
            .I(N__7264));
    Span4Mux_v I__1084 (
            .O(N__7267),
            .I(N__7261));
    Span12Mux_h I__1083 (
            .O(N__7264),
            .I(N__7258));
    Odrv4 I__1082 (
            .O(N__7261),
            .I(write_address_c_9));
    Odrv12 I__1081 (
            .O(N__7258),
            .I(write_address_c_9));
    CascadeMux I__1080 (
            .O(N__7253),
            .I(N__7250));
    CascadeBuf I__1079 (
            .O(N__7250),
            .I(N__7247));
    CascadeMux I__1078 (
            .O(N__7247),
            .I(N__7244));
    CascadeBuf I__1077 (
            .O(N__7244),
            .I(N__7240));
    CascadeMux I__1076 (
            .O(N__7243),
            .I(N__7237));
    CascadeMux I__1075 (
            .O(N__7240),
            .I(N__7234));
    CascadeBuf I__1074 (
            .O(N__7237),
            .I(N__7231));
    CascadeBuf I__1073 (
            .O(N__7234),
            .I(N__7228));
    CascadeMux I__1072 (
            .O(N__7231),
            .I(N__7225));
    CascadeMux I__1071 (
            .O(N__7228),
            .I(N__7222));
    CascadeBuf I__1070 (
            .O(N__7225),
            .I(N__7219));
    CascadeBuf I__1069 (
            .O(N__7222),
            .I(N__7216));
    CascadeMux I__1068 (
            .O(N__7219),
            .I(N__7213));
    CascadeMux I__1067 (
            .O(N__7216),
            .I(N__7210));
    CascadeBuf I__1066 (
            .O(N__7213),
            .I(N__7207));
    CascadeBuf I__1065 (
            .O(N__7210),
            .I(N__7204));
    CascadeMux I__1064 (
            .O(N__7207),
            .I(N__7201));
    CascadeMux I__1063 (
            .O(N__7204),
            .I(N__7198));
    CascadeBuf I__1062 (
            .O(N__7201),
            .I(N__7195));
    CascadeBuf I__1061 (
            .O(N__7198),
            .I(N__7192));
    CascadeMux I__1060 (
            .O(N__7195),
            .I(N__7189));
    CascadeMux I__1059 (
            .O(N__7192),
            .I(N__7186));
    CascadeBuf I__1058 (
            .O(N__7189),
            .I(N__7183));
    CascadeBuf I__1057 (
            .O(N__7186),
            .I(N__7180));
    CascadeMux I__1056 (
            .O(N__7183),
            .I(N__7177));
    CascadeMux I__1055 (
            .O(N__7180),
            .I(N__7174));
    CascadeBuf I__1054 (
            .O(N__7177),
            .I(N__7171));
    CascadeBuf I__1053 (
            .O(N__7174),
            .I(N__7168));
    CascadeMux I__1052 (
            .O(N__7171),
            .I(N__7165));
    CascadeMux I__1051 (
            .O(N__7168),
            .I(N__7162));
    CascadeBuf I__1050 (
            .O(N__7165),
            .I(N__7159));
    CascadeBuf I__1049 (
            .O(N__7162),
            .I(N__7156));
    CascadeMux I__1048 (
            .O(N__7159),
            .I(N__7153));
    CascadeMux I__1047 (
            .O(N__7156),
            .I(N__7150));
    CascadeBuf I__1046 (
            .O(N__7153),
            .I(N__7147));
    CascadeBuf I__1045 (
            .O(N__7150),
            .I(N__7144));
    CascadeMux I__1044 (
            .O(N__7147),
            .I(N__7141));
    CascadeMux I__1043 (
            .O(N__7144),
            .I(N__7138));
    CascadeBuf I__1042 (
            .O(N__7141),
            .I(N__7135));
    CascadeBuf I__1041 (
            .O(N__7138),
            .I(N__7132));
    CascadeMux I__1040 (
            .O(N__7135),
            .I(N__7129));
    CascadeMux I__1039 (
            .O(N__7132),
            .I(N__7126));
    CascadeBuf I__1038 (
            .O(N__7129),
            .I(N__7123));
    CascadeBuf I__1037 (
            .O(N__7126),
            .I(N__7120));
    CascadeMux I__1036 (
            .O(N__7123),
            .I(N__7117));
    CascadeMux I__1035 (
            .O(N__7120),
            .I(N__7114));
    CascadeBuf I__1034 (
            .O(N__7117),
            .I(N__7111));
    CascadeBuf I__1033 (
            .O(N__7114),
            .I(N__7108));
    CascadeMux I__1032 (
            .O(N__7111),
            .I(N__7105));
    CascadeMux I__1031 (
            .O(N__7108),
            .I(N__7102));
    CascadeBuf I__1030 (
            .O(N__7105),
            .I(N__7099));
    CascadeBuf I__1029 (
            .O(N__7102),
            .I(N__7096));
    CascadeMux I__1028 (
            .O(N__7099),
            .I(N__7093));
    CascadeMux I__1027 (
            .O(N__7096),
            .I(N__7090));
    CascadeBuf I__1026 (
            .O(N__7093),
            .I(N__7087));
    CascadeBuf I__1025 (
            .O(N__7090),
            .I(N__7084));
    CascadeMux I__1024 (
            .O(N__7087),
            .I(N__7081));
    CascadeMux I__1023 (
            .O(N__7084),
            .I(N__7078));
    InMux I__1022 (
            .O(N__7081),
            .I(N__7075));
    InMux I__1021 (
            .O(N__7078),
            .I(N__7072));
    LocalMux I__1020 (
            .O(N__7075),
            .I(N__7069));
    LocalMux I__1019 (
            .O(N__7072),
            .I(N__7066));
    Span4Mux_v I__1018 (
            .O(N__7069),
            .I(N__7063));
    IoSpan4Mux I__1017 (
            .O(N__7066),
            .I(N__7060));
    IoSpan4Mux I__1016 (
            .O(N__7063),
            .I(N__7057));
    IoSpan4Mux I__1015 (
            .O(N__7060),
            .I(N__7054));
    IoSpan4Mux I__1014 (
            .O(N__7057),
            .I(N__7051));
    IoSpan4Mux I__1013 (
            .O(N__7054),
            .I(N__7048));
    Odrv4 I__1012 (
            .O(N__7051),
            .I(write_address_c_8));
    Odrv4 I__1011 (
            .O(N__7048),
            .I(write_address_c_8));
    CascadeMux I__1010 (
            .O(N__7043),
            .I(N__7040));
    CascadeBuf I__1009 (
            .O(N__7040),
            .I(N__7037));
    CascadeMux I__1008 (
            .O(N__7037),
            .I(N__7034));
    CascadeBuf I__1007 (
            .O(N__7034),
            .I(N__7031));
    CascadeMux I__1006 (
            .O(N__7031),
            .I(N__7027));
    CascadeMux I__1005 (
            .O(N__7030),
            .I(N__7024));
    CascadeBuf I__1004 (
            .O(N__7027),
            .I(N__7021));
    CascadeBuf I__1003 (
            .O(N__7024),
            .I(N__7018));
    CascadeMux I__1002 (
            .O(N__7021),
            .I(N__7015));
    CascadeMux I__1001 (
            .O(N__7018),
            .I(N__7012));
    CascadeBuf I__1000 (
            .O(N__7015),
            .I(N__7009));
    CascadeBuf I__999 (
            .O(N__7012),
            .I(N__7006));
    CascadeMux I__998 (
            .O(N__7009),
            .I(N__7003));
    CascadeMux I__997 (
            .O(N__7006),
            .I(N__7000));
    CascadeBuf I__996 (
            .O(N__7003),
            .I(N__6997));
    CascadeBuf I__995 (
            .O(N__7000),
            .I(N__6994));
    CascadeMux I__994 (
            .O(N__6997),
            .I(N__6991));
    CascadeMux I__993 (
            .O(N__6994),
            .I(N__6988));
    CascadeBuf I__992 (
            .O(N__6991),
            .I(N__6985));
    CascadeBuf I__991 (
            .O(N__6988),
            .I(N__6982));
    CascadeMux I__990 (
            .O(N__6985),
            .I(N__6979));
    CascadeMux I__989 (
            .O(N__6982),
            .I(N__6976));
    CascadeBuf I__988 (
            .O(N__6979),
            .I(N__6973));
    CascadeBuf I__987 (
            .O(N__6976),
            .I(N__6970));
    CascadeMux I__986 (
            .O(N__6973),
            .I(N__6967));
    CascadeMux I__985 (
            .O(N__6970),
            .I(N__6964));
    CascadeBuf I__984 (
            .O(N__6967),
            .I(N__6961));
    CascadeBuf I__983 (
            .O(N__6964),
            .I(N__6958));
    CascadeMux I__982 (
            .O(N__6961),
            .I(N__6955));
    CascadeMux I__981 (
            .O(N__6958),
            .I(N__6952));
    CascadeBuf I__980 (
            .O(N__6955),
            .I(N__6949));
    CascadeBuf I__979 (
            .O(N__6952),
            .I(N__6946));
    CascadeMux I__978 (
            .O(N__6949),
            .I(N__6943));
    CascadeMux I__977 (
            .O(N__6946),
            .I(N__6940));
    CascadeBuf I__976 (
            .O(N__6943),
            .I(N__6937));
    CascadeBuf I__975 (
            .O(N__6940),
            .I(N__6934));
    CascadeMux I__974 (
            .O(N__6937),
            .I(N__6931));
    CascadeMux I__973 (
            .O(N__6934),
            .I(N__6928));
    CascadeBuf I__972 (
            .O(N__6931),
            .I(N__6925));
    CascadeBuf I__971 (
            .O(N__6928),
            .I(N__6922));
    CascadeMux I__970 (
            .O(N__6925),
            .I(N__6919));
    CascadeMux I__969 (
            .O(N__6922),
            .I(N__6916));
    CascadeBuf I__968 (
            .O(N__6919),
            .I(N__6913));
    CascadeBuf I__967 (
            .O(N__6916),
            .I(N__6910));
    CascadeMux I__966 (
            .O(N__6913),
            .I(N__6907));
    CascadeMux I__965 (
            .O(N__6910),
            .I(N__6904));
    CascadeBuf I__964 (
            .O(N__6907),
            .I(N__6901));
    CascadeBuf I__963 (
            .O(N__6904),
            .I(N__6898));
    CascadeMux I__962 (
            .O(N__6901),
            .I(N__6895));
    CascadeMux I__961 (
            .O(N__6898),
            .I(N__6892));
    CascadeBuf I__960 (
            .O(N__6895),
            .I(N__6889));
    CascadeBuf I__959 (
            .O(N__6892),
            .I(N__6886));
    CascadeMux I__958 (
            .O(N__6889),
            .I(N__6883));
    CascadeMux I__957 (
            .O(N__6886),
            .I(N__6880));
    CascadeBuf I__956 (
            .O(N__6883),
            .I(N__6877));
    CascadeBuf I__955 (
            .O(N__6880),
            .I(N__6874));
    CascadeMux I__954 (
            .O(N__6877),
            .I(N__6871));
    CascadeMux I__953 (
            .O(N__6874),
            .I(N__6868));
    InMux I__952 (
            .O(N__6871),
            .I(N__6865));
    InMux I__951 (
            .O(N__6868),
            .I(N__6862));
    LocalMux I__950 (
            .O(N__6865),
            .I(N__6859));
    LocalMux I__949 (
            .O(N__6862),
            .I(N__6856));
    Span4Mux_s2_v I__948 (
            .O(N__6859),
            .I(N__6853));
    Span4Mux_h I__947 (
            .O(N__6856),
            .I(N__6850));
    Sp12to4 I__946 (
            .O(N__6853),
            .I(N__6847));
    Sp12to4 I__945 (
            .O(N__6850),
            .I(N__6842));
    Span12Mux_h I__944 (
            .O(N__6847),
            .I(N__6842));
    Span12Mux_v I__943 (
            .O(N__6842),
            .I(N__6839));
    Span12Mux_v I__942 (
            .O(N__6839),
            .I(N__6836));
    Odrv12 I__941 (
            .O(N__6836),
            .I(write_address_c_7));
    CascadeMux I__940 (
            .O(N__6833),
            .I(N__6830));
    CascadeBuf I__939 (
            .O(N__6830),
            .I(N__6827));
    CascadeMux I__938 (
            .O(N__6827),
            .I(N__6824));
    CascadeBuf I__937 (
            .O(N__6824),
            .I(N__6821));
    CascadeMux I__936 (
            .O(N__6821),
            .I(N__6818));
    CascadeBuf I__935 (
            .O(N__6818),
            .I(N__6815));
    CascadeMux I__934 (
            .O(N__6815),
            .I(N__6811));
    CascadeMux I__933 (
            .O(N__6814),
            .I(N__6808));
    CascadeBuf I__932 (
            .O(N__6811),
            .I(N__6805));
    CascadeBuf I__931 (
            .O(N__6808),
            .I(N__6802));
    CascadeMux I__930 (
            .O(N__6805),
            .I(N__6799));
    CascadeMux I__929 (
            .O(N__6802),
            .I(N__6796));
    CascadeBuf I__928 (
            .O(N__6799),
            .I(N__6793));
    CascadeBuf I__927 (
            .O(N__6796),
            .I(N__6790));
    CascadeMux I__926 (
            .O(N__6793),
            .I(N__6787));
    CascadeMux I__925 (
            .O(N__6790),
            .I(N__6784));
    CascadeBuf I__924 (
            .O(N__6787),
            .I(N__6781));
    CascadeBuf I__923 (
            .O(N__6784),
            .I(N__6778));
    CascadeMux I__922 (
            .O(N__6781),
            .I(N__6775));
    CascadeMux I__921 (
            .O(N__6778),
            .I(N__6772));
    CascadeBuf I__920 (
            .O(N__6775),
            .I(N__6769));
    CascadeBuf I__919 (
            .O(N__6772),
            .I(N__6766));
    CascadeMux I__918 (
            .O(N__6769),
            .I(N__6763));
    CascadeMux I__917 (
            .O(N__6766),
            .I(N__6760));
    CascadeBuf I__916 (
            .O(N__6763),
            .I(N__6757));
    CascadeBuf I__915 (
            .O(N__6760),
            .I(N__6754));
    CascadeMux I__914 (
            .O(N__6757),
            .I(N__6751));
    CascadeMux I__913 (
            .O(N__6754),
            .I(N__6748));
    CascadeBuf I__912 (
            .O(N__6751),
            .I(N__6745));
    CascadeBuf I__911 (
            .O(N__6748),
            .I(N__6742));
    CascadeMux I__910 (
            .O(N__6745),
            .I(N__6739));
    CascadeMux I__909 (
            .O(N__6742),
            .I(N__6736));
    CascadeBuf I__908 (
            .O(N__6739),
            .I(N__6733));
    CascadeBuf I__907 (
            .O(N__6736),
            .I(N__6730));
    CascadeMux I__906 (
            .O(N__6733),
            .I(N__6727));
    CascadeMux I__905 (
            .O(N__6730),
            .I(N__6724));
    CascadeBuf I__904 (
            .O(N__6727),
            .I(N__6721));
    CascadeBuf I__903 (
            .O(N__6724),
            .I(N__6718));
    CascadeMux I__902 (
            .O(N__6721),
            .I(N__6715));
    CascadeMux I__901 (
            .O(N__6718),
            .I(N__6712));
    CascadeBuf I__900 (
            .O(N__6715),
            .I(N__6709));
    CascadeBuf I__899 (
            .O(N__6712),
            .I(N__6706));
    CascadeMux I__898 (
            .O(N__6709),
            .I(N__6703));
    CascadeMux I__897 (
            .O(N__6706),
            .I(N__6700));
    CascadeBuf I__896 (
            .O(N__6703),
            .I(N__6697));
    CascadeBuf I__895 (
            .O(N__6700),
            .I(N__6694));
    CascadeMux I__894 (
            .O(N__6697),
            .I(N__6691));
    CascadeMux I__893 (
            .O(N__6694),
            .I(N__6688));
    CascadeBuf I__892 (
            .O(N__6691),
            .I(N__6685));
    CascadeBuf I__891 (
            .O(N__6688),
            .I(N__6682));
    CascadeMux I__890 (
            .O(N__6685),
            .I(N__6679));
    CascadeMux I__889 (
            .O(N__6682),
            .I(N__6676));
    CascadeBuf I__888 (
            .O(N__6679),
            .I(N__6673));
    CascadeBuf I__887 (
            .O(N__6676),
            .I(N__6670));
    CascadeMux I__886 (
            .O(N__6673),
            .I(N__6667));
    CascadeMux I__885 (
            .O(N__6670),
            .I(N__6664));
    InMux I__884 (
            .O(N__6667),
            .I(N__6661));
    CascadeBuf I__883 (
            .O(N__6664),
            .I(N__6658));
    LocalMux I__882 (
            .O(N__6661),
            .I(N__6655));
    CascadeMux I__881 (
            .O(N__6658),
            .I(N__6652));
    Span4Mux_v I__880 (
            .O(N__6655),
            .I(N__6649));
    InMux I__879 (
            .O(N__6652),
            .I(N__6646));
    Sp12to4 I__878 (
            .O(N__6649),
            .I(N__6643));
    LocalMux I__877 (
            .O(N__6646),
            .I(N__6640));
    Span12Mux_h I__876 (
            .O(N__6643),
            .I(N__6637));
    Span12Mux_h I__875 (
            .O(N__6640),
            .I(N__6634));
    Span12Mux_v I__874 (
            .O(N__6637),
            .I(N__6631));
    Span12Mux_v I__873 (
            .O(N__6634),
            .I(N__6626));
    Span12Mux_h I__872 (
            .O(N__6631),
            .I(N__6626));
    Odrv12 I__871 (
            .O(N__6626),
            .I(write_address_c_6));
    CascadeMux I__870 (
            .O(N__6623),
            .I(N__6620));
    CascadeBuf I__869 (
            .O(N__6620),
            .I(N__6617));
    CascadeMux I__868 (
            .O(N__6617),
            .I(N__6614));
    CascadeBuf I__867 (
            .O(N__6614),
            .I(N__6611));
    CascadeMux I__866 (
            .O(N__6611),
            .I(N__6608));
    CascadeBuf I__865 (
            .O(N__6608),
            .I(N__6605));
    CascadeMux I__864 (
            .O(N__6605),
            .I(N__6601));
    CascadeMux I__863 (
            .O(N__6604),
            .I(N__6598));
    CascadeBuf I__862 (
            .O(N__6601),
            .I(N__6595));
    CascadeBuf I__861 (
            .O(N__6598),
            .I(N__6592));
    CascadeMux I__860 (
            .O(N__6595),
            .I(N__6589));
    CascadeMux I__859 (
            .O(N__6592),
            .I(N__6586));
    CascadeBuf I__858 (
            .O(N__6589),
            .I(N__6583));
    CascadeBuf I__857 (
            .O(N__6586),
            .I(N__6580));
    CascadeMux I__856 (
            .O(N__6583),
            .I(N__6577));
    CascadeMux I__855 (
            .O(N__6580),
            .I(N__6574));
    CascadeBuf I__854 (
            .O(N__6577),
            .I(N__6571));
    CascadeBuf I__853 (
            .O(N__6574),
            .I(N__6568));
    CascadeMux I__852 (
            .O(N__6571),
            .I(N__6565));
    CascadeMux I__851 (
            .O(N__6568),
            .I(N__6562));
    CascadeBuf I__850 (
            .O(N__6565),
            .I(N__6559));
    CascadeBuf I__849 (
            .O(N__6562),
            .I(N__6556));
    CascadeMux I__848 (
            .O(N__6559),
            .I(N__6553));
    CascadeMux I__847 (
            .O(N__6556),
            .I(N__6550));
    CascadeBuf I__846 (
            .O(N__6553),
            .I(N__6547));
    CascadeBuf I__845 (
            .O(N__6550),
            .I(N__6544));
    CascadeMux I__844 (
            .O(N__6547),
            .I(N__6541));
    CascadeMux I__843 (
            .O(N__6544),
            .I(N__6538));
    CascadeBuf I__842 (
            .O(N__6541),
            .I(N__6535));
    CascadeBuf I__841 (
            .O(N__6538),
            .I(N__6532));
    CascadeMux I__840 (
            .O(N__6535),
            .I(N__6529));
    CascadeMux I__839 (
            .O(N__6532),
            .I(N__6526));
    CascadeBuf I__838 (
            .O(N__6529),
            .I(N__6523));
    CascadeBuf I__837 (
            .O(N__6526),
            .I(N__6520));
    CascadeMux I__836 (
            .O(N__6523),
            .I(N__6517));
    CascadeMux I__835 (
            .O(N__6520),
            .I(N__6514));
    CascadeBuf I__834 (
            .O(N__6517),
            .I(N__6511));
    CascadeBuf I__833 (
            .O(N__6514),
            .I(N__6508));
    CascadeMux I__832 (
            .O(N__6511),
            .I(N__6505));
    CascadeMux I__831 (
            .O(N__6508),
            .I(N__6502));
    CascadeBuf I__830 (
            .O(N__6505),
            .I(N__6499));
    CascadeBuf I__829 (
            .O(N__6502),
            .I(N__6496));
    CascadeMux I__828 (
            .O(N__6499),
            .I(N__6493));
    CascadeMux I__827 (
            .O(N__6496),
            .I(N__6490));
    CascadeBuf I__826 (
            .O(N__6493),
            .I(N__6487));
    CascadeBuf I__825 (
            .O(N__6490),
            .I(N__6484));
    CascadeMux I__824 (
            .O(N__6487),
            .I(N__6481));
    CascadeMux I__823 (
            .O(N__6484),
            .I(N__6478));
    CascadeBuf I__822 (
            .O(N__6481),
            .I(N__6475));
    CascadeBuf I__821 (
            .O(N__6478),
            .I(N__6472));
    CascadeMux I__820 (
            .O(N__6475),
            .I(N__6469));
    CascadeMux I__819 (
            .O(N__6472),
            .I(N__6466));
    CascadeBuf I__818 (
            .O(N__6469),
            .I(N__6463));
    CascadeBuf I__817 (
            .O(N__6466),
            .I(N__6460));
    CascadeMux I__816 (
            .O(N__6463),
            .I(N__6457));
    CascadeMux I__815 (
            .O(N__6460),
            .I(N__6454));
    InMux I__814 (
            .O(N__6457),
            .I(N__6451));
    CascadeBuf I__813 (
            .O(N__6454),
            .I(N__6448));
    LocalMux I__812 (
            .O(N__6451),
            .I(N__6445));
    CascadeMux I__811 (
            .O(N__6448),
            .I(N__6442));
    Span4Mux_s3_v I__810 (
            .O(N__6445),
            .I(N__6439));
    InMux I__809 (
            .O(N__6442),
            .I(N__6436));
    Span4Mux_v I__808 (
            .O(N__6439),
            .I(N__6433));
    LocalMux I__807 (
            .O(N__6436),
            .I(N__6430));
    Span4Mux_v I__806 (
            .O(N__6433),
            .I(N__6427));
    Sp12to4 I__805 (
            .O(N__6430),
            .I(N__6424));
    Sp12to4 I__804 (
            .O(N__6427),
            .I(N__6421));
    Span12Mux_s11_v I__803 (
            .O(N__6424),
            .I(N__6418));
    Span12Mux_h I__802 (
            .O(N__6421),
            .I(N__6415));
    Odrv12 I__801 (
            .O(N__6418),
            .I(write_address_c_5));
    Odrv12 I__800 (
            .O(N__6415),
            .I(write_address_c_5));
    CascadeMux I__799 (
            .O(N__6410),
            .I(N__6407));
    CascadeBuf I__798 (
            .O(N__6407),
            .I(N__6404));
    CascadeMux I__797 (
            .O(N__6404),
            .I(N__6401));
    CascadeBuf I__796 (
            .O(N__6401),
            .I(N__6398));
    CascadeMux I__795 (
            .O(N__6398),
            .I(N__6395));
    CascadeBuf I__794 (
            .O(N__6395),
            .I(N__6391));
    CascadeMux I__793 (
            .O(N__6394),
            .I(N__6388));
    CascadeMux I__792 (
            .O(N__6391),
            .I(N__6385));
    CascadeBuf I__791 (
            .O(N__6388),
            .I(N__6382));
    CascadeBuf I__790 (
            .O(N__6385),
            .I(N__6379));
    CascadeMux I__789 (
            .O(N__6382),
            .I(N__6376));
    CascadeMux I__788 (
            .O(N__6379),
            .I(N__6373));
    CascadeBuf I__787 (
            .O(N__6376),
            .I(N__6370));
    CascadeBuf I__786 (
            .O(N__6373),
            .I(N__6367));
    CascadeMux I__785 (
            .O(N__6370),
            .I(N__6364));
    CascadeMux I__784 (
            .O(N__6367),
            .I(N__6361));
    CascadeBuf I__783 (
            .O(N__6364),
            .I(N__6358));
    CascadeBuf I__782 (
            .O(N__6361),
            .I(N__6355));
    CascadeMux I__781 (
            .O(N__6358),
            .I(N__6352));
    CascadeMux I__780 (
            .O(N__6355),
            .I(N__6349));
    CascadeBuf I__779 (
            .O(N__6352),
            .I(N__6346));
    CascadeBuf I__778 (
            .O(N__6349),
            .I(N__6343));
    CascadeMux I__777 (
            .O(N__6346),
            .I(N__6340));
    CascadeMux I__776 (
            .O(N__6343),
            .I(N__6337));
    CascadeBuf I__775 (
            .O(N__6340),
            .I(N__6334));
    CascadeBuf I__774 (
            .O(N__6337),
            .I(N__6331));
    CascadeMux I__773 (
            .O(N__6334),
            .I(N__6328));
    CascadeMux I__772 (
            .O(N__6331),
            .I(N__6325));
    CascadeBuf I__771 (
            .O(N__6328),
            .I(N__6322));
    CascadeBuf I__770 (
            .O(N__6325),
            .I(N__6319));
    CascadeMux I__769 (
            .O(N__6322),
            .I(N__6316));
    CascadeMux I__768 (
            .O(N__6319),
            .I(N__6313));
    CascadeBuf I__767 (
            .O(N__6316),
            .I(N__6310));
    CascadeBuf I__766 (
            .O(N__6313),
            .I(N__6307));
    CascadeMux I__765 (
            .O(N__6310),
            .I(N__6304));
    CascadeMux I__764 (
            .O(N__6307),
            .I(N__6301));
    CascadeBuf I__763 (
            .O(N__6304),
            .I(N__6298));
    CascadeBuf I__762 (
            .O(N__6301),
            .I(N__6295));
    CascadeMux I__761 (
            .O(N__6298),
            .I(N__6292));
    CascadeMux I__760 (
            .O(N__6295),
            .I(N__6289));
    CascadeBuf I__759 (
            .O(N__6292),
            .I(N__6286));
    CascadeBuf I__758 (
            .O(N__6289),
            .I(N__6283));
    CascadeMux I__757 (
            .O(N__6286),
            .I(N__6280));
    CascadeMux I__756 (
            .O(N__6283),
            .I(N__6277));
    CascadeBuf I__755 (
            .O(N__6280),
            .I(N__6274));
    CascadeBuf I__754 (
            .O(N__6277),
            .I(N__6271));
    CascadeMux I__753 (
            .O(N__6274),
            .I(N__6268));
    CascadeMux I__752 (
            .O(N__6271),
            .I(N__6265));
    CascadeBuf I__751 (
            .O(N__6268),
            .I(N__6262));
    CascadeBuf I__750 (
            .O(N__6265),
            .I(N__6259));
    CascadeMux I__749 (
            .O(N__6262),
            .I(N__6256));
    CascadeMux I__748 (
            .O(N__6259),
            .I(N__6253));
    CascadeBuf I__747 (
            .O(N__6256),
            .I(N__6250));
    CascadeBuf I__746 (
            .O(N__6253),
            .I(N__6247));
    CascadeMux I__745 (
            .O(N__6250),
            .I(N__6244));
    CascadeMux I__744 (
            .O(N__6247),
            .I(N__6241));
    CascadeBuf I__743 (
            .O(N__6244),
            .I(N__6238));
    InMux I__742 (
            .O(N__6241),
            .I(N__6235));
    CascadeMux I__741 (
            .O(N__6238),
            .I(N__6232));
    LocalMux I__740 (
            .O(N__6235),
            .I(N__6229));
    InMux I__739 (
            .O(N__6232),
            .I(N__6226));
    Span4Mux_v I__738 (
            .O(N__6229),
            .I(N__6223));
    LocalMux I__737 (
            .O(N__6226),
            .I(N__6220));
    Span4Mux_v I__736 (
            .O(N__6223),
            .I(N__6217));
    Span4Mux_v I__735 (
            .O(N__6220),
            .I(N__6214));
    Sp12to4 I__734 (
            .O(N__6217),
            .I(N__6211));
    Sp12to4 I__733 (
            .O(N__6214),
            .I(N__6206));
    Span12Mux_h I__732 (
            .O(N__6211),
            .I(N__6206));
    Odrv12 I__731 (
            .O(N__6206),
            .I(write_address_c_4));
    CascadeMux I__730 (
            .O(N__6203),
            .I(N__6200));
    CascadeBuf I__729 (
            .O(N__6200),
            .I(N__6197));
    CascadeMux I__728 (
            .O(N__6197),
            .I(N__6194));
    CascadeBuf I__727 (
            .O(N__6194),
            .I(N__6191));
    CascadeMux I__726 (
            .O(N__6191),
            .I(N__6188));
    CascadeBuf I__725 (
            .O(N__6188),
            .I(N__6184));
    CascadeMux I__724 (
            .O(N__6187),
            .I(N__6181));
    CascadeMux I__723 (
            .O(N__6184),
            .I(N__6178));
    CascadeBuf I__722 (
            .O(N__6181),
            .I(N__6175));
    CascadeBuf I__721 (
            .O(N__6178),
            .I(N__6172));
    CascadeMux I__720 (
            .O(N__6175),
            .I(N__6169));
    CascadeMux I__719 (
            .O(N__6172),
            .I(N__6166));
    CascadeBuf I__718 (
            .O(N__6169),
            .I(N__6163));
    CascadeBuf I__717 (
            .O(N__6166),
            .I(N__6160));
    CascadeMux I__716 (
            .O(N__6163),
            .I(N__6157));
    CascadeMux I__715 (
            .O(N__6160),
            .I(N__6154));
    CascadeBuf I__714 (
            .O(N__6157),
            .I(N__6151));
    CascadeBuf I__713 (
            .O(N__6154),
            .I(N__6148));
    CascadeMux I__712 (
            .O(N__6151),
            .I(N__6145));
    CascadeMux I__711 (
            .O(N__6148),
            .I(N__6142));
    CascadeBuf I__710 (
            .O(N__6145),
            .I(N__6139));
    CascadeBuf I__709 (
            .O(N__6142),
            .I(N__6136));
    CascadeMux I__708 (
            .O(N__6139),
            .I(N__6133));
    CascadeMux I__707 (
            .O(N__6136),
            .I(N__6130));
    CascadeBuf I__706 (
            .O(N__6133),
            .I(N__6127));
    CascadeBuf I__705 (
            .O(N__6130),
            .I(N__6124));
    CascadeMux I__704 (
            .O(N__6127),
            .I(N__6121));
    CascadeMux I__703 (
            .O(N__6124),
            .I(N__6118));
    CascadeBuf I__702 (
            .O(N__6121),
            .I(N__6115));
    CascadeBuf I__701 (
            .O(N__6118),
            .I(N__6112));
    CascadeMux I__700 (
            .O(N__6115),
            .I(N__6109));
    CascadeMux I__699 (
            .O(N__6112),
            .I(N__6106));
    CascadeBuf I__698 (
            .O(N__6109),
            .I(N__6103));
    CascadeBuf I__697 (
            .O(N__6106),
            .I(N__6100));
    CascadeMux I__696 (
            .O(N__6103),
            .I(N__6097));
    CascadeMux I__695 (
            .O(N__6100),
            .I(N__6094));
    CascadeBuf I__694 (
            .O(N__6097),
            .I(N__6091));
    CascadeBuf I__693 (
            .O(N__6094),
            .I(N__6088));
    CascadeMux I__692 (
            .O(N__6091),
            .I(N__6085));
    CascadeMux I__691 (
            .O(N__6088),
            .I(N__6082));
    CascadeBuf I__690 (
            .O(N__6085),
            .I(N__6079));
    CascadeBuf I__689 (
            .O(N__6082),
            .I(N__6076));
    CascadeMux I__688 (
            .O(N__6079),
            .I(N__6073));
    CascadeMux I__687 (
            .O(N__6076),
            .I(N__6070));
    CascadeBuf I__686 (
            .O(N__6073),
            .I(N__6067));
    CascadeBuf I__685 (
            .O(N__6070),
            .I(N__6064));
    CascadeMux I__684 (
            .O(N__6067),
            .I(N__6061));
    CascadeMux I__683 (
            .O(N__6064),
            .I(N__6058));
    CascadeBuf I__682 (
            .O(N__6061),
            .I(N__6055));
    CascadeBuf I__681 (
            .O(N__6058),
            .I(N__6052));
    CascadeMux I__680 (
            .O(N__6055),
            .I(N__6049));
    CascadeMux I__679 (
            .O(N__6052),
            .I(N__6046));
    CascadeBuf I__678 (
            .O(N__6049),
            .I(N__6043));
    CascadeBuf I__677 (
            .O(N__6046),
            .I(N__6040));
    CascadeMux I__676 (
            .O(N__6043),
            .I(N__6037));
    CascadeMux I__675 (
            .O(N__6040),
            .I(N__6034));
    CascadeBuf I__674 (
            .O(N__6037),
            .I(N__6031));
    InMux I__673 (
            .O(N__6034),
            .I(N__6028));
    CascadeMux I__672 (
            .O(N__6031),
            .I(N__6025));
    LocalMux I__671 (
            .O(N__6028),
            .I(N__6022));
    InMux I__670 (
            .O(N__6025),
            .I(N__6019));
    Span4Mux_s1_v I__669 (
            .O(N__6022),
            .I(N__6016));
    LocalMux I__668 (
            .O(N__6019),
            .I(N__6013));
    Sp12to4 I__667 (
            .O(N__6016),
            .I(N__6010));
    Span4Mux_v I__666 (
            .O(N__6013),
            .I(N__6007));
    Span12Mux_h I__665 (
            .O(N__6010),
            .I(N__6004));
    Span4Mux_h I__664 (
            .O(N__6007),
            .I(N__6001));
    Span12Mux_h I__663 (
            .O(N__6004),
            .I(N__5998));
    Odrv4 I__662 (
            .O(N__6001),
            .I(write_address_c_3));
    Odrv12 I__661 (
            .O(N__5998),
            .I(write_address_c_3));
    CascadeMux I__660 (
            .O(N__5993),
            .I(N__5990));
    CascadeBuf I__659 (
            .O(N__5990),
            .I(N__5987));
    CascadeMux I__658 (
            .O(N__5987),
            .I(N__5983));
    CascadeMux I__657 (
            .O(N__5986),
            .I(N__5980));
    CascadeBuf I__656 (
            .O(N__5983),
            .I(N__5977));
    CascadeBuf I__655 (
            .O(N__5980),
            .I(N__5974));
    CascadeMux I__654 (
            .O(N__5977),
            .I(N__5971));
    CascadeMux I__653 (
            .O(N__5974),
            .I(N__5968));
    CascadeBuf I__652 (
            .O(N__5971),
            .I(N__5965));
    CascadeBuf I__651 (
            .O(N__5968),
            .I(N__5962));
    CascadeMux I__650 (
            .O(N__5965),
            .I(N__5959));
    CascadeMux I__649 (
            .O(N__5962),
            .I(N__5956));
    CascadeBuf I__648 (
            .O(N__5959),
            .I(N__5953));
    CascadeBuf I__647 (
            .O(N__5956),
            .I(N__5950));
    CascadeMux I__646 (
            .O(N__5953),
            .I(N__5947));
    CascadeMux I__645 (
            .O(N__5950),
            .I(N__5944));
    CascadeBuf I__644 (
            .O(N__5947),
            .I(N__5941));
    CascadeBuf I__643 (
            .O(N__5944),
            .I(N__5938));
    CascadeMux I__642 (
            .O(N__5941),
            .I(N__5935));
    CascadeMux I__641 (
            .O(N__5938),
            .I(N__5932));
    CascadeBuf I__640 (
            .O(N__5935),
            .I(N__5929));
    CascadeBuf I__639 (
            .O(N__5932),
            .I(N__5926));
    CascadeMux I__638 (
            .O(N__5929),
            .I(N__5923));
    CascadeMux I__637 (
            .O(N__5926),
            .I(N__5920));
    CascadeBuf I__636 (
            .O(N__5923),
            .I(N__5917));
    CascadeBuf I__635 (
            .O(N__5920),
            .I(N__5914));
    CascadeMux I__634 (
            .O(N__5917),
            .I(N__5911));
    CascadeMux I__633 (
            .O(N__5914),
            .I(N__5908));
    CascadeBuf I__632 (
            .O(N__5911),
            .I(N__5905));
    CascadeBuf I__631 (
            .O(N__5908),
            .I(N__5902));
    CascadeMux I__630 (
            .O(N__5905),
            .I(N__5899));
    CascadeMux I__629 (
            .O(N__5902),
            .I(N__5896));
    CascadeBuf I__628 (
            .O(N__5899),
            .I(N__5893));
    CascadeBuf I__627 (
            .O(N__5896),
            .I(N__5890));
    CascadeMux I__626 (
            .O(N__5893),
            .I(N__5887));
    CascadeMux I__625 (
            .O(N__5890),
            .I(N__5884));
    CascadeBuf I__624 (
            .O(N__5887),
            .I(N__5881));
    CascadeBuf I__623 (
            .O(N__5884),
            .I(N__5878));
    CascadeMux I__622 (
            .O(N__5881),
            .I(N__5875));
    CascadeMux I__621 (
            .O(N__5878),
            .I(N__5872));
    CascadeBuf I__620 (
            .O(N__5875),
            .I(N__5869));
    CascadeBuf I__619 (
            .O(N__5872),
            .I(N__5866));
    CascadeMux I__618 (
            .O(N__5869),
            .I(N__5863));
    CascadeMux I__617 (
            .O(N__5866),
            .I(N__5860));
    CascadeBuf I__616 (
            .O(N__5863),
            .I(N__5857));
    CascadeBuf I__615 (
            .O(N__5860),
            .I(N__5854));
    CascadeMux I__614 (
            .O(N__5857),
            .I(N__5851));
    CascadeMux I__613 (
            .O(N__5854),
            .I(N__5848));
    CascadeBuf I__612 (
            .O(N__5851),
            .I(N__5845));
    CascadeBuf I__611 (
            .O(N__5848),
            .I(N__5842));
    CascadeMux I__610 (
            .O(N__5845),
            .I(N__5839));
    CascadeMux I__609 (
            .O(N__5842),
            .I(N__5836));
    CascadeBuf I__608 (
            .O(N__5839),
            .I(N__5833));
    CascadeBuf I__607 (
            .O(N__5836),
            .I(N__5830));
    CascadeMux I__606 (
            .O(N__5833),
            .I(N__5827));
    CascadeMux I__605 (
            .O(N__5830),
            .I(N__5824));
    CascadeBuf I__604 (
            .O(N__5827),
            .I(N__5821));
    InMux I__603 (
            .O(N__5824),
            .I(N__5818));
    CascadeMux I__602 (
            .O(N__5821),
            .I(N__5815));
    LocalMux I__601 (
            .O(N__5818),
            .I(N__5812));
    InMux I__600 (
            .O(N__5815),
            .I(N__5809));
    Span4Mux_v I__599 (
            .O(N__5812),
            .I(N__5806));
    LocalMux I__598 (
            .O(N__5809),
            .I(N__5803));
    Sp12to4 I__597 (
            .O(N__5806),
            .I(N__5800));
    Span12Mux_s1_v I__596 (
            .O(N__5803),
            .I(N__5797));
    Span12Mux_h I__595 (
            .O(N__5800),
            .I(N__5792));
    Span12Mux_h I__594 (
            .O(N__5797),
            .I(N__5792));
    Odrv12 I__593 (
            .O(N__5792),
            .I(write_address_c_2));
    CascadeMux I__592 (
            .O(N__5789),
            .I(N__5786));
    CascadeBuf I__591 (
            .O(N__5786),
            .I(N__5783));
    CascadeMux I__590 (
            .O(N__5783),
            .I(N__5780));
    CascadeBuf I__589 (
            .O(N__5780),
            .I(N__5777));
    CascadeMux I__588 (
            .O(N__5777),
            .I(N__5773));
    CascadeMux I__587 (
            .O(N__5776),
            .I(N__5770));
    CascadeBuf I__586 (
            .O(N__5773),
            .I(N__5767));
    CascadeBuf I__585 (
            .O(N__5770),
            .I(N__5764));
    CascadeMux I__584 (
            .O(N__5767),
            .I(N__5761));
    CascadeMux I__583 (
            .O(N__5764),
            .I(N__5758));
    CascadeBuf I__582 (
            .O(N__5761),
            .I(N__5755));
    CascadeBuf I__581 (
            .O(N__5758),
            .I(N__5752));
    CascadeMux I__580 (
            .O(N__5755),
            .I(N__5749));
    CascadeMux I__579 (
            .O(N__5752),
            .I(N__5746));
    CascadeBuf I__578 (
            .O(N__5749),
            .I(N__5743));
    CascadeBuf I__577 (
            .O(N__5746),
            .I(N__5740));
    CascadeMux I__576 (
            .O(N__5743),
            .I(N__5737));
    CascadeMux I__575 (
            .O(N__5740),
            .I(N__5734));
    CascadeBuf I__574 (
            .O(N__5737),
            .I(N__5731));
    CascadeBuf I__573 (
            .O(N__5734),
            .I(N__5728));
    CascadeMux I__572 (
            .O(N__5731),
            .I(N__5725));
    CascadeMux I__571 (
            .O(N__5728),
            .I(N__5722));
    CascadeBuf I__570 (
            .O(N__5725),
            .I(N__5719));
    CascadeBuf I__569 (
            .O(N__5722),
            .I(N__5716));
    CascadeMux I__568 (
            .O(N__5719),
            .I(N__5713));
    CascadeMux I__567 (
            .O(N__5716),
            .I(N__5710));
    CascadeBuf I__566 (
            .O(N__5713),
            .I(N__5707));
    CascadeBuf I__565 (
            .O(N__5710),
            .I(N__5704));
    CascadeMux I__564 (
            .O(N__5707),
            .I(N__5701));
    CascadeMux I__563 (
            .O(N__5704),
            .I(N__5698));
    CascadeBuf I__562 (
            .O(N__5701),
            .I(N__5695));
    CascadeBuf I__561 (
            .O(N__5698),
            .I(N__5692));
    CascadeMux I__560 (
            .O(N__5695),
            .I(N__5689));
    CascadeMux I__559 (
            .O(N__5692),
            .I(N__5686));
    CascadeBuf I__558 (
            .O(N__5689),
            .I(N__5683));
    CascadeBuf I__557 (
            .O(N__5686),
            .I(N__5680));
    CascadeMux I__556 (
            .O(N__5683),
            .I(N__5677));
    CascadeMux I__555 (
            .O(N__5680),
            .I(N__5674));
    CascadeBuf I__554 (
            .O(N__5677),
            .I(N__5671));
    CascadeBuf I__553 (
            .O(N__5674),
            .I(N__5668));
    CascadeMux I__552 (
            .O(N__5671),
            .I(N__5665));
    CascadeMux I__551 (
            .O(N__5668),
            .I(N__5662));
    CascadeBuf I__550 (
            .O(N__5665),
            .I(N__5659));
    CascadeBuf I__549 (
            .O(N__5662),
            .I(N__5656));
    CascadeMux I__548 (
            .O(N__5659),
            .I(N__5653));
    CascadeMux I__547 (
            .O(N__5656),
            .I(N__5650));
    CascadeBuf I__546 (
            .O(N__5653),
            .I(N__5647));
    CascadeBuf I__545 (
            .O(N__5650),
            .I(N__5644));
    CascadeMux I__544 (
            .O(N__5647),
            .I(N__5641));
    CascadeMux I__543 (
            .O(N__5644),
            .I(N__5638));
    CascadeBuf I__542 (
            .O(N__5641),
            .I(N__5635));
    CascadeBuf I__541 (
            .O(N__5638),
            .I(N__5632));
    CascadeMux I__540 (
            .O(N__5635),
            .I(N__5629));
    CascadeMux I__539 (
            .O(N__5632),
            .I(N__5626));
    CascadeBuf I__538 (
            .O(N__5629),
            .I(N__5623));
    CascadeBuf I__537 (
            .O(N__5626),
            .I(N__5620));
    CascadeMux I__536 (
            .O(N__5623),
            .I(N__5617));
    CascadeMux I__535 (
            .O(N__5620),
            .I(N__5614));
    InMux I__534 (
            .O(N__5617),
            .I(N__5611));
    InMux I__533 (
            .O(N__5614),
            .I(N__5608));
    LocalMux I__532 (
            .O(N__5611),
            .I(N__5605));
    LocalMux I__531 (
            .O(N__5608),
            .I(N__5602));
    Span4Mux_s1_v I__530 (
            .O(N__5605),
            .I(N__5599));
    Span4Mux_v I__529 (
            .O(N__5602),
            .I(N__5596));
    Sp12to4 I__528 (
            .O(N__5599),
            .I(N__5593));
    IoSpan4Mux I__527 (
            .O(N__5596),
            .I(N__5590));
    Span12Mux_h I__526 (
            .O(N__5593),
            .I(N__5587));
    Odrv4 I__525 (
            .O(N__5590),
            .I(write_address_c_10));
    Odrv12 I__524 (
            .O(N__5587),
            .I(write_address_c_10));
    CascadeMux I__523 (
            .O(N__5582),
            .I(N__5579));
    CascadeBuf I__522 (
            .O(N__5579),
            .I(N__5576));
    CascadeMux I__521 (
            .O(N__5576),
            .I(N__5573));
    CascadeBuf I__520 (
            .O(N__5573),
            .I(N__5570));
    CascadeMux I__519 (
            .O(N__5570),
            .I(N__5567));
    CascadeBuf I__518 (
            .O(N__5567),
            .I(N__5564));
    CascadeMux I__517 (
            .O(N__5564),
            .I(N__5561));
    CascadeBuf I__516 (
            .O(N__5561),
            .I(N__5557));
    CascadeMux I__515 (
            .O(N__5560),
            .I(N__5554));
    CascadeMux I__514 (
            .O(N__5557),
            .I(N__5551));
    CascadeBuf I__513 (
            .O(N__5554),
            .I(N__5548));
    CascadeBuf I__512 (
            .O(N__5551),
            .I(N__5545));
    CascadeMux I__511 (
            .O(N__5548),
            .I(N__5542));
    CascadeMux I__510 (
            .O(N__5545),
            .I(N__5539));
    CascadeBuf I__509 (
            .O(N__5542),
            .I(N__5536));
    CascadeBuf I__508 (
            .O(N__5539),
            .I(N__5533));
    CascadeMux I__507 (
            .O(N__5536),
            .I(N__5530));
    CascadeMux I__506 (
            .O(N__5533),
            .I(N__5527));
    CascadeBuf I__505 (
            .O(N__5530),
            .I(N__5524));
    CascadeBuf I__504 (
            .O(N__5527),
            .I(N__5521));
    CascadeMux I__503 (
            .O(N__5524),
            .I(N__5518));
    CascadeMux I__502 (
            .O(N__5521),
            .I(N__5515));
    CascadeBuf I__501 (
            .O(N__5518),
            .I(N__5512));
    CascadeBuf I__500 (
            .O(N__5515),
            .I(N__5509));
    CascadeMux I__499 (
            .O(N__5512),
            .I(N__5506));
    CascadeMux I__498 (
            .O(N__5509),
            .I(N__5503));
    CascadeBuf I__497 (
            .O(N__5506),
            .I(N__5500));
    CascadeBuf I__496 (
            .O(N__5503),
            .I(N__5497));
    CascadeMux I__495 (
            .O(N__5500),
            .I(N__5494));
    CascadeMux I__494 (
            .O(N__5497),
            .I(N__5491));
    CascadeBuf I__493 (
            .O(N__5494),
            .I(N__5488));
    CascadeBuf I__492 (
            .O(N__5491),
            .I(N__5485));
    CascadeMux I__491 (
            .O(N__5488),
            .I(N__5482));
    CascadeMux I__490 (
            .O(N__5485),
            .I(N__5479));
    CascadeBuf I__489 (
            .O(N__5482),
            .I(N__5476));
    CascadeBuf I__488 (
            .O(N__5479),
            .I(N__5473));
    CascadeMux I__487 (
            .O(N__5476),
            .I(N__5470));
    CascadeMux I__486 (
            .O(N__5473),
            .I(N__5467));
    CascadeBuf I__485 (
            .O(N__5470),
            .I(N__5464));
    CascadeBuf I__484 (
            .O(N__5467),
            .I(N__5461));
    CascadeMux I__483 (
            .O(N__5464),
            .I(N__5458));
    CascadeMux I__482 (
            .O(N__5461),
            .I(N__5455));
    CascadeBuf I__481 (
            .O(N__5458),
            .I(N__5452));
    CascadeBuf I__480 (
            .O(N__5455),
            .I(N__5449));
    CascadeMux I__479 (
            .O(N__5452),
            .I(N__5446));
    CascadeMux I__478 (
            .O(N__5449),
            .I(N__5443));
    CascadeBuf I__477 (
            .O(N__5446),
            .I(N__5440));
    CascadeBuf I__476 (
            .O(N__5443),
            .I(N__5437));
    CascadeMux I__475 (
            .O(N__5440),
            .I(N__5434));
    CascadeMux I__474 (
            .O(N__5437),
            .I(N__5431));
    CascadeBuf I__473 (
            .O(N__5434),
            .I(N__5428));
    CascadeBuf I__472 (
            .O(N__5431),
            .I(N__5425));
    CascadeMux I__471 (
            .O(N__5428),
            .I(N__5422));
    CascadeMux I__470 (
            .O(N__5425),
            .I(N__5419));
    CascadeBuf I__469 (
            .O(N__5422),
            .I(N__5416));
    InMux I__468 (
            .O(N__5419),
            .I(N__5413));
    CascadeMux I__467 (
            .O(N__5416),
            .I(N__5410));
    LocalMux I__466 (
            .O(N__5413),
            .I(N__5407));
    CascadeBuf I__465 (
            .O(N__5410),
            .I(N__5404));
    Span4Mux_s3_v I__464 (
            .O(N__5407),
            .I(N__5401));
    CascadeMux I__463 (
            .O(N__5404),
            .I(N__5398));
    Span4Mux_h I__462 (
            .O(N__5401),
            .I(N__5395));
    InMux I__461 (
            .O(N__5398),
            .I(N__5392));
    Sp12to4 I__460 (
            .O(N__5395),
            .I(N__5389));
    LocalMux I__459 (
            .O(N__5392),
            .I(N__5386));
    Span12Mux_h I__458 (
            .O(N__5389),
            .I(N__5383));
    Odrv12 I__457 (
            .O(N__5386),
            .I(write_address_c_1));
    Odrv12 I__456 (
            .O(N__5383),
            .I(write_address_c_1));
    CascadeMux I__455 (
            .O(N__5378),
            .I(N__5375));
    CascadeBuf I__454 (
            .O(N__5375),
            .I(N__5372));
    CascadeMux I__453 (
            .O(N__5372),
            .I(N__5368));
    CascadeMux I__452 (
            .O(N__5371),
            .I(N__5365));
    CascadeBuf I__451 (
            .O(N__5368),
            .I(N__5362));
    CascadeBuf I__450 (
            .O(N__5365),
            .I(N__5359));
    CascadeMux I__449 (
            .O(N__5362),
            .I(N__5356));
    CascadeMux I__448 (
            .O(N__5359),
            .I(N__5353));
    CascadeBuf I__447 (
            .O(N__5356),
            .I(N__5350));
    CascadeBuf I__446 (
            .O(N__5353),
            .I(N__5347));
    CascadeMux I__445 (
            .O(N__5350),
            .I(N__5344));
    CascadeMux I__444 (
            .O(N__5347),
            .I(N__5341));
    CascadeBuf I__443 (
            .O(N__5344),
            .I(N__5338));
    CascadeBuf I__442 (
            .O(N__5341),
            .I(N__5335));
    CascadeMux I__441 (
            .O(N__5338),
            .I(N__5332));
    CascadeMux I__440 (
            .O(N__5335),
            .I(N__5329));
    CascadeBuf I__439 (
            .O(N__5332),
            .I(N__5326));
    CascadeBuf I__438 (
            .O(N__5329),
            .I(N__5323));
    CascadeMux I__437 (
            .O(N__5326),
            .I(N__5320));
    CascadeMux I__436 (
            .O(N__5323),
            .I(N__5317));
    CascadeBuf I__435 (
            .O(N__5320),
            .I(N__5314));
    CascadeBuf I__434 (
            .O(N__5317),
            .I(N__5311));
    CascadeMux I__433 (
            .O(N__5314),
            .I(N__5308));
    CascadeMux I__432 (
            .O(N__5311),
            .I(N__5305));
    CascadeBuf I__431 (
            .O(N__5308),
            .I(N__5302));
    CascadeBuf I__430 (
            .O(N__5305),
            .I(N__5299));
    CascadeMux I__429 (
            .O(N__5302),
            .I(N__5296));
    CascadeMux I__428 (
            .O(N__5299),
            .I(N__5293));
    CascadeBuf I__427 (
            .O(N__5296),
            .I(N__5290));
    CascadeBuf I__426 (
            .O(N__5293),
            .I(N__5287));
    CascadeMux I__425 (
            .O(N__5290),
            .I(N__5284));
    CascadeMux I__424 (
            .O(N__5287),
            .I(N__5281));
    CascadeBuf I__423 (
            .O(N__5284),
            .I(N__5278));
    CascadeBuf I__422 (
            .O(N__5281),
            .I(N__5275));
    CascadeMux I__421 (
            .O(N__5278),
            .I(N__5272));
    CascadeMux I__420 (
            .O(N__5275),
            .I(N__5269));
    CascadeBuf I__419 (
            .O(N__5272),
            .I(N__5266));
    CascadeBuf I__418 (
            .O(N__5269),
            .I(N__5263));
    CascadeMux I__417 (
            .O(N__5266),
            .I(N__5260));
    CascadeMux I__416 (
            .O(N__5263),
            .I(N__5257));
    CascadeBuf I__415 (
            .O(N__5260),
            .I(N__5254));
    CascadeBuf I__414 (
            .O(N__5257),
            .I(N__5251));
    CascadeMux I__413 (
            .O(N__5254),
            .I(N__5248));
    CascadeMux I__412 (
            .O(N__5251),
            .I(N__5245));
    CascadeBuf I__411 (
            .O(N__5248),
            .I(N__5242));
    CascadeBuf I__410 (
            .O(N__5245),
            .I(N__5239));
    CascadeMux I__409 (
            .O(N__5242),
            .I(N__5236));
    CascadeMux I__408 (
            .O(N__5239),
            .I(N__5233));
    CascadeBuf I__407 (
            .O(N__5236),
            .I(N__5230));
    CascadeBuf I__406 (
            .O(N__5233),
            .I(N__5227));
    CascadeMux I__405 (
            .O(N__5230),
            .I(N__5224));
    CascadeMux I__404 (
            .O(N__5227),
            .I(N__5221));
    CascadeBuf I__403 (
            .O(N__5224),
            .I(N__5218));
    CascadeBuf I__402 (
            .O(N__5221),
            .I(N__5215));
    CascadeMux I__401 (
            .O(N__5218),
            .I(N__5212));
    CascadeMux I__400 (
            .O(N__5215),
            .I(N__5209));
    CascadeBuf I__399 (
            .O(N__5212),
            .I(N__5206));
    InMux I__398 (
            .O(N__5209),
            .I(N__5203));
    CascadeMux I__397 (
            .O(N__5206),
            .I(N__5200));
    LocalMux I__396 (
            .O(N__5203),
            .I(N__5197));
    InMux I__395 (
            .O(N__5200),
            .I(N__5194));
    Span4Mux_v I__394 (
            .O(N__5197),
            .I(N__5191));
    LocalMux I__393 (
            .O(N__5194),
            .I(N__5188));
    Sp12to4 I__392 (
            .O(N__5191),
            .I(N__5185));
    Span4Mux_h I__391 (
            .O(N__5188),
            .I(N__5182));
    Span12Mux_h I__390 (
            .O(N__5185),
            .I(N__5179));
    Span4Mux_h I__389 (
            .O(N__5182),
            .I(N__5176));
    Odrv12 I__388 (
            .O(N__5179),
            .I(write_address_c_0));
    Odrv4 I__387 (
            .O(N__5176),
            .I(write_address_c_0));
    InMux I__386 (
            .O(N__5171),
            .I(N__5168));
    LocalMux I__385 (
            .O(N__5168),
            .I(N__5165));
    Span4Mux_s3_v I__384 (
            .O(N__5165),
            .I(N__5161));
    InMux I__383 (
            .O(N__5164),
            .I(N__5158));
    Span4Mux_v I__382 (
            .O(N__5161),
            .I(N__5151));
    LocalMux I__381 (
            .O(N__5158),
            .I(N__5151));
    InMux I__380 (
            .O(N__5157),
            .I(N__5148));
    InMux I__379 (
            .O(N__5156),
            .I(N__5145));
    Span4Mux_v I__378 (
            .O(N__5151),
            .I(N__5139));
    LocalMux I__377 (
            .O(N__5148),
            .I(N__5139));
    LocalMux I__376 (
            .O(N__5145),
            .I(N__5136));
    InMux I__375 (
            .O(N__5144),
            .I(N__5133));
    Span4Mux_v I__374 (
            .O(N__5139),
            .I(N__5130));
    Span4Mux_v I__373 (
            .O(N__5136),
            .I(N__5125));
    LocalMux I__372 (
            .O(N__5133),
            .I(N__5125));
    Span4Mux_v I__371 (
            .O(N__5130),
            .I(N__5119));
    Span4Mux_v I__370 (
            .O(N__5125),
            .I(N__5119));
    InMux I__369 (
            .O(N__5124),
            .I(N__5114));
    Span4Mux_h I__368 (
            .O(N__5119),
            .I(N__5109));
    InMux I__367 (
            .O(N__5118),
            .I(N__5106));
    InMux I__366 (
            .O(N__5117),
            .I(N__5103));
    LocalMux I__365 (
            .O(N__5114),
            .I(N__5100));
    InMux I__364 (
            .O(N__5113),
            .I(N__5097));
    InMux I__363 (
            .O(N__5112),
            .I(N__5094));
    Sp12to4 I__362 (
            .O(N__5109),
            .I(N__5091));
    LocalMux I__361 (
            .O(N__5106),
            .I(N__5086));
    LocalMux I__360 (
            .O(N__5103),
            .I(N__5086));
    Span12Mux_s7_v I__359 (
            .O(N__5100),
            .I(N__5079));
    LocalMux I__358 (
            .O(N__5097),
            .I(N__5079));
    LocalMux I__357 (
            .O(N__5094),
            .I(N__5079));
    Span12Mux_h I__356 (
            .O(N__5091),
            .I(N__5072));
    Span12Mux_v I__355 (
            .O(N__5086),
            .I(N__5072));
    Span12Mux_v I__354 (
            .O(N__5079),
            .I(N__5072));
    Odrv12 I__353 (
            .O(N__5072),
            .I(write_data_c_5));
    InMux I__352 (
            .O(N__5069),
            .I(N__5066));
    LocalMux I__351 (
            .O(N__5066),
            .I(N__5062));
    InMux I__350 (
            .O(N__5065),
            .I(N__5059));
    Span4Mux_v I__349 (
            .O(N__5062),
            .I(N__5054));
    LocalMux I__348 (
            .O(N__5059),
            .I(N__5054));
    Span4Mux_v I__347 (
            .O(N__5054),
            .I(N__5051));
    Span4Mux_v I__346 (
            .O(N__5051),
            .I(N__5047));
    InMux I__345 (
            .O(N__5050),
            .I(N__5044));
    Span4Mux_v I__344 (
            .O(N__5047),
            .I(N__5038));
    LocalMux I__343 (
            .O(N__5044),
            .I(N__5038));
    InMux I__342 (
            .O(N__5043),
            .I(N__5033));
    Span4Mux_v I__341 (
            .O(N__5038),
            .I(N__5030));
    InMux I__340 (
            .O(N__5037),
            .I(N__5026));
    InMux I__339 (
            .O(N__5036),
            .I(N__5022));
    LocalMux I__338 (
            .O(N__5033),
            .I(N__5019));
    Span4Mux_h I__337 (
            .O(N__5030),
            .I(N__5016));
    InMux I__336 (
            .O(N__5029),
            .I(N__5013));
    LocalMux I__335 (
            .O(N__5026),
            .I(N__5010));
    InMux I__334 (
            .O(N__5025),
            .I(N__5007));
    LocalMux I__333 (
            .O(N__5022),
            .I(N__5004));
    Span12Mux_h I__332 (
            .O(N__5019),
            .I(N__4999));
    Span4Mux_v I__331 (
            .O(N__5016),
            .I(N__4996));
    LocalMux I__330 (
            .O(N__5013),
            .I(N__4993));
    Span12Mux_s4_v I__329 (
            .O(N__5010),
            .I(N__4988));
    LocalMux I__328 (
            .O(N__5007),
            .I(N__4988));
    Span4Mux_v I__327 (
            .O(N__5004),
            .I(N__4985));
    InMux I__326 (
            .O(N__5003),
            .I(N__4982));
    InMux I__325 (
            .O(N__5002),
            .I(N__4979));
    Span12Mux_v I__324 (
            .O(N__4999),
            .I(N__4972));
    Sp12to4 I__323 (
            .O(N__4996),
            .I(N__4972));
    Span12Mux_h I__322 (
            .O(N__4993),
            .I(N__4972));
    Span12Mux_v I__321 (
            .O(N__4988),
            .I(N__4963));
    Sp12to4 I__320 (
            .O(N__4985),
            .I(N__4963));
    LocalMux I__319 (
            .O(N__4982),
            .I(N__4963));
    LocalMux I__318 (
            .O(N__4979),
            .I(N__4963));
    Span12Mux_h I__317 (
            .O(N__4972),
            .I(N__4958));
    Span12Mux_v I__316 (
            .O(N__4963),
            .I(N__4958));
    Odrv12 I__315 (
            .O(N__4958),
            .I(write_data_c_4));
    InMux I__314 (
            .O(N__4955),
            .I(N__4951));
    InMux I__313 (
            .O(N__4954),
            .I(N__4948));
    LocalMux I__312 (
            .O(N__4951),
            .I(N__4945));
    LocalMux I__311 (
            .O(N__4948),
            .I(N__4941));
    Span4Mux_s2_v I__310 (
            .O(N__4945),
            .I(N__4937));
    InMux I__309 (
            .O(N__4944),
            .I(N__4934));
    Span4Mux_s3_v I__308 (
            .O(N__4941),
            .I(N__4931));
    InMux I__307 (
            .O(N__4940),
            .I(N__4928));
    Span4Mux_v I__306 (
            .O(N__4937),
            .I(N__4921));
    LocalMux I__305 (
            .O(N__4934),
            .I(N__4921));
    Span4Mux_v I__304 (
            .O(N__4931),
            .I(N__4914));
    LocalMux I__303 (
            .O(N__4928),
            .I(N__4914));
    InMux I__302 (
            .O(N__4927),
            .I(N__4911));
    InMux I__301 (
            .O(N__4926),
            .I(N__4908));
    Span4Mux_h I__300 (
            .O(N__4921),
            .I(N__4904));
    InMux I__299 (
            .O(N__4920),
            .I(N__4901));
    InMux I__298 (
            .O(N__4919),
            .I(N__4898));
    Span4Mux_v I__297 (
            .O(N__4914),
            .I(N__4893));
    LocalMux I__296 (
            .O(N__4911),
            .I(N__4893));
    LocalMux I__295 (
            .O(N__4908),
            .I(N__4890));
    InMux I__294 (
            .O(N__4907),
            .I(N__4887));
    Span4Mux_v I__293 (
            .O(N__4904),
            .I(N__4882));
    LocalMux I__292 (
            .O(N__4901),
            .I(N__4882));
    LocalMux I__291 (
            .O(N__4898),
            .I(N__4879));
    Span4Mux_v I__290 (
            .O(N__4893),
            .I(N__4875));
    Span4Mux_v I__289 (
            .O(N__4890),
            .I(N__4870));
    LocalMux I__288 (
            .O(N__4887),
            .I(N__4870));
    Span4Mux_v I__287 (
            .O(N__4882),
            .I(N__4867));
    Span4Mux_v I__286 (
            .O(N__4879),
            .I(N__4864));
    InMux I__285 (
            .O(N__4878),
            .I(N__4861));
    Span4Mux_v I__284 (
            .O(N__4875),
            .I(N__4856));
    Span4Mux_v I__283 (
            .O(N__4870),
            .I(N__4856));
    Span4Mux_v I__282 (
            .O(N__4867),
            .I(N__4849));
    Span4Mux_v I__281 (
            .O(N__4864),
            .I(N__4849));
    LocalMux I__280 (
            .O(N__4861),
            .I(N__4849));
    Sp12to4 I__279 (
            .O(N__4856),
            .I(N__4846));
    Span4Mux_h I__278 (
            .O(N__4849),
            .I(N__4843));
    Span12Mux_h I__277 (
            .O(N__4846),
            .I(N__4840));
    IoSpan4Mux I__276 (
            .O(N__4843),
            .I(N__4837));
    Odrv12 I__275 (
            .O(N__4840),
            .I(write_data_c_3));
    Odrv4 I__274 (
            .O(N__4837),
            .I(write_data_c_3));
    InMux I__273 (
            .O(N__4832),
            .I(N__4829));
    LocalMux I__272 (
            .O(N__4829),
            .I(N__4825));
    InMux I__271 (
            .O(N__4828),
            .I(N__4822));
    Span4Mux_v I__270 (
            .O(N__4825),
            .I(N__4817));
    LocalMux I__269 (
            .O(N__4822),
            .I(N__4817));
    Span4Mux_v I__268 (
            .O(N__4817),
            .I(N__4812));
    InMux I__267 (
            .O(N__4816),
            .I(N__4809));
    InMux I__266 (
            .O(N__4815),
            .I(N__4805));
    Span4Mux_v I__265 (
            .O(N__4812),
            .I(N__4799));
    LocalMux I__264 (
            .O(N__4809),
            .I(N__4799));
    InMux I__263 (
            .O(N__4808),
            .I(N__4796));
    LocalMux I__262 (
            .O(N__4805),
            .I(N__4793));
    InMux I__261 (
            .O(N__4804),
            .I(N__4790));
    Span4Mux_v I__260 (
            .O(N__4799),
            .I(N__4785));
    LocalMux I__259 (
            .O(N__4796),
            .I(N__4785));
    Span4Mux_v I__258 (
            .O(N__4793),
            .I(N__4779));
    LocalMux I__257 (
            .O(N__4790),
            .I(N__4779));
    Span4Mux_v I__256 (
            .O(N__4785),
            .I(N__4775));
    InMux I__255 (
            .O(N__4784),
            .I(N__4772));
    Span4Mux_v I__254 (
            .O(N__4779),
            .I(N__4769));
    InMux I__253 (
            .O(N__4778),
            .I(N__4766));
    Span4Mux_v I__252 (
            .O(N__4775),
            .I(N__4760));
    LocalMux I__251 (
            .O(N__4772),
            .I(N__4760));
    Span4Mux_v I__250 (
            .O(N__4769),
            .I(N__4755));
    LocalMux I__249 (
            .O(N__4766),
            .I(N__4755));
    InMux I__248 (
            .O(N__4765),
            .I(N__4752));
    Span4Mux_v I__247 (
            .O(N__4760),
            .I(N__4749));
    Span4Mux_v I__246 (
            .O(N__4755),
            .I(N__4744));
    LocalMux I__245 (
            .O(N__4752),
            .I(N__4744));
    Span4Mux_h I__244 (
            .O(N__4749),
            .I(N__4740));
    Span4Mux_v I__243 (
            .O(N__4744),
            .I(N__4737));
    InMux I__242 (
            .O(N__4743),
            .I(N__4734));
    Sp12to4 I__241 (
            .O(N__4740),
            .I(N__4731));
    Span4Mux_v I__240 (
            .O(N__4737),
            .I(N__4726));
    LocalMux I__239 (
            .O(N__4734),
            .I(N__4726));
    Span12Mux_h I__238 (
            .O(N__4731),
            .I(N__4723));
    Span4Mux_v I__237 (
            .O(N__4726),
            .I(N__4720));
    Odrv12 I__236 (
            .O(N__4723),
            .I(write_data_c_2));
    Odrv4 I__235 (
            .O(N__4720),
            .I(write_data_c_2));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_6_cry_7 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_6_THRU_CO ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\this_vga_signals.address_1_0_8 ),
            .carryinitout(bfn_13_18_0_));
    ICE_GB \this_reset_cond.M_stage_q_RNI6VB7_3  (
            .USERSIGNALTOGLOBALBUFFER(N__12070),
            .GLOBALBUFFEROUTPUT(N_112_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_0_LC_1_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_0_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_0_LC_1_16_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \this_vga_signals.M_hstate_q_RNI1P4R_0_0_LC_1_16_2  (
            .in0(N__11797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12139),
            .lcout(this_vga_signals_N_170_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_1_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_1_17_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_hstate_q_RNI1P4R_0_LC_1_17_4  (
            .in0(N__11784),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12126),
            .lcout(this_vga_signals_N_171_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNIUAUT_0_LC_1_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNIUAUT_0_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNIUAUT_0_LC_1_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_hstate_q_RNIUAUT_0_LC_1_18_0  (
            .in0(N__12140),
            .in1(N__10471),
            .in2(N__10520),
            .in3(N__11798),
            .lcout(rgb5_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_0_LC_1_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_0_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_0_LC_1_18_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_vstate_q_RNITHP2_0_0_LC_1_18_7  (
            .in0(N__10472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10519),
            .lcout(vsync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_LC_2_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNITHP2_0_LC_2_18_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_vstate_q_RNITHP2_0_LC_2_18_4  (
            .in0(N__10465),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10515),
            .lcout(this_vga_signals_N_94_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNILGF11_LC_7_7_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNILGF11_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNILGF11_LC_7_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_0_0_RNILGF11_LC_7_7_2  (
            .in0(N__14436),
            .in1(N__7808),
            .in2(_gnd_net_),
            .in3(N__7796),
            .lcout(\this_vram.mem_mem_0_0_RNILGFZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNINGF11_LC_7_9_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNINGF11_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNINGF11_LC_7_9_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_0_1_RNINGF11_LC_7_9_2  (
            .in0(N__7790),
            .in1(N__14477),
            .in2(_gnd_net_),
            .in3(N__7778),
            .lcout(\this_vram.mem_mem_0_1_RNINGFZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_1_RNINGF11_0_LC_7_9_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_1_RNINGF11_0_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_1_RNINGF11_0_LC_7_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_0_1_RNINGF11_0_LC_7_9_7  (
            .in0(N__14476),
            .in1(N__8036),
            .in2(_gnd_net_),
            .in3(N__8024),
            .lcout(\this_vram.mem_mem_0_1_RNINGF11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_2_RNIPGF11_LC_7_11_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_2_RNIPGF11_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_2_RNIPGF11_LC_7_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_0_2_RNIPGF11_LC_7_11_4  (
            .in0(N__8018),
            .in1(N__14463),
            .in2(_gnd_net_),
            .in3(N__8006),
            .lcout(\this_vram.mem_mem_0_2_RNIPGFZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_2_RNIPGF11_0_LC_7_11_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_2_RNIPGF11_0_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_2_RNIPGF11_0_LC_7_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_0_2_RNIPGF11_0_LC_7_11_5  (
            .in0(N__14462),
            .in1(N__8000),
            .in2(_gnd_net_),
            .in3(N__7994),
            .lcout(\this_vram.mem_mem_0_2_RNIPGF11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIPOJ11_LC_7_13_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIPOJ11_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIPOJ11_LC_7_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_2_0_RNIPOJ11_LC_7_13_0  (
            .in0(N__7982),
            .in1(N__14456),
            .in2(_gnd_net_),
            .in3(N__7970),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_0_RNIPOJZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNINVA72_0_12_LC_7_13_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNINVA72_0_12_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNINVA72_0_12_LC_7_13_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vram.mem_radreg_RNINVA72_0_12_LC_7_13_1  (
            .in0(N__7964),
            .in1(_gnd_net_),
            .in2(N__7955),
            .in3(N__14175),
            .lcout(\this_vram.mem_N_2362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OEJ4_0_13_LC_7_15_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OEJ4_0_13_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OEJ4_0_13_LC_7_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNI9OEJ4_0_13_LC_7_15_2  (
            .in0(N__8381),
            .in1(N__7952),
            .in2(_gnd_net_),
            .in3(N__10273),
            .lcout(),
            .ltout(\this_vram.mem_N_2364_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIN7E66_0_14_LC_7_15_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIN7E66_0_14_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIN7E66_0_14_LC_7_15_3 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \this_vram.mem_radreg_RNIN7E66_0_14_LC_7_15_3  (
            .in0(N__8732),
            .in1(N__13946),
            .in2(N__7943),
            .in3(N__10202),
            .lcout(M_this_vram_read_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNIROJ11_0_LC_7_15_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNIROJ11_0_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNIROJ11_0_LC_7_15_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_2_1_RNIROJ11_0_LC_7_15_4  (
            .in0(N__7928),
            .in1(N__14361),
            .in2(_gnd_net_),
            .in3(N__7916),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_1_RNIROJ11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIRVA72_12_LC_7_15_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIRVA72_12_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIRVA72_12_LC_7_15_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vram.mem_radreg_RNIRVA72_12_LC_7_15_5  (
            .in0(N__8165),
            .in1(_gnd_net_),
            .in2(N__8156),
            .in3(N__14097),
            .lcout(\this_vram.mem_N_2335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_1_RNI14P11_0_LC_7_16_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_1_RNI14P11_0_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_1_RNI14P11_0_LC_7_16_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_4_1_RNI14P11_0_LC_7_16_1  (
            .in0(N__14171),
            .in1(N__8153),
            .in2(_gnd_net_),
            .in3(N__8138),
            .lcout(),
            .ltout(\this_vram.mem_mem_4_1_RNI14P11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIC1S72_11_LC_7_16_2 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIC1S72_11_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIC1S72_11_LC_7_16_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vram.mem_radreg_RNIC1S72_11_LC_7_16_2  (
            .in0(N__12749),
            .in1(_gnd_net_),
            .in2(N__8117),
            .in3(N__14453),
            .lcout(),
            .ltout(\this_vram.mem_N_2336_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIHOEJ4_13_LC_7_16_3 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIHOEJ4_13_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIHOEJ4_13_LC_7_16_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNIHOEJ4_13_LC_7_16_3  (
            .in0(N__10293),
            .in1(_gnd_net_),
            .in2(N__8114),
            .in3(N__8111),
            .lcout(\this_vram.mem_N_2337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_1_RNIROJ11_LC_7_16_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_1_RNIROJ11_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_1_RNIROJ11_LC_7_16_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_2_1_RNIROJ11_LC_7_16_6  (
            .in0(N__8105),
            .in1(N__14452),
            .in2(_gnd_net_),
            .in3(N__8093),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_1_RNIROJZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIRVA72_0_12_LC_7_16_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIRVA72_0_12_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIRVA72_0_12_LC_7_16_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNIRVA72_0_12_LC_7_16_7  (
            .in0(N__14172),
            .in1(_gnd_net_),
            .in2(N__8087),
            .in3(N__8084),
            .lcout(\this_vram.mem_N_2344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_2_RNITOJ11_0_LC_7_17_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_2_RNITOJ11_0_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_2_RNITOJ11_0_LC_7_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_2_2_RNITOJ11_0_LC_7_17_4  (
            .in0(N__8072),
            .in1(N__14454),
            .in2(_gnd_net_),
            .in3(N__8060),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_2_RNITOJ11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIVVA72_12_LC_7_17_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIVVA72_12_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIVVA72_12_LC_7_17_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vram.mem_radreg_RNIVVA72_12_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__8054),
            .in2(N__8042),
            .in3(N__14173),
            .lcout(),
            .ltout(\this_vram.mem_N_2371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIPOEJ4_13_LC_7_17_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIPOEJ4_13_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIPOEJ4_13_LC_7_17_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vram.mem_radreg_RNIPOEJ4_13_LC_7_17_6  (
            .in0(N__10294),
            .in1(_gnd_net_),
            .in2(N__8039),
            .in3(N__13466),
            .lcout(\this_vram.mem_N_2373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_2_RNITOJ11_LC_7_18_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_2_RNITOJ11_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_2_RNITOJ11_LC_7_18_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_2_2_RNITOJ11_LC_7_18_5  (
            .in0(N__8318),
            .in1(N__14455),
            .in2(_gnd_net_),
            .in3(N__8312),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_2_RNITOJZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIVVA72_0_12_LC_7_18_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIVVA72_0_12_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIVVA72_0_12_LC_7_18_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \this_vram.mem_radreg_RNIVVA72_0_12_LC_7_18_6  (
            .in0(N__14174),
            .in1(N__8300),
            .in2(N__8288),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_vram.mem_N_2326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIPOEJ4_0_13_LC_7_18_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIPOEJ4_0_13_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIPOEJ4_0_13_LC_7_18_7 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \this_vram.mem_radreg_RNIPOEJ4_0_13_LC_7_18_7  (
            .in0(N__10295),
            .in1(N__8765),
            .in2(N__8285),
            .in3(_gnd_net_),
            .lcout(\this_vram.mem_N_2328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIB8E66_14_LC_7_20_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIB8E66_14_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIB8E66_14_LC_7_20_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \this_vram.mem_radreg_RNIB8E66_14_LC_7_20_1  (
            .in0(N__10230),
            .in1(N__12827),
            .in2(N__8282),
            .in3(N__8733),
            .lcout(M_this_vram_read_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIB8E66_0_14_LC_7_21_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIB8E66_0_14_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIB8E66_0_14_LC_7_21_0 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \this_vram.mem_radreg_RNIB8E66_0_14_LC_7_21_0  (
            .in0(N__8252),
            .in1(N__14267),
            .in2(N__8741),
            .in3(N__10232),
            .lcout(M_this_vram_read_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI18E66_14_LC_7_21_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI18E66_14_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI18E66_14_LC_7_21_6 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \this_vram.mem_radreg_RNI18E66_14_LC_7_21_6  (
            .in0(N__8225),
            .in1(N__14492),
            .in2(N__8740),
            .in3(N__10231),
            .lcout(M_this_vram_read_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_RNILGF11_0_LC_9_7_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_RNILGF11_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_RNILGF11_0_LC_9_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_0_0_RNILGF11_0_LC_9_7_7  (
            .in0(N__14435),
            .in1(N__8201),
            .in2(_gnd_net_),
            .in3(N__8189),
            .lcout(\this_vram.mem_mem_0_0_RNILGF11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_RNIPOJ11_0_LC_9_13_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_RNIPOJ11_0_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_RNIPOJ11_0_LC_9_13_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_2_0_RNIPOJ11_0_LC_9_13_3  (
            .in0(N__8183),
            .in1(N__14425),
            .in2(_gnd_net_),
            .in3(N__8171),
            .lcout(),
            .ltout(\this_vram.mem_mem_2_0_RNIPOJ11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNINVA72_12_LC_9_13_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNINVA72_12_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNINVA72_12_LC_9_13_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \this_vram.mem_radreg_RNINVA72_12_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__8507),
            .in2(N__8498),
            .in3(N__14157),
            .lcout(\this_vram.mem_N_2353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_RNIV3P11_LC_9_15_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_RNIV3P11_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_RNIV3P11_LC_9_15_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_4_0_RNIV3P11_LC_9_15_1  (
            .in0(N__8495),
            .in1(N__14095),
            .in2(_gnd_net_),
            .in3(N__8474),
            .lcout(\this_vram.mem_mem_4_0_RNIV3PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_0_0_wclke_0_a2_LC_9_15_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_0_0_wclke_0_a2_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_0_0_wclke_0_a2_LC_9_15_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vram.mem_mem_0_0_wclke_0_a2_LC_9_15_5  (
            .in0(N__14804),
            .in1(N__14900),
            .in2(N__14681),
            .in3(N__13864),
            .lcout(\this_vram.mem_WE_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_0_RNI18R11_LC_9_15_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_0_RNI18R11_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_0_RNI18R11_LC_9_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_5_0_RNI18R11_LC_9_15_6  (
            .in0(N__14096),
            .in1(N__8429),
            .in2(_gnd_net_),
            .in3(N__8408),
            .lcout(),
            .ltout(\this_vram.mem_mem_5_0_RNI18RZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI81S72_0_11_LC_9_15_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI81S72_0_11_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI81S72_0_11_LC_9_15_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vram.mem_radreg_RNI81S72_0_11_LC_9_15_7  (
            .in0(N__14357),
            .in1(_gnd_net_),
            .in2(N__8390),
            .in3(N__8387),
            .lcout(\this_vram.mem_N_2363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIHOEJ4_0_13_LC_9_16_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIHOEJ4_0_13_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIHOEJ4_0_13_LC_9_16_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_radreg_RNIHOEJ4_0_13_LC_9_16_0  (
            .in0(N__10281),
            .in1(N__8813),
            .in2(_gnd_net_),
            .in3(N__8369),
            .lcout(\this_vram.mem_N_2346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIU5NC_13_LC_9_17_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIU5NC_13_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIU5NC_13_LC_9_17_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \this_vram.mem_radreg_RNIU5NC_13_LC_9_17_5  (
            .in0(N__10215),
            .in1(N__10282),
            .in2(_gnd_net_),
            .in3(N__14161),
            .lcout(\this_vram.mem_G_25_0 ),
            .ltout(\this_vram.mem_G_25_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI18E66_0_14_LC_9_17_6 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI18E66_0_14_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI18E66_0_14_LC_9_17_6 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \this_vram.mem_radreg_RNI18E66_0_14_LC_9_17_6  (
            .in0(N__13880),
            .in1(N__8360),
            .in2(N__8354),
            .in3(N__10214),
            .lcout(M_this_vram_read_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_2_0_wclke_0_a2_LC_9_17_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_2_0_wclke_0_a2_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_2_0_wclke_0_a2_LC_9_17_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vram.mem_mem_2_0_wclke_0_a2_LC_9_17_7  (
            .in0(N__14803),
            .in1(N__14895),
            .in2(N__13860),
            .in3(N__14676),
            .lcout(\this_vram.mem_WE_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIG1S72_0_11_LC_9_18_0 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIG1S72_0_11_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIG1S72_0_11_LC_9_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_radreg_RNIG1S72_0_11_LC_9_18_0  (
            .in0(N__14201),
            .in1(N__8654),
            .in2(_gnd_net_),
            .in3(N__14431),
            .lcout(\this_vram.mem_N_2327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI9OEJ4_13_LC_9_18_4 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI9OEJ4_13_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI9OEJ4_13_LC_9_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_radreg_RNI9OEJ4_13_LC_9_18_4  (
            .in0(N__10283),
            .in1(N__8543),
            .in2(_gnd_net_),
            .in3(N__8756),
            .lcout(),
            .ltout(\this_vram.mem_N_2355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIN7E66_14_LC_9_18_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIN7E66_14_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIN7E66_14_LC_9_18_5 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \this_vram.mem_radreg_RNIN7E66_14_LC_9_18_5  (
            .in0(N__10216),
            .in1(N__13913),
            .in2(N__8744),
            .in3(N__8712),
            .lcout(M_this_vram_read_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_2_RNI34P11_LC_9_19_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_2_RNI34P11_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_2_RNI34P11_LC_9_19_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_4_2_RNI34P11_LC_9_19_0  (
            .in0(N__8690),
            .in1(N__14170),
            .in2(_gnd_net_),
            .in3(N__8675),
            .lcout(\this_vram.mem_mem_4_2_RNI34PZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_3_0_wclke_0_a2_LC_9_19_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_3_0_wclke_0_a2_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_3_0_wclke_0_a2_LC_9_19_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vram.mem_mem_3_0_wclke_0_a2_LC_9_19_1  (
            .in0(N__14793),
            .in1(N__14885),
            .in2(N__13859),
            .in3(N__14675),
            .lcout(\this_vram.mem_WE_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_RNIV3P11_0_LC_9_20_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_RNIV3P11_0_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_RNIV3P11_0_LC_9_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_4_0_RNIV3P11_0_LC_9_20_3  (
            .in0(N__8621),
            .in1(N__8600),
            .in2(_gnd_net_),
            .in3(N__14176),
            .lcout(\this_vram.mem_mem_4_0_RNIV3P11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_0_RNI18R11_0_LC_9_20_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_0_RNI18R11_0_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_0_RNI18R11_0_LC_9_20_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_5_0_RNI18R11_0_LC_9_20_6  (
            .in0(N__8588),
            .in1(N__14177),
            .in2(_gnd_net_),
            .in3(N__8573),
            .lcout(),
            .ltout(\this_vram.mem_mem_5_0_RNI18R11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNI81S72_11_LC_9_20_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNI81S72_11_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNI81S72_11_LC_9_20_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vram.mem_radreg_RNI81S72_11_LC_9_20_7  (
            .in0(N__8552),
            .in1(_gnd_net_),
            .in2(N__8546),
            .in3(N__14464),
            .lcout(\this_vram.mem_N_2354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_1_0_wclke_0_a2_LC_10_15_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_1_0_wclke_0_a2_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_1_0_wclke_0_a2_LC_10_15_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_vram.mem_mem_1_0_wclke_0_a2_LC_10_15_5  (
            .in0(N__14680),
            .in1(N__14899),
            .in2(N__13865),
            .in3(N__14784),
            .lcout(\this_vram.mem_WE_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_1_RNI14P11_LC_10_16_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_1_RNI14P11_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_1_RNI14P11_LC_10_16_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_4_1_RNI14P11_LC_10_16_0  (
            .in0(N__8852),
            .in1(N__14141),
            .in2(_gnd_net_),
            .in3(N__8837),
            .lcout(),
            .ltout(\this_vram.mem_mem_4_1_RNI14PZ0Z11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIC1S72_0_11_LC_10_16_1 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIC1S72_0_11_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIC1S72_0_11_LC_10_16_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vram.mem_radreg_RNIC1S72_0_11_LC_10_16_1  (
            .in0(N__12788),
            .in1(_gnd_net_),
            .in2(N__8816),
            .in3(N__14407),
            .lcout(\this_vram.mem_N_2345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_wclke_0_a2_LC_10_21_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_wclke_0_a2_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_wclke_0_a2_LC_10_21_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_vram.mem_mem_4_0_wclke_0_a2_LC_10_21_1  (
            .in0(N__14774),
            .in1(N__14864),
            .in2(N__13858),
            .in3(N__14659),
            .lcout(\this_vram.mem_WE_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_o2_LC_12_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_o2_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_o2_LC_12_17_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m24_0_o2_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__10792),
            .in2(_gnd_net_),
            .in3(N__10729),
            .lcout(\this_vga_signals.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_1_LC_12_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_1_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_1_LC_12_17_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_1_LC_12_17_2  (
            .in0(N__10730),
            .in1(N__10834),
            .in2(_gnd_net_),
            .in3(N__10793),
            .lcout(\this_vga_signals.m27_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_LC_12_18_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_LC_12_18_0  (
            .in0(N__10539),
            .in1(N__10409),
            .in2(N__10462),
            .in3(N__10309),
            .lcout(),
            .ltout(\this_vga_signals.m24_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_LC_12_18_1 .LUT_INIT=16'b1111010111111001;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m24_0_LC_12_18_1  (
            .in0(N__10500),
            .in1(N__8771),
            .in2(N__8777),
            .in3(N__9715),
            .lcout(),
            .ltout(\this_vga_signals.N_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_0_LC_12_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_0_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_0_LC_12_18_2 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \this_vga_signals.M_vstate_q_0_LC_12_18_2  (
            .in0(N__12076),
            .in1(N__10501),
            .in2(N__8774),
            .in3(N__10680),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13692),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_0_LC_12_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_0_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_0_LC_12_18_3 .LUT_INIT=16'b0000001001010110;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m24_0_1_0_LC_12_18_3  (
            .in0(N__10498),
            .in1(N__9730),
            .in2(N__10464),
            .in3(N__10842),
            .lcout(\this_vga_signals.m24_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_0_LC_12_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_0_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_0_LC_12_18_4 .LUT_INIT=16'b1000101100000011;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m27_0_0_LC_12_18_4  (
            .in0(N__10540),
            .in1(N__10499),
            .in2(N__10463),
            .in3(N__10310),
            .lcout(),
            .ltout(\this_vga_signals.m27_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_LC_12_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_LC_12_18_5 .LUT_INIT=16'b1111010111110100;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m27_0_LC_12_18_5  (
            .in0(N__10453),
            .in1(N__9731),
            .in2(N__9722),
            .in3(N__9716),
            .lcout(),
            .ltout(\this_vga_signals.i9_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_1_LC_12_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_1_LC_12_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vstate_q_1_LC_12_18_6 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \this_vga_signals.M_vstate_q_1_LC_12_18_6  (
            .in0(N__12077),
            .in1(N__10454),
            .in2(N__9719),
            .in3(N__10681),
            .lcout(\this_vga_signals.M_vstate_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13692),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_LC_12_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_LC_12_18_7 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_LC_12_18_7  (
            .in0(N__11986),
            .in1(N__10933),
            .in2(_gnd_net_),
            .in3(N__10322),
            .lcout(\this_vga_signals.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI8NSN1_2_LC_13_15_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_RNI8NSN1_2_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI8NSN1_2_LC_13_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI8NSN1_2_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__10788),
            .in2(N__9758),
            .in3(_gnd_net_),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\this_vga_signals.address_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_cry_0_c_RNI17SC1_LC_13_15_1 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_cry_0_c_RNI17SC1_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_cry_0_c_RNI17SC1_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.address_1_cry_0_c_RNI17SC1_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__10728),
            .in2(N__9743),
            .in3(N__9293),
            .lcout(M_this_vga_signals_address_8),
            .ltout(),
            .carryin(\this_vga_signals.address_1_cry_0 ),
            .carryout(\this_vga_signals.address_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_cry_1_c_RNI5DUC1_LC_13_15_2 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_cry_1_c_RNI5DUC1_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_cry_1_c_RNI5DUC1_LC_13_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.address_1_cry_1_c_RNI5DUC1_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__10682),
            .in2(N__10388),
            .in3(N__9074),
            .lcout(M_this_vga_signals_address_9),
            .ltout(),
            .carryin(\this_vga_signals.address_1_cry_1 ),
            .carryout(\this_vga_signals.address_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_cry_2_c_RNI9J0D1_LC_13_15_3 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_cry_2_c_RNI9J0D1_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_cry_2_c_RNI9J0D1_LC_13_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.address_1_cry_2_c_RNI9J0D1_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__10637),
            .in2(N__10373),
            .in3(N__8858),
            .lcout(M_this_vga_signals_address_10),
            .ltout(),
            .carryin(\this_vga_signals.address_1_cry_2 ),
            .carryout(\this_vga_signals.address_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_11_LC_13_15_4 .C_ON=1'b1;
    defparam \this_vram.mem_radreg_11_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_11_LC_13_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vram.mem_radreg_11_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__10358),
            .in2(N__10601),
            .in3(N__8855),
            .lcout(\this_vram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_cry_3 ),
            .carryout(\this_vga_signals.address_1_cry_4 ),
            .clk(N__13676),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_12_LC_13_15_5 .C_ON=1'b1;
    defparam \this_vram.mem_radreg_12_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_12_LC_13_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vram.mem_radreg_12_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__10346),
            .in2(N__10973),
            .in3(N__10298),
            .lcout(\this_vram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_cry_4 ),
            .carryout(\this_vga_signals.address_1_cry_5 ),
            .clk(N__13676),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_13_LC_13_15_6 .C_ON=1'b1;
    defparam \this_vram.mem_radreg_13_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_13_LC_13_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vram.mem_radreg_13_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__10331),
            .in2(N__10934),
            .in3(N__10238),
            .lcout(\this_vram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_cry_5 ),
            .carryout(\this_vga_signals.address_1_cry_6 ),
            .clk(N__13676),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_14_LC_13_15_7 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_14_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \this_vram.mem_radreg_14_LC_13_15_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vram.mem_radreg_14_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__11987),
            .in2(_gnd_net_),
            .in3(N__10235),
            .lcout(\this_vram.mem_radregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13676),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_13_16_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_13_16_0  (
            .in0(N__12015),
            .in1(N__10797),
            .in2(N__11936),
            .in3(N__10751),
            .lcout(\this_vga_signals.address_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13681),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_16_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_13_16_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_13_16_5  (
            .in0(N__10737),
            .in1(N__12016),
            .in2(N__10697),
            .in3(N__11933),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13681),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNINV7N_9_LC_13_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_RNINV7N_9_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNINV7N_9_LC_13_17_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNINV7N_9_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__10787),
            .in2(N__11747),
            .in3(_gnd_net_),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\this_vga_signals.address_1_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_cry_0_c_RNIM2N91_LC_13_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_0_cry_0_c_RNIM2N91_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_cry_0_c_RNIM2N91_LC_13_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.address_1_0_cry_0_c_RNIM2N91_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__10727),
            .in2(N__11712),
            .in3(N__9761),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(\this_vga_signals.address_1_0_cry_0 ),
            .carryout(\this_vga_signals.address_1_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_cry_1_c_RNIP6O91_LC_13_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_0_cry_1_c_RNIP6O91_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_cry_1_c_RNIP6O91_LC_13_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.address_1_0_cry_1_c_RNIP6O91_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__10666),
            .in2(N__12490),
            .in3(N__9746),
            .lcout(\this_vga_signals.address_1 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_0_cry_1 ),
            .carryout(\this_vga_signals.address_1_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_cry_2_c_RNIADGT_LC_13_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_0_cry_2_c_RNIADGT_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_cry_2_c_RNIADGT_LC_13_17_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.address_1_0_cry_2_c_RNIADGT_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10636),
            .in3(N__10391),
            .lcout(\this_vga_signals.address_1_0_3 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_0_cry_2 ),
            .carryout(\this_vga_signals.address_1_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_cry_3_c_RNICGHT_LC_13_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_0_cry_3_c_RNICGHT_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_cry_3_c_RNICGHT_LC_13_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.address_1_0_cry_3_c_RNICGHT_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__10588),
            .in2(_gnd_net_),
            .in3(N__10376),
            .lcout(\this_vga_signals.address_1_0_4 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_0_cry_3 ),
            .carryout(\this_vga_signals.address_1_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_cry_4_c_RNIEJIT_LC_13_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_0_cry_4_c_RNIEJIT_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_cry_4_c_RNIEJIT_LC_13_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.address_1_0_cry_4_c_RNIEJIT_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__10960),
            .in2(_gnd_net_),
            .in3(N__10361),
            .lcout(\this_vga_signals.address_1_0_5 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_0_cry_4 ),
            .carryout(\this_vga_signals.address_1_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_cry_5_c_RNIGMJT_LC_13_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_0_cry_5_c_RNIGMJT_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_cry_5_c_RNIGMJT_LC_13_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.address_1_0_cry_5_c_RNIGMJT_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__10923),
            .in2(_gnd_net_),
            .in3(N__10349),
            .lcout(\this_vga_signals.address_1_0_6 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_0_cry_5 ),
            .carryout(\this_vga_signals.address_1_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_cry_6_c_RNIIPKT_LC_13_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.address_1_0_cry_6_c_RNIIPKT_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_cry_6_c_RNIIPKT_LC_13_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.address_1_0_cry_6_c_RNIIPKT_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__11984),
            .in2(_gnd_net_),
            .in3(N__10337),
            .lcout(\this_vga_signals.address_1_0_7 ),
            .ltout(),
            .carryin(\this_vga_signals.address_1_0_cry_6 ),
            .carryout(\this_vga_signals.address_1_0_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.address_1_0_8_THRU_LUT4_0_LC_13_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.address_1_0_8_THRU_LUT4_0_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.address_1_0_8_THRU_LUT4_0_LC_13_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.address_1_0_8_THRU_LUT4_0_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10334),
            .lcout(\this_vga_signals.address_1_0_8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_3_LC_13_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_3_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_3_LC_13_18_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m27_0_o2_0_3_LC_13_18_1  (
            .in0(N__10961),
            .in1(N__10589),
            .in2(N__10869),
            .in3(N__10630),
            .lcout(\this_vga_signals.m27_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_5_LC_13_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_5_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_5_LC_13_18_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_5_LC_13_18_2  (
            .in0(N__10631),
            .in1(N__10862),
            .in2(N__10843),
            .in3(N__10316),
            .lcout(\this_vga_signals.m27_0_a2_1_5 ),
            .ltout(\this_vga_signals.m27_0_a2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNICG7G4_1_LC_13_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNICG7G4_1_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNICG7G4_1_LC_13_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_vstate_q_RNICG7G4_1_LC_13_18_3  (
            .in0(N__10443),
            .in1(N__10526),
            .in2(N__10301),
            .in3(N__10541),
            .lcout(\this_vga_signals.N_68 ),
            .ltout(\this_vga_signals.N_68_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_13_18_4 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_13_18_4  (
            .in0(N__10838),
            .in1(N__11929),
            .in2(N__10544),
            .in3(N__10811),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13688),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_4_LC_13_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_4_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_4_LC_13_18_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m27_0_a2_1_4_LC_13_18_5  (
            .in0(N__10962),
            .in1(N__10918),
            .in2(N__11985),
            .in3(N__10590),
            .lcout(\this_vga_signals.m27_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_RNIVAHF_0_LC_13_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_RNIVAHF_0_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_RNIVAHF_0_LC_13_18_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_vstate_q_RNIVAHF_0_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__10496),
            .in2(_gnd_net_),
            .in3(N__10670),
            .lcout(\this_vga_signals.M_vcounter_q_0_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_0_LC_13_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_0_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vstate_q_ns_1_0__m24_0_0_LC_13_18_7 .LUT_INIT=16'b0001010101010100;
    LogicCell40 \this_vga_signals.M_vstate_q_ns_1_0__m24_0_0_LC_13_18_7  (
            .in0(N__10497),
            .in1(N__10799),
            .in2(N__10461),
            .in3(N__10739),
            .lcout(\this_vga_signals.m24_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_14_15_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__11865),
            .in2(N__11834),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_14_15_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_14_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__11846),
            .in2(_gnd_net_),
            .in3(N__10403),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__13673),
            .ce(),
            .sr(N__11908));
    defparam \this_vga_signals.M_hcounter_q_3_LC_14_15_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_14_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__11810),
            .in2(_gnd_net_),
            .in3(N__10400),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__13673),
            .ce(),
            .sr(N__11908));
    defparam \this_vga_signals.M_hcounter_q_4_LC_14_15_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_14_15_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_14_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__12520),
            .in2(_gnd_net_),
            .in3(N__10397),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__13673),
            .ce(),
            .sr(N__11908));
    defparam \this_vga_signals.M_hcounter_q_5_LC_14_15_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_14_15_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_14_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__12271),
            .in2(_gnd_net_),
            .in3(N__10394),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__13673),
            .ce(),
            .sr(N__11908));
    defparam \this_vga_signals.M_hcounter_q_6_LC_14_15_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_14_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__11481),
            .in2(_gnd_net_),
            .in3(N__10562),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__13673),
            .ce(),
            .sr(N__11908));
    defparam \this_vga_signals.M_hcounter_q_7_LC_14_15_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_14_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_14_15_6  (
            .in0(N__12227),
            .in1(N__11251),
            .in2(_gnd_net_),
            .in3(N__10559),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__13673),
            .ce(),
            .sr(N__11908));
    defparam \this_vga_signals.M_hcounter_q_8_LC_14_15_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_14_15_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_14_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__11010),
            .in2(_gnd_net_),
            .in3(N__10556),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__13673),
            .ce(),
            .sr(N__11908));
    defparam \this_vga_signals.M_hcounter_q_9_LC_14_16_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_9_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_9_LC_14_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_9_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__11745),
            .in2(_gnd_net_),
            .in3(N__10553),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_9 ),
            .clk(N__13677),
            .ce(),
            .sr(N__11906));
    defparam \this_vga_signals.M_hcounter_q_10_LC_14_16_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_10_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_10_LC_14_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_10_LC_14_16_1  (
            .in0(N__12224),
            .in1(N__11711),
            .in2(_gnd_net_),
            .in3(N__10550),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_10 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_9 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_10 ),
            .clk(N__13677),
            .ce(),
            .sr(N__11906));
    defparam \this_vga_signals.M_hcounter_q_11_LC_14_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_11_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_11_LC_14_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_11_LC_14_16_2  (
            .in0(N__12223),
            .in1(N__12489),
            .in2(_gnd_net_),
            .in3(N__10547),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13677),
            .ce(),
            .sr(N__11906));
    defparam \this_vga_signals.M_vcounter_q_0_LC_14_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_0_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_14_17_1 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_14_17_1  (
            .in0(N__10871),
            .in1(N__12011),
            .in2(N__11935),
            .in3(N__12225),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13682),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_2_0_LC_14_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_2_0_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_2_0_LC_14_17_2 .LUT_INIT=16'b0001000110001000;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_2_0_LC_14_17_2  (
            .in0(N__12111),
            .in1(N__11744),
            .in2(_gnd_net_),
            .in3(N__11493),
            .lcout(\this_vga_signals.M_hstate_q_ns_i_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_1_0_LC_14_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_1_0_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_1_0_LC_14_17_5 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_1_0_LC_14_17_5  (
            .in0(N__11255),
            .in1(N__11018),
            .in2(N__11714),
            .in3(N__11768),
            .lcout(),
            .ltout(\this_vga_signals.N_76_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_0_LC_14_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_0_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_0_LC_14_17_6 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_0_LC_14_17_6  (
            .in0(N__11769),
            .in1(N__10886),
            .in2(N__10877),
            .in3(N__12731),
            .lcout(),
            .ltout(\this_vga_signals.N_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_0_LC_14_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_0_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_0_LC_14_17_7 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \this_vga_signals.M_hstate_q_0_LC_14_17_7  (
            .in0(N__12066),
            .in1(N__12191),
            .in2(N__10874),
            .in3(N__11770),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13682),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_0_c_LC_14_18_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_0_c_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_0_c_LC_14_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_0_c_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__10870),
            .in2(N__12226),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_LUT4_0_LC_14_18_1 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_LUT4_0_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_LUT4_0_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_LUT4_0_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10844),
            .in3(N__10802),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_LUT4_0_LC_14_18_2 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_LUT4_0_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_LUT4_0_LC_14_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_LUT4_0_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__10798),
            .in2(_gnd_net_),
            .in3(N__10742),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_LUT4_0_LC_14_18_3 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_LUT4_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_LUT4_0_LC_14_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_LUT4_0_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__10738),
            .in2(_gnd_net_),
            .in3(N__10685),
            .lcout(\this_vga_signals.un1_M_vcounter_q_6_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_LC_14_18_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_4_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_LC_14_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__10671),
            .in2(_gnd_net_),
            .in3(N__10640),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_4 ),
            .clk(N__13685),
            .ce(),
            .sr(N__11905));
    defparam \this_vga_signals.M_vcounter_q_5_LC_14_18_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_5_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_LC_14_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__10632),
            .in2(_gnd_net_),
            .in3(N__10604),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_5 ),
            .clk(N__13685),
            .ce(),
            .sr(N__11905));
    defparam \this_vga_signals.M_vcounter_q_6_LC_14_18_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_6_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_LC_14_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__10591),
            .in2(_gnd_net_),
            .in3(N__10565),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_6 ),
            .clk(N__13685),
            .ce(),
            .sr(N__11905));
    defparam \this_vga_signals.M_vcounter_q_7_LC_14_18_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_7_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_LC_14_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__10963),
            .in2(_gnd_net_),
            .in3(N__10937),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_7 ),
            .clk(N__13685),
            .ce(),
            .sr(N__11905));
    defparam \this_vga_signals.M_vcounter_q_8_LC_14_19_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_8_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_LC_14_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__10922),
            .in2(_gnd_net_),
            .in3(N__10889),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8 ),
            .clk(N__13689),
            .ce(),
            .sr(N__11904));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_0_LC_14_19_1 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_0_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_0_LC_14_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_0_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__13017),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_8 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_1_LC_14_19_2 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_1_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_1_LC_14_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_1_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__13084),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_0_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_2_LC_14_19_3 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_2_LC_14_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_2_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__13021),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_1_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_3_LC_14_19_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_3_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_3_LC_14_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_3_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__13085),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_2_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_3_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_4_LC_14_19_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_4_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_4_LC_14_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_4_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__13025),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_3_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_4_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_5_LC_14_19_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_5_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_5_LC_14_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_5_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__13086),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_4_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_5_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_6_LC_14_19_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_6_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_6_LC_14_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_6_cry_8_c_THRU_CRY_6_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__13029),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_5_THRU_CO ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_6_cry_8_THRU_CRY_6_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_LC_14_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_LC_14_20_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_LC_14_20_0 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_LC_14_20_0  (
            .in0(N__11971),
            .in1(N__12017),
            .in2(N__11934),
            .in3(N__11990),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13693),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_15_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_15_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_15_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__11866),
            .in2(_gnd_net_),
            .in3(N__11832),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13669),
            .ce(),
            .sr(N__11907));
    defparam \this_vga_signals.M_hcounter_q_0_LC_15_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_15_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_15_15_6  (
            .in0(N__11867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13669),
            .ce(),
            .sr(N__11907));
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_1_LC_15_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_1_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_1_LC_15_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI2UC41_1_LC_15_16_0  (
            .in0(N__11864),
            .in1(N__11845),
            .in2(N__11833),
            .in3(N__11809),
            .lcout(\this_vga_signals.N_169_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNITMFU_0_9_LC_15_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNITMFU_0_9_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNITMFU_0_9_LC_15_16_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNITMFU_0_9_LC_15_16_3  (
            .in0(N__11704),
            .in1(_gnd_net_),
            .in2(N__11746),
            .in3(N__11486),
            .lcout(\this_vga_signals.N_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNID7PV_0_LC_15_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNID7PV_0_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNID7PV_0_LC_15_16_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \this_vga_signals.M_hstate_q_RNID7PV_0_LC_15_16_6  (
            .in0(N__11767),
            .in1(N__11250),
            .in2(_gnd_net_),
            .in3(N__11014),
            .lcout(\this_vga_signals.N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNITMFU_9_LC_15_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNITMFU_9_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNITMFU_9_LC_15_16_7 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNITMFU_9_LC_15_16_7  (
            .in0(N__11740),
            .in1(_gnd_net_),
            .in2(N__11713),
            .in3(N__11485),
            .lcout(\this_vga_signals.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_4_0_LC_15_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_4_0_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_4_0_LC_15_17_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_4_0_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__11259),
            .in2(_gnd_net_),
            .in3(N__11022),
            .lcout(),
            .ltout(\this_vga_signals.N_37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_3_0_LC_15_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_3_0_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_3_0_LC_15_17_1 .LUT_INIT=16'b0000101000000011;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_3_0_LC_15_17_1  (
            .in0(N__12151),
            .in1(N__12163),
            .in2(N__12734),
            .in3(N__12108),
            .lcout(\this_vga_signals.M_hstate_q_ns_i_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_15_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_15_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIQFS22_11_LC_15_17_2  (
            .in0(N__12539),
            .in1(N__12278),
            .in2(N__12491),
            .in3(N__12236),
            .lcout(\this_vga_signals.N_169 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIPU1C1_11_LC_15_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIPU1C1_11_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIPU1C1_11_LC_15_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIPU1C1_11_LC_15_17_3  (
            .in0(N__12540),
            .in1(N__12485),
            .in2(N__12288),
            .in3(N__12107),
            .lcout(),
            .ltout(\this_vga_signals.M_hstate_d_0_sqmuxa_0_a2_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_15_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_15_17_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI5RNE4_11_LC_15_17_4  (
            .in0(N__12175),
            .in1(N__12150),
            .in2(N__12239),
            .in3(N__12235),
            .lcout(\this_vga_signals.M_hstate_d_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_1_LC_15_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_1_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hstate_q_1_LC_15_17_5 .LUT_INIT=16'b0000011100000010;
    LogicCell40 \this_vga_signals.M_hstate_q_1_LC_15_17_5  (
            .in0(N__12187),
            .in1(N__12083),
            .in2(N__12065),
            .in3(N__12110),
            .lcout(\this_vga_signals.M_hstate_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13678),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_15_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hstate_q_RNO_0_1_LC_15_17_7 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \this_vga_signals.M_hstate_q_RNO_0_1_LC_15_17_7  (
            .in0(N__12176),
            .in1(N__12164),
            .in2(N__12155),
            .in3(N__12109),
            .lcout(\this_vga_signals.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_16_17_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_16_17_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__13758),
            .in2(_gnd_net_),
            .in3(N__13733),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13672),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_16_17_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_16_17_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__13760),
            .in2(_gnd_net_),
            .in3(N__12023),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13672),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_16_17_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_16_17_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_16_17_5  (
            .in0(N__13759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12029),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13672),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_16_17_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_16_17_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_16_17_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_16_17_7  (
            .in0(N__13757),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13672),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_2_RNI34P11_0_LC_17_16_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_2_RNI34P11_0_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_2_RNI34P11_0_LC_17_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vram.mem_mem_4_2_RNI34P11_0_LC_17_16_4  (
            .in0(N__13502),
            .in1(N__13490),
            .in2(_gnd_net_),
            .in3(N__14156),
            .lcout(),
            .ltout(\this_vram.mem_mem_4_2_RNI34P11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_radreg_RNIG1S72_11_LC_17_16_5 .C_ON=1'b0;
    defparam \this_vram.mem_radreg_RNIG1S72_11_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_radreg_RNIG1S72_11_LC_17_16_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \this_vram.mem_radreg_RNIG1S72_11_LC_17_16_5  (
            .in0(N__14009),
            .in1(_gnd_net_),
            .in2(N__13469),
            .in3(N__14406),
            .lcout(\this_vram.mem_N_2372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_0_wclke_0_a2_LC_19_18_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_0_wclke_0_a2_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_0_wclke_0_a2_LC_19_18_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vram.mem_mem_5_0_wclke_0_a2_LC_19_18_7  (
            .in0(N__14650),
            .in1(N__14870),
            .in2(N__13828),
            .in3(N__14802),
            .lcout(\this_vram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_22_5_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_22_5_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_22_5_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_22_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_2_RNI9H021_0_LC_23_21_4 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_2_RNI9H021_0_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_2_RNI9H021_0_LC_23_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_vram.mem_mem_8_2_RNI9H021_0_LC_23_21_4  (
            .in0(N__14478),
            .in1(N__12851),
            .in2(_gnd_net_),
            .in3(N__12836),
            .lcout(\this_vram.mem_mem_8_2_RNI9H021Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_1_RNI38R11_LC_24_13_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_1_RNI38R11_LC_24_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_1_RNI38R11_LC_24_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \this_vram.mem_mem_5_1_RNI38R11_LC_24_13_2  (
            .in0(N__14169),
            .in1(N__12809),
            .in2(_gnd_net_),
            .in3(N__12794),
            .lcout(\this_vram.mem_mem_5_1_RNI38RZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_1_RNI38R11_0_LC_24_13_3 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_1_RNI38R11_0_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_1_RNI38R11_0_LC_24_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_5_1_RNI38R11_0_LC_24_13_3  (
            .in0(N__12770),
            .in1(N__14168),
            .in2(_gnd_net_),
            .in3(N__12755),
            .lcout(\this_vram.mem_mem_5_1_RNI38R11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_6_0_wclke_0_a2_LC_24_15_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_6_0_wclke_0_a2_LC_24_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_6_0_wclke_0_a2_LC_24_15_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vram.mem_mem_6_0_wclke_0_a2_LC_24_15_0  (
            .in0(N__14800),
            .in1(N__14845),
            .in2(N__13804),
            .in3(N__14629),
            .lcout(\this_vram.mem_WE_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_2_RNI58R11_LC_24_15_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_2_RNI58R11_LC_24_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_2_RNI58R11_LC_24_15_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_5_2_RNI58R11_LC_24_15_1  (
            .in0(N__14225),
            .in1(N__14140),
            .in2(_gnd_net_),
            .in3(N__14216),
            .lcout(\this_vram.mem_mem_5_2_RNI58RZ0Z11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_5_2_RNI58R11_0_LC_24_15_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_5_2_RNI58R11_0_LC_24_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_5_2_RNI58R11_0_LC_24_15_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_5_2_RNI58R11_0_LC_24_15_2  (
            .in0(N__14183),
            .in1(N__14139),
            .in2(_gnd_net_),
            .in3(N__14024),
            .lcout(\this_vram.mem_mem_5_2_RNI58R11Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_7_0_wclke_0_a2_LC_24_15_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_7_0_wclke_0_a2_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_7_0_wclke_0_a2_LC_24_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vram.mem_mem_7_0_wclke_0_a2_LC_24_15_6  (
            .in0(N__14801),
            .in1(N__14846),
            .in2(N__13805),
            .in3(N__14630),
            .lcout(\this_vram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_0_RNI5H021_LC_24_17_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_0_RNI5H021_LC_24_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_0_RNI5H021_LC_24_17_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_8_0_RNI5H021_LC_24_17_1  (
            .in0(N__13964),
            .in1(N__14465),
            .in2(_gnd_net_),
            .in3(N__13952),
            .lcout(\this_vram.mem_mem_8_0_RNI5HZ0Z021 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_0_RNI5H021_0_LC_24_18_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_0_RNI5H021_0_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_0_RNI5H021_0_LC_24_18_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_8_0_RNI5H021_0_LC_24_18_6  (
            .in0(N__13931),
            .in1(N__14466),
            .in2(_gnd_net_),
            .in3(N__13925),
            .lcout(\this_vram.mem_mem_8_0_RNI5H021Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_1_RNI7H021_LC_24_19_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_1_RNI7H021_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_1_RNI7H021_LC_24_19_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vram.mem_mem_8_1_RNI7H021_LC_24_19_7  (
            .in0(N__13898),
            .in1(N__14467),
            .in2(_gnd_net_),
            .in3(N__13892),
            .lcout(\this_vram.mem_mem_8_1_RNI7HZ0Z021 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_4_0_wclke_0_a2_1_LC_24_20_0 .C_ON=1'b0;
    defparam \this_vram.mem_mem_4_0_wclke_0_a2_1_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_4_0_wclke_0_a2_1_LC_24_20_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vram.mem_mem_4_0_wclke_0_a2_1_LC_24_20_0  (
            .in0(N__14565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14697),
            .lcout(\this_vram.mem_N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_9_0_wclke_0_a2_LC_24_20_1 .C_ON=1'b0;
    defparam \this_vram.mem_mem_9_0_wclke_0_a2_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_9_0_wclke_0_a2_LC_24_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vram.mem_mem_9_0_wclke_0_a2_LC_24_20_1  (
            .in0(N__14699),
            .in1(N__14705),
            .in2(N__14570),
            .in3(N__14614),
            .lcout(\this_vram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_0_wclke_0_a2_0_LC_24_20_6 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_0_wclke_0_a2_0_LC_24_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_0_wclke_0_a2_0_LC_24_20_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vram.mem_mem_8_0_wclke_0_a2_0_LC_24_20_6  (
            .in0(N__14844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14767),
            .lcout(\this_vram.mem_N_29 ),
            .ltout(\this_vram.mem_N_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_0_wclke_0_a2_LC_24_20_7 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_0_wclke_0_a2_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_0_wclke_0_a2_LC_24_20_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vram.mem_mem_8_0_wclke_0_a2_LC_24_20_7  (
            .in0(N__14698),
            .in1(N__14613),
            .in2(N__14573),
            .in3(N__14566),
            .lcout(\this_vram.mem_WE_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_1_RNI7H021_0_LC_24_21_2 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_1_RNI7H021_0_LC_24_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_1_RNI7H021_0_LC_24_21_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \this_vram.mem_mem_8_1_RNI7H021_0_LC_24_21_2  (
            .in0(N__14513),
            .in1(N__14479),
            .in2(_gnd_net_),
            .in3(N__14501),
            .lcout(\this_vram.mem_mem_8_1_RNI7H021Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vram.mem_mem_8_2_RNI9H021_LC_24_21_5 .C_ON=1'b0;
    defparam \this_vram.mem_mem_8_2_RNI9H021_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vram.mem_mem_8_2_RNI9H021_LC_24_21_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \this_vram.mem_mem_8_2_RNI9H021_LC_24_21_5  (
            .in0(N__14480),
            .in1(_gnd_net_),
            .in2(N__14288),
            .in3(N__14279),
            .lcout(\this_vram.mem_mem_8_2_RNI9HZ0Z021 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
